
`default_nettype none

module my_chip (
    input logic [11:0] io_in,
    input logic clock, reset,
    output logic [11:0] io_out
);

wire [7:0] val;
reg [11:0] index;

always_ff @(posedge clock) begin
    index <= io_in;
    io_out <= {4'b0000, val};
end

assign val[0] = (~index[0] & index[1] & index[2] & index[3] & index[4] & ~index[8] & index[10]) | (~index[0] & index[1] & ~index[4] & ~index[5] & ~index[6] & index[7] & index[9] & ~index[10] & ~index[11]) | (index[0] & index[1] & index[3] & index[5] & ~index[6] & ~index[7]) | (index[0] & ~index[1] & ~index[3] & index[5] & index[6] & index[7] & ~index[8] & index[10]) | (~index[0] & index[1] & ~index[2] & index[4] & index[6] & index[8] & ~index[9] & index[10]) | (index[0] & ~index[1] & ~index[2] & ~index[3] & index[4] & index[7] & ~index[9] & ~index[10] & ~index[11]) | (~index[0] & index[1] & index[2] & index[5] & ~index[6] & ~index[8]) | (index[0] & index[1] & index[2] & ~index[3] & ~index[4] & ~index[5] & ~index[7] & index[8] & ~index[9] & index[10]) | (index[0] & ~index[1] & index[2] & index[3] & ~index[4] & ~index[5] & ~index[7] & index[9] & index[10]) | (~index[0] & index[3] & index[6] & index[7] & index[8] & ~index[10] & index[11]) | (~index[0] & ~index[1] & ~index[3] & ~index[6] & index[7] & ~index[8] & ~index[9] & index[10] & ~index[11]) | (index[0] & ~index[1] & ~index[2] & index[3] & index[4] & index[7] & index[8] & ~index[10] & index[11]) | (index[1] & index[2] & ~index[3] & ~index[4] & ~index[5] & index[6] & ~index[7] & index[10] & index[11]) | (index[0] & ~index[1] & index[2] & ~index[3] & index[5] & index[6] & index[7] & index[10] & ~index[11]) | (index[0] & index[1] & ~index[3] & index[5] & index[6] & ~index[7] & index[11]) | (~index[0] & index[1] & ~index[2] & ~index[3] & ~index[5] & index[6] & index[7] & ~index[8] & ~index[9]) | (index[1] & ~index[2] & ~index[4] & ~index[5] & index[6] & index[7] & ~index[8] & index[9] & index[10]) | (index[0] & index[3] & index[5] & index[9] & ~index[10]) | (index[0] & ~index[2] & ~index[4] & ~index[5] & ~index[7] & index[8] & ~index[9] & ~index[10] & ~index[11]) | (index[1] & index[2] & ~index[3] & index[4] & ~index[7] & ~index[8] & ~index[9] & index[10]) | (index[0] & ~index[3] & ~index[4] & ~index[6] & ~index[8] & index[9] & ~index[10] & ~index[11]) | (index[0] & ~index[1] & ~index[3] & ~index[5] & index[6] & ~index[7] & ~index[8] & index[9]) | (~index[0] & ~index[3] & index[4] & ~index[6] & index[7] & index[8] & index[9] & index[10] & ~index[11]) | (~index[0] & ~index[2] & ~index[3] & index[6] & ~index[7] & index[8] & index[9] & index[10] & index[11]) | (~index[0] & index[1] & index[2] & index[3] & ~index[6] & ~index[8] & ~index[9] & index[11]) | (~index[0] & index[1] & index[2] & ~index[3] & ~index[4] & index[7] & index[8] & ~index[9] & ~index[10] & ~index[11]) | (index[2] & index[3] & ~index[4] & ~index[6] & index[7] & ~index[8] & index[9] & ~index[10]) | (~index[0] & index[3] & ~index[4] & index[6] & index[7] & ~index[9] & index[11]) | (index[0] & ~index[1] & ~index[4] & index[6] & index[7] & index[8] & ~index[9] & index[10]) | (~index[0] & ~index[1] & ~index[3] & ~index[4] & ~index[5] & ~index[6] & index[8] & index[9] & index[10] & index[11]) | (index[0] & index[1] & ~index[4] & ~index[6] & index[7] & index[8] & index[9] & index[10] & ~index[11]) | (~index[1] & ~index[2] & index[4] & ~index[6] & index[7] & index[9] & ~index[10] & index[11]) | (~index[0] & index[2] & index[3] & ~index[4] & index[6] & index[8] & index[9] & index[10] & ~index[11]) | (~index[0] & index[2] & ~index[3] & ~index[4] & index[6] & ~index[7] & index[8] & ~index[10] & index[11]) | (~index[1] & ~index[2] & ~index[3] & index[4] & index[5] & ~index[7]) | (index[1] & index[4] & index[6] & index[7] & index[9] & ~index[10] & index[11]) | (index[0] & index[1] & ~index[2] & index[3] & ~index[6] & index[7] & index[9] & index[10] & ~index[11]) | (~index[1] & ~index[2] & index[3] & index[4] & index[6] & ~index[8] & ~index[9] & index[10]) | (index[0] & ~index[1] & index[2] & ~index[3] & index[4] & ~index[6] & ~index[7] & index[8] & index[10]) | (~index[0] & ~index[1] & index[2] & index[3] & index[4] & ~index[8] & index[9] & index[11]) | (index[0] & index[2] & ~index[3] & ~index[4] & ~index[5] & index[6] & index[7] & index[8] & index[11]) | (~index[0] & index[2] & ~index[4] & ~index[5] & ~index[6] & index[7] & index[8] & ~index[9] & index[10]) | (index[0] & ~index[1] & ~index[2] & index[5] & ~index[6] & index[7] & index[9] & ~index[11]) | (index[0] & ~index[1] & ~index[2] & ~index[3] & ~index[4] & ~index[5] & ~index[7] & ~index[8] & ~index[11]) | (index[0] & ~index[1] & index[2] & index[3] & ~index[4] & ~index[5] & index[7] & ~index[9] & index[10]) | (index[0] & ~index[1] & index[2] & index[3] & ~index[7] & index[8] & index[9] & index[10] & ~index[11]) | (~index[0] & index[2] & index[3] & ~index[4] & index[6] & ~index[7] & index[8] & index[9] & ~index[11]) | (~index[0] & index[1] & ~index[3] & ~index[6] & index[7] & index[8] & ~index[9] & index[11]) | (~index[0] & ~index[1] & index[2] & index[3] & ~index[4] & ~index[7] & ~index[10] & ~index[11]) | (index[0] & ~index[1] & index[2] & ~index[4] & ~index[5] & index[6] & ~index[7] & ~index[8] & index[10]) | (index[0] & ~index[1] & index[2] & ~index[3] & ~index[5] & index[6] & index[7] & index[8] & ~index[10] & ~index[11]) | (index[0] & index[1] & index[2] & index[3] & ~index[6] & ~index[7] & index[11]) | (~index[1] & ~index[2] & index[3] & index[6] & ~index[7] & ~index[8] & ~index[9] & index[10]) | (~index[0] & index[1] & index[2] & ~index[4] & ~index[6] & ~index[7] & ~index[8] & ~index[9] & index[11]) | (index[0] & index[1] & ~index[3] & ~index[4] & ~index[5] & index[6] & ~index[8] & ~index[10] & ~index[11]) | (~index[0] & index[1] & index[2] & index[4] & index[6] & ~index[7] & index[9] & ~index[10]) | (index[0] & ~index[1] & ~index[2] & index[4] & index[6] & ~index[7] & index[9] & index[11]) | (~index[0] & ~index[1] & index[2] & index[3] & index[4] & index[8] & ~index[9] & index[10]) | (~index[0] & ~index[1] & index[2] & index[4] & ~index[6] & ~index[8] & ~index[10] & ~index[11]) | (~index[0] & index[1] & index[2] & ~index[3] & index[4] & index[7] & ~index[8] & index[9] & index[11]) | (~index[0] & index[1] & ~index[2] & index[4] & ~index[5] & ~index[6] & index[8] & index[9] & index[10]) | (index[0] & index[1] & ~index[2] & ~index[3] & ~index[4] & ~index[5] & index[6] & index[8] & index[10] & ~index[11]) | (index[0] & index[1] & index[2] & ~index[3] & ~index[4] & ~index[5] & index[7] & ~index[8] & ~index[9] & ~index[11]) | (~index[0] & index[1] & index[2] & index[5] & ~index[6] & ~index[9] & index[10]) | (~index[0] & index[1] & ~index[2] & ~index[5] & ~index[6] & index[10] & index[11]) | (index[1] & ~index[3] & ~index[4] & ~index[8] & index[9] & ~index[10] & ~index[11]) | (index[0] & ~index[1] & index[4] & index[6] & index[7] & ~index[8] & index[9] & index[10]) | (index[0] & ~index[2] & ~index[3] & index[4] & index[6] & ~index[7] & ~index[10] & index[11]) | (index[0] & ~index[1] & ~index[2] & ~index[4] & ~index[6] & index[7] & index[10] & index[11]) | (~index[0] & ~index[1] & ~index[2] & ~index[4] & index[6] & ~index[7] & ~index[9] & ~index[10] & index[11]) | (~index[1] & index[3] & ~index[4] & ~index[7] & index[8] & ~index[9] & ~index[10] & ~index[11]) | (~index[1] & ~index[2] & index[3] & ~index[5] & index[6] & index[7] & index[8] & index[9] & index[10] & ~index[11]) | (~index[0] & index[1] & ~index[2] & index[3] & ~index[4] & ~index[5] & ~index[7] & ~index[8] & ~index[11]) | (~index[0] & index[1] & ~index[2] & ~index[3] & index[6] & index[10] & index[11]) | (index[0] & ~index[2] & ~index[3] & ~index[4] & index[6] & ~index[7] & index[8] & ~index[9]) | (index[0] & ~index[1] & index[4] & ~index[6] & index[7] & index[8] & ~index[9] & index[10]) | (~index[0] & ~index[1] & ~index[2] & ~index[3] & index[4] & ~index[6] & index[8] & ~index[9] & index[11]) | (index[0] & index[1] & ~index[2] & ~index[3] & index[4] & ~index[6] & index[8] & index[9] & ~index[10]) | (index[2] & index[4] & index[6] & ~index[7] & index[8] & ~index[9] & ~index[10] & ~index[11]) | (index[2] & index[3] & index[4] & ~index[7] & ~index[8] & ~index[10] & ~index[11]) | (~index[0] & ~index[2] & index[3] & ~index[5] & index[6] & ~index[7] & ~index[8] & ~index[9] & index[11]) | (index[0] & index[1] & ~index[2] & ~index[4] & index[6] & index[7] & index[8] & index[9] & ~index[10]) | (~index[0] & index[1] & ~index[2] & index[3] & ~index[4] & ~index[6] & index[9] & ~index[10]) | (~index[0] & ~index[1] & ~index[2] & ~index[3] & index[4] & index[6] & index[8] & ~index[10] & ~index[11]) | (~index[0] & ~index[1] & index[3] & index[5] & ~index[7] & ~index[8]) | (~index[0] & ~index[1] & index[2] & ~index[4] & ~index[5] & ~index[6] & index[10] & index[11]) | (~index[0] & ~index[1] & ~index[4] & ~index[6] & ~index[7] & index[8] & ~index[9] & ~index[10] & ~index[11]) | (index[0] & ~index[1] & index[2] & index[3] & ~index[4] & ~index[5] & index[8] & index[9] & index[10] & ~index[11]) | (index[0] & ~index[1] & index[3] & index[4] & index[6] & ~index[8] & index[11]) | (~index[0] & ~index[1] & ~index[3] & index[6] & index[7] & index[8] & ~index[9] & ~index[10] & ~index[11]) | (~index[0] & index[2] & index[4] & index[6] & index[7] & index[9] & ~index[10] & index[11]) | (~index[0] & ~index[1] & index[2] & index[5] & index[6] & ~index[9] & index[10]) | (~index[0] & ~index[1] & index[2] & index[3] & ~index[4] & index[6] & ~index[8] & index[11]) | (index[0] & ~index[1] & ~index[2] & ~index[3] & ~index[4] & ~index[5] & ~index[6] & index[8] & index[10] & ~index[11]) | (index[0] & index[1] & ~index[2] & index[3] & index[6] & ~index[7] & index[8] & ~index[10]) | (~index[0] & ~index[1] & ~index[2] & index[3] & index[6] & ~index[7] & ~index[8] & index[10]) | (index[0] & ~index[1] & index[2] & index[3] & ~index[5] & ~index[6] & index[7] & ~index[9] & index[10]) | (~index[2] & index[3] & index[4] & index[7] & index[9] & ~index[10] & index[11]) | (index[0] & ~index[2] & ~index[3] & ~index[4] & ~index[5] & index[6] & index[7] & index[8] & index[9] & ~index[11]) | (index[0] & ~index[1] & ~index[2] & index[3] & ~index[4] & ~index[5] & index[6] & index[9] & index[11]) | (index[0] & index[1] & ~index[2] & index[4] & index[6] & ~index[7] & ~index[8] & index[9] & index[10]) | (~index[0] & index[1] & ~index[3] & index[4] & ~index[5] & ~index[6] & index[7] & index[9] & index[10]) | (index[1] & index[2] & ~index[4] & ~index[7] & ~index[8] & ~index[10] & ~index[11]) | (~index[0] & index[1] & ~index[2] & index[4] & index[6] & index[7] & ~index[10] & ~index[11]) | (index[0] & index[1] & index[3] & index[4] & index[7] & ~index[9] & ~index[10] & ~index[11]) | (index[0] & index[1] & ~index[2] & ~index[3] & ~index[4] & ~index[6] & ~index[7] & ~index[8]) | (~index[0] & index[2] & index[3] & index[4] & index[6] & ~index[7] & index[9] & index[11]) | (~index[0] & index[2] & ~index[4] & ~index[6] & index[7] & index[8] & ~index[9] & index[11]) | (~index[0] & index[1] & ~index[2] & ~index[4] & ~index[5] & ~index[6] & ~index[7] & index[8] & index[11]) | (~index[0] & ~index[1] & index[3] & ~index[4] & ~index[5] & index[7] & ~index[9] & index[11]) | (index[0] & index[1] & index[3] & ~index[6] & ~index[7] & ~index[8] & ~index[9]) | (~index[0] & ~index[1] & ~index[2] & index[3] & index[4] & ~index[6] & ~index[7] & index[10] & index[11]) | (~index[0] & ~index[1] & index[2] & ~index[4] & index[6] & index[8] & ~index[9] & ~index[10] & ~index[11]) | (~index[0] & ~index[1] & index[2] & ~index[3] & ~index[4] & index[7] & ~index[8] & ~index[9] & index[10]) | (~index[0] & index[2] & index[5] & index[6] & ~index[7] & ~index[11]) | (~index[0] & ~index[1] & index[5] & ~index[7] & index[9] & ~index[11]) | (~index[1] & index[2] & index[3] & ~index[4] & index[7] & ~index[8] & index[9] & index[11]) | (index[0] & ~index[2] & index[3] & ~index[4] & index[6] & index[7] & index[9] & index[11]) | (~index[0] & index[1] & ~index[2] & ~index[3] & ~index[7] & index[10] & index[11]) | (~index[1] & index[2] & ~index[3] & index[6] & index[8] & ~index[9] & ~index[10] & ~index[11]) | (index[0] & index[2] & index[3] & index[5] & ~index[8] & index[9]) | (index[0] & ~index[1] & ~index[2] & index[3] & ~index[4] & index[6] & index[7] & index[8] & ~index[9] & ~index[11]) | (~index[0] & index[1] & ~index[2] & index[3] & index[5] & index[6] & index[10]) | (~index[1] & ~index[2] & ~index[4] & ~index[5] & ~index[6] & index[7] & ~index[9] & index[10] & ~index[11]) | (~index[0] & ~index[1] & index[3] & ~index[5] & index[6] & index[7] & index[8] & index[9] & ~index[11]) | (~index[0] & ~index[1] & ~index[2] & index[3] & ~index[6] & ~index[9] & ~index[10] & ~index[11]) | (index[0] & ~index[1] & index[2] & ~index[3] & index[4] & index[6] & index[7] & ~index[9] & ~index[11]) | (~index[0] & ~index[2] & index[4] & ~index[6] & ~index[7] & ~index[8] & index[9] & index[10]) | (index[0] & index[1] & index[2] & ~index[3] & ~index[5] & index[7] & index[10] & index[11]) | (index[0] & ~index[1] & ~index[2] & ~index[3] & ~index[4] & ~index[5] & index[7] & index[11]) | (index[0] & index[1] & index[2] & index[3] & ~index[4] & ~index[6] & ~index[7] & ~index[9]) | (~index[1] & index[2] & index[4] & index[5] & ~index[6]) | (index[1] & ~index[2] & ~index[3] & ~index[4] & ~index[5] & index[7] & ~index[8] & index[9] & ~index[11]) | (~index[0] & index[1] & index[2] & index[3] & index[4] & ~index[6] & ~index[7] & ~index[9]) | (~index[1] & index[2] & index[3] & ~index[4] & index[6] & ~index[7] & index[8] & index[9] & ~index[11]) | (index[0] & index[1] & index[2] & index[3] & ~index[7] & ~index[8] & ~index[10]) | (~index[0] & ~index[1] & index[2] & ~index[3] & index[6] & ~index[7] & index[8] & ~index[9] & ~index[10]) | (~index[0] & index[1] & index[2] & ~index[3] & ~index[5] & index[6] & ~index[8] & ~index[9] & index[11]) | (index[0] & ~index[1] & index[2] & index[3] & index[6] & ~index[7] & ~index[9] & index[11]) | (~index[0] & ~index[1] & index[3] & index[5] & ~index[7] & index[11]) | (index[0] & ~index[1] & ~index[2] & index[3] & index[5] & index[6] & ~index[9]) | (index[1] & index[2] & index[3] & ~index[6] & index[7] & index[8] & index[9] & ~index[11]) | (~index[0] & index[1] & index[2] & index[3] & ~index[4] & index[6] & index[7] & ~index[8] & ~index[9] & ~index[10]) | (~index[1] & index[2] & ~index[3] & ~index[4] & ~index[6] & ~index[7] & index[8] & index[9] & index[10] & ~index[11]) | (~index[0] & ~index[1] & index[2] & index[3] & index[4] & ~index[6] & index[8] & index[10] & ~index[11]) | (~index[0] & ~index[1] & ~index[2] & ~index[4] & ~index[5] & index[7] & ~index[8] & ~index[9] & index[10] & ~index[11]) | (index[0] & index[1] & ~index[2] & ~index[4] & ~index[6] & index[8] & ~index[9] & ~index[10] & ~index[11]) | (~index[0] & ~index[1] & ~index[2] & ~index[3] & ~index[4] & ~index[7] & index[8] & index[10] & ~index[11]) | (index[0] & ~index[3] & index[4] & ~index[6] & index[7] & ~index[8] & ~index[9] & index[11]) | (index[0] & ~index[1] & ~index[3] & ~index[6] & index[7] & index[8] & ~index[9] & ~index[10] & ~index[11]) | (~index[0] & ~index[2] & index[3] & index[4] & index[6] & index[7] & index[9] & ~index[10]) | (~index[0] & index[2] & ~index[4] & index[6] & index[7] & ~index[8] & ~index[9] & index[11]) | (~index[0] & ~index[1] & index[4] & ~index[6] & ~index[7] & index[8] & index[9] & ~index[10]) | (index[1] & ~index[2] & index[5] & index[6] & index[7] & index[8] & index[10] & ~index[11]) | (index[1] & ~index[2] & ~index[3] & index[4] & ~index[6] & ~index[7] & index[8] & index[9] & ~index[11]) | (~index[0] & ~index[1] & ~index[4] & ~index[5] & ~index[6] & index[7] & ~index[8] & ~index[9] & ~index[10]) | (~index[0] & index[1] & index[2] & index[4] & index[6] & index[7] & index[8] & ~index[9] & index[11]) | (~index[0] & ~index[1] & index[2] & ~index[4] & index[5] & index[6] & index[11]) | (index[0] & ~index[2] & ~index[3] & index[4] & index[6] & ~index[7] & index[9] & index[10] & ~index[11]) | (~index[1] & ~index[2] & index[4] & index[6] & index[7] & index[8] & ~index[9] & index[11]) | (index[0] & index[1] & index[2] & index[3] & ~index[4] & ~index[6] & ~index[8] & index[11]) | (index[1] & index[2] & ~index[3] & ~index[6] & index[7] & index[8] & ~index[9] & ~index[10] & ~index[11]) | (index[0] & index[1] & ~index[4] & ~index[5] & index[6] & index[7] & ~index[8] & index[9] & index[10]) | (index[0] & index[1] & ~index[5] & ~index[6] & ~index[7] & index[8] & ~index[10] & index[11]) | (~index[0] & index[1] & ~index[3] & index[4] & index[7] & ~index[8] & ~index[9] & ~index[11]) | (index[0] & index[1] & index[2] & ~index[3] & index[4] & index[6] & ~index[7] & ~index[9]) | (~index[0] & index[1] & ~index[2] & index[3] & index[4] & index[7] & index[8] & ~index[10]) | (index[0] & index[2] & index[3] & index[4] & ~index[6] & index[8] & ~index[10] & ~index[11]) | (~index[0] & ~index[1] & ~index[2] & index[3] & ~index[4] & ~index[5] & ~index[6] & index[8] & index[10] & ~index[11]) | (~index[0] & index[1] & ~index[2] & ~index[8] & index[9] & ~index[10] & ~index[11]) | (index[0] & index[1] & index[2] & ~index[3] & ~index[4] & ~index[8] & ~index[10] & ~index[11]) | (~index[0] & index[2] & index[3] & index[4] & index[6] & ~index[8] & index[9] & index[10]) | (~index[0] & ~index[2] & index[4] & ~index[5] & index[6] & index[7] & index[8] & index[10] & ~index[11]) | (index[0] & index[1] & index[2] & index[3] & index[4] & ~index[6] & index[8] & index[11]) | (~index[1] & index[2] & index[3] & ~index[4] & ~index[6] & ~index[7] & ~index[8] & index[9] & index[10]) | (~index[0] & index[2] & index[3] & index[4] & index[6] & index[7] & ~index[8] & index[10]) | (~index[0] & index[1] & ~index[2] & index[4] & index[6] & index[7] & index[8] & index[9]) | (~index[0] & ~index[1] & ~index[2] & index[3] & ~index[4] & ~index[6] & ~index[8] & index[11]) | (index[0] & index[2] & ~index[3] & ~index[5] & index[6] & index[7] & ~index[8] & index[9] & index[10]) | (~index[0] & ~index[1] & ~index[2] & index[3] & ~index[7] & ~index[8] & ~index[9] & index[11]) | (index[0] & index[1] & index[2] & ~index[3] & index[4] & index[7] & index[8] & index[9] & index[10]) | (~index[1] & ~index[2] & ~index[3] & ~index[4] & ~index[5] & index[6] & index[7] & ~index[8] & ~index[10] & index[11]) | (~index[1] & ~index[2] & index[5] & index[6] & ~index[7] & index[8] & index[10] & ~index[11]) | (index[0] & ~index[2] & ~index[3] & ~index[4] & index[5] & ~index[6] & index[10] & index[11]) | (index[0] & index[2] & index[3] & ~index[6] & index[7] & index[8] & index[10] & ~index[11]) | (index[0] & index[2] & ~index[4] & ~index[6] & index[7] & ~index[8] & index[9] & ~index[10]) | (index[0] & index[1] & ~index[2] & ~index[3] & ~index[5] & ~index[7] & ~index[9] & index[11]) | (~index[0] & ~index[2] & ~index[3] & ~index[5] & ~index[6] & ~index[7] & ~index[8] & index[9] & ~index[10] & index[11]) | (index[1] & ~index[2] & index[3] & ~index[4] & index[6] & ~index[7] & ~index[8] & index[9]) | (~index[0] & index[1] & ~index[2] & index[3] & ~index[6] & index[7] & index[8] & ~index[10] & ~index[11]) | (index[1] & index[2] & index[4] & ~index[6] & ~index[7] & index[8] & ~index[10] & index[11]) | (~index[0] & ~index[1] & index[3] & ~index[4] & ~index[5] & index[6] & index[9] & ~index[10] & ~index[11]) | (~index[0] & ~index[2] & index[4] & index[6] & ~index[7] & ~index[8] & ~index[9] & index[10]) | (~index[0] & ~index[1] & ~index[2] & index[3] & ~index[6] & index[7] & ~index[8] & index[9] & index[10]) | (~index[1] & index[2] & ~index[3] & ~index[4] & ~index[5] & index[6] & ~index[7] & ~index[8] & index[10]) | (index[0] & ~index[1] & index[2] & ~index[3] & ~index[4] & ~index[5] & index[7] & index[8] & ~index[10]) | (index[0] & index[1] & index[2] & ~index[5] & ~index[6] & ~index[7] & ~index[8] & index[9] & index[11]) | (~index[0] & index[1] & index[2] & index[3] & ~index[6] & ~index[8] & index[9] & index[10]) | (index[1] & index[2] & ~index[3] & index[5] & ~index[6] & index[7] & ~index[8] & ~index[9] & index[10]) | (~index[0] & index[1] & ~index[2] & ~index[3] & index[7] & ~index[8] & ~index[10] & ~index[11]) | (~index[0] & ~index[1] & index[2] & index[4] & ~index[7] & ~index[8] & ~index[10] & ~index[11]) | (index[0] & index[2] & ~index[3] & ~index[4] & ~index[6] & ~index[7] & index[8] & index[9] & ~index[10]) | (index[0] & index[1] & ~index[2] & ~index[4] & index[6] & index[8] & ~index[9] & index[10]) | (~index[0] & index[1] & ~index[3] & index[4] & index[6] & index[7] & index[8] & index[9] & ~index[10]) | (~index[0] & index[1] & index[2] & index[4] & ~index[6] & ~index[9] & ~index[10] & ~index[11]) | (~index[0] & index[1] & ~index[2] & index[3] & index[4] & index[6] & index[8] & ~index[11]) | (index[0] & index[1] & ~index[2] & index[3] & index[6] & index[7] & ~index[8] & index[11]) | (index[0] & ~index[1] & index[2] & ~index[4] & ~index[5] & ~index[6] & index[7] & ~index[8] & index[9]) | (~index[0] & ~index[1] & index[4] & ~index[6] & ~index[7] & index[8] & ~index[9] & index[10]) | (~index[0] & ~index[1] & ~index[2] & index[3] & index[6] & ~index[9] & index[11]) | (~index[0] & ~index[1] & ~index[2] & index[3] & ~index[4] & ~index[8] & ~index[9] & ~index[10]) | (~index[0] & ~index[1] & index[2] & ~index[3] & ~index[5] & index[7] & index[10] & index[11]) | (index[0] & index[1] & index[2] & index[3] & ~index[6] & index[7] & index[9] & ~index[10]) | (index[0] & index[2] & ~index[3] & ~index[6] & ~index[8] & index[9] & ~index[10] & ~index[11]) | (~index[0] & ~index[1] & index[2] & ~index[3] & ~index[4] & ~index[5] & index[6] & index[7] & index[8] & index[9] & index[10]) | (index[0] & ~index[1] & index[2] & ~index[3] & index[4] & index[8] & ~index[9] & ~index[11]) | (index[0] & index[1] & index[2] & ~index[8] & index[9] & ~index[10] & ~index[11]) | (~index[0] & index[1] & ~index[2] & index[5] & index[7] & ~index[9] & ~index[10]) | (index[0] & ~index[1] & ~index[2] & index[4] & ~index[6] & ~index[8] & index[9] & index[11]) | (~index[0] & ~index[1] & index[2] & index[4] & ~index[6] & ~index[7] & ~index[8] & index[11]) | (~index[0] & index[1] & ~index[3] & index[5] & ~index[7] & ~index[8] & ~index[9] & index[10]) | (index[0] & ~index[1] & ~index[2] & index[3] & ~index[4] & ~index[6] & index[7] & index[9] & ~index[10] & ~index[11]) | (~index[0] & index[1] & ~index[3] & ~index[5] & ~index[6] & ~index[7] & index[8] & index[9] & index[10] & ~index[11]) | (~index[0] & index[1] & ~index[2] & index[3] & index[6] & ~index[7] & index[8] & index[9] & index[10] & ~index[11]) | (index[0] & index[1] & ~index[2] & index[3] & ~index[4] & ~index[5] & index[7] & ~index[8] & index[10]) | (index[0] & index[1] & index[2] & ~index[3] & ~index[4] & ~index[7] & index[8] & index[9] & ~index[10]) | (index[0] & index[1] & index[3] & index[4] & index[6] & index[7] & ~index[8] & ~index[10]) | (index[0] & ~index[2] & ~index[3] & index[5] & ~index[8] & ~index[9] & index[11]) | (index[0] & ~index[1] & index[2] & ~index[3] & ~index[4] & ~index[6] & index[8] & ~index[10] & index[11]) | (index[0] & index[1] & ~index[2] & index[3] & ~index[5] & ~index[6] & ~index[9] & index[11]) | (~index[0] & ~index[1] & ~index[2] & index[5] & index[6] & ~index[8] & index[9]) | (~index[0] & ~index[1] & index[2] & ~index[3] & ~index[6] & ~index[7] & ~index[8] & index[9]) | (~index[1] & ~index[2] & index[5] & index[6] & index[8] & ~index[9]) | (index[0] & ~index[1] & ~index[3] & ~index[4] & ~index[5] & index[7] & index[9] & index[11]) | (index[0] & ~index[1] & index[3] & ~index[4] & ~index[6] & ~index[7] & ~index[8] & index[9]) | (~index[0] & index[1] & index[2] & ~index[3] & index[4] & index[6] & ~index[7] & index[9] & ~index[11]) | (~index[0] & ~index[1] & ~index[2] & ~index[3] & ~index[7] & index[8] & index[9] & ~index[10] & ~index[11]) | (index[0] & index[1] & index[3] & index[4] & ~index[6] & index[7] & index[8] & index[10]) | (~index[0] & index[1] & index[2] & index[3] & ~index[4] & ~index[6] & index[7] & index[9]) | (~index[0] & ~index[1] & index[5] & ~index[6] & index[7] & index[9] & ~index[10]) | (~index[0] & ~index[1] & ~index[2] & ~index[3] & index[4] & index[7] & index[8] & ~index[9] & ~index[10]) | (~index[0] & index[2] & index[3] & ~index[4] & ~index[5] & index[7] & ~index[10] & index[11]) | (~index[0] & ~index[1] & ~index[2] & index[5] & ~index[7] & index[8] & ~index[10]) | (~index[1] & ~index[2] & ~index[3] & index[4] & ~index[6] & ~index[7] & ~index[8] & ~index[9] & index[10]) | (~index[0] & index[1] & ~index[3] & ~index[4] & index[5] & ~index[6] & ~index[7] & index[10] & index[11]) | (index[1] & ~index[2] & ~index[3] & index[4] & ~index[6] & ~index[8] & ~index[9] & ~index[10]) | (index[1] & index[3] & index[5] & index[8] & index[10] & ~index[11]) | (~index[0] & index[1] & index[3] & ~index[5] & ~index[6] & index[7] & ~index[8] & ~index[9] & index[10]) | (index[0] & ~index[1] & index[2] & index[3] & index[4] & index[7] & index[10] & index[11]) | (~index[0] & index[1] & ~index[2] & ~index[3] & ~index[5] & index[6] & index[9] & index[11]) | (index[0] & index[2] & index[3] & index[4] & ~index[6] & ~index[7] & index[9] & ~index[11]) | (~index[0] & index[2] & index[3] & index[4] & index[7] & ~index[8] & index[9] & index[10]) | (index[0] & index[1] & ~index[2] & index[3] & ~index[4] & ~index[6] & index[9] & index[10] & ~index[11]) | (index[0] & index[2] & ~index[3] & index[6] & index[7] & index[8] & ~index[9] & index[10]) | (~index[1] & ~index[2] & index[3] & ~index[4] & index[7] & index[8] & ~index[9] & index[10]) | (~index[0] & index[3] & ~index[4] & ~index[5] & ~index[6] & index[7] & ~index[8] & index[11]) | (index[0] & index[1] & index[2] & index[3] & ~index[4] & index[6] & index[7] & index[8] & ~index[10]) | (index[0] & ~index[1] & index[2] & index[4] & index[6] & index[8] & ~index[9] & index[10]) | (index[0] & ~index[1] & index[2] & index[5] & ~index[6] & index[8] & ~index[9]) | (~index[0] & index[1] & ~index[2] & ~index[3] & ~index[5] & index[6] & index[7] & index[9] & ~index[10]) | (~index[0] & ~index[1] & ~index[4] & index[5] & index[6] & ~index[7] & index[10]) | (index[0] & ~index[1] & index[2] & ~index[3] & ~index[4] & index[5] & ~index[7] & index[8] & index[11]) | (index[0] & ~index[1] & ~index[2] & ~index[3] & ~index[7] & ~index[8] & ~index[10] & ~index[11]) | (~index[0] & index[1] & index[2] & index[5] & index[6] & index[9] & ~index[10]) | (index[0] & index[1] & ~index[2] & index[3] & index[6] & ~index[7] & index[8] & ~index[9]) | (index[2] & index[3] & ~index[4] & index[6] & index[7] & index[8] & ~index[9] & index[11]) | (~index[1] & ~index[2] & index[3] & ~index[4] & ~index[5] & ~index[6] & index[7] & ~index[8] & ~index[9]) | (index[0] & ~index[1] & ~index[3] & ~index[4] & ~index[5] & ~index[6] & ~index[7] & ~index[9] & index[10]) | (~index[1] & ~index[3] & index[5] & ~index[7] & index[8] & ~index[9] & index[10]) | (index[0] & index[1] & index[4] & index[5] & index[7]) | (~index[0] & ~index[2] & index[5] & index[7] & index[8] & ~index[9] & ~index[11]) | (~index[0] & ~index[1] & ~index[2] & index[4] & index[6] & index[7] & ~index[9] & index[11]) | (~index[0] & ~index[1] & index[2] & ~index[3] & index[4] & ~index[8] & index[9] & ~index[10] & ~index[11]) | (~index[0] & ~index[1] & ~index[2] & ~index[3] & ~index[4] & index[5] & index[8] & ~index[11]) | (~index[0] & index[1] & index[2] & ~index[4] & index[6] & ~index[7] & index[8] & ~index[9] & index[10]) | (index[0] & ~index[1] & ~index[3] & index[4] & ~index[5] & index[6] & index[10] & index[11]) | (index[0] & index[1] & index[2] & ~index[3] & index[6] & ~index[7] & ~index[9] & index[10]) | (~index[0] & index[1] & index[2] & index[3] & ~index[5] & index[6] & ~index[7] & index[10] & index[11]) | (index[0] & index[1] & ~index[2] & index[3] & ~index[4] & ~index[6] & ~index[8] & index[10]) | (~index[0] & index[2] & ~index[3] & index[5] & index[7] & ~index[8] & index[10]) | (index[1] & ~index[2] & ~index[3] & index[4] & index[6] & index[7] & ~index[9] & index[10]) | (~index[0] & index[1] & index[2] & ~index[3] & ~index[5] & ~index[6] & index[7] & index[8] & ~index[10]) | (index[0] & index[1] & ~index[2] & index[4] & ~index[6] & index[8] & ~index[9] & index[10]) | (~index[0] & ~index[1] & index[2] & index[3] & ~index[4] & ~index[6] & ~index[9] & index[10]) | (index[0] & ~index[1] & ~index[2] & ~index[3] & index[4] & index[6] & index[7] & ~index[8] & ~index[11]) | (~index[0] & ~index[2] & ~index[3] & ~index[6] & ~index[7] & index[8] & index[9] & ~index[11]) | (index[0] & ~index[2] & ~index[3] & ~index[4] & ~index[5] & ~index[6] & ~index[7] & ~index[8] & ~index[9]) | (~index[0] & index[1] & ~index[2] & ~index[3] & ~index[5] & ~index[6] & ~index[7] & ~index[9] & ~index[11]) | (index[0] & ~index[1] & ~index[2] & index[4] & index[6] & ~index[7] & index[9] & ~index[10]);

assign val[1] = (~index[0] & index[1] & ~index[2] & ~index[4] & ~index[6] & index[7] & index[8] & index[10] & ~index[11]) | (index[0] & index[1] & ~index[4] & index[6] & ~index[7] & index[8] & ~index[9] & index[10]) | (~index[0] & ~index[1] & ~index[2] & index[3] & index[4] & index[6] & index[7] & ~index[8] & index[10]) | (index[0] & index[1] & ~index[2] & index[4] & ~index[7] & ~index[8] & index[9] & index[11]) | (index[0] & index[1] & index[2] & index[3] & index[4] & ~index[7] & index[8] & ~index[10]) | (index[0] & index[5] & index[7] & ~index[8] & index[9] & index[11]) | (index[0] & ~index[2] & index[3] & index[4] & ~index[7] & index[8] & index[9] & index[10] & ~index[11]) | (index[1] & index[2] & index[3] & ~index[6] & ~index[7] & ~index[8] & index[9] & index[11]) | (index[1] & ~index[2] & ~index[3] & index[4] & ~index[6] & index[7] & ~index[8] & index[9] & index[10]) | (index[0] & index[2] & index[3] & ~index[4] & ~index[6] & ~index[7] & ~index[8] & index[9]) | (~index[0] & ~index[1] & ~index[2] & ~index[3] & index[4] & index[6] & ~index[7] & index[8] & ~index[10]) | (index[0] & ~index[1] & index[2] & ~index[3] & ~index[6] & index[7] & index[9] & ~index[10] & index[11]) | (index[1] & ~index[2] & ~index[5] & index[6] & index[7] & ~index[8] & ~index[9] & index[11]) | (~index[0] & index[1] & ~index[2] & index[3] & index[5] & index[6] & index[9] & index[11]) | (~index[0] & index[1] & ~index[4] & ~index[6] & ~index[7] & ~index[8] & ~index[9] & index[11]) | (~index[0] & index[1] & ~index[2] & ~index[3] & index[5] & ~index[6] & index[7] & ~index[8] & index[9] & index[10]) | (~index[0] & ~index[1] & ~index[3] & ~index[4] & ~index[6] & index[7] & index[8] & index[9] & index[10] & index[11]) | (index[1] & ~index[2] & ~index[3] & ~index[4] & ~index[5] & ~index[7] & ~index[8] & index[9]) | (~index[0] & index[1] & index[2] & index[4] & index[6] & index[7] & ~index[8] & ~index[10] & ~index[11]) | (index[0] & ~index[1] & ~index[2] & ~index[3] & ~index[5] & ~index[6] & index[7] & ~index[8] & index[9] & index[10]) | (~index[0] & ~index[1] & index[2] & index[3] & ~index[4] & ~index[5] & index[6] & index[7] & ~index[8] & index[10]) | (index[0] & index[1] & index[3] & ~index[4] & index[7] & index[8] & ~index[10] & index[11]) | (~index[0] & ~index[1] & index[2] & index[3] & index[4] & ~index[6] & index[8] & index[9]) | (index[0] & index[1] & index[2] & index[3] & ~index[4] & index[7] & index[8] & ~index[9] & ~index[10]) | (index[0] & index[1] & ~index[2] & index[3] & ~index[4] & index[6] & index[7] & index[8] & ~index[10]) | (index[0] & ~index[1] & ~index[2] & index[3] & ~index[4] & ~index[6] & index[7] & ~index[8] & index[9] & ~index[10]) | (~index[1] & index[3] & ~index[4] & ~index[6] & ~index[7] & ~index[8] & index[9] & index[10]) | (index[0] & index[1] & index[2] & ~index[3] & index[4] & ~index[6] & ~index[7] & ~index[9] & index[10]) | (~index[0] & index[1] & ~index[2] & index[4] & index[7] & ~index[9] & index[11]) | (~index[0] & ~index[1] & index[3] & index[5] & ~index[6] & index[7] & ~index[11]) | (index[0] & index[2] & ~index[4] & ~index[6] & index[7] & index[9] & ~index[10] & index[11]) | (index[0] & index[1] & ~index[3] & index[4] & ~index[6] & ~index[7] & ~index[8] & index[9] & index[10]) | (index[0] & index[1] & index[2] & ~index[3] & index[6] & ~index[7] & ~index[8] & ~index[9] & index[11]) | (index[0] & ~index[1] & ~index[2] & index[3] & index[4] & index[7] & index[8] & index[9] & ~index[10]) | (~index[0] & ~index[1] & ~index[2] & ~index[3] & index[4] & index[7] & index[8] & index[9] & index[10] & ~index[11]) | (~index[0] & ~index[1] & index[2] & ~index[4] & ~index[6] & ~index[8] & index[9] & index[10]) | (~index[0] & ~index[1] & index[2] & ~index[3] & ~index[4] & index[5] & index[9] & index[11]) | (~index[1] & index[2] & index[3] & ~index[4] & ~index[6] & ~index[8] & index[9] & index[10]) | (index[0] & index[1] & index[2] & ~index[3] & ~index[5] & ~index[6] & index[7] & index[10] & index[11]) | (~index[0] & index[2] & ~index[3] & index[4] & index[6] & ~index[7] & ~index[8] & index[9] & index[10]) | (index[0] & ~index[1] & index[2] & index[3] & index[4] & index[6] & index[7] & index[10] & ~index[11]) | (~index[2] & index[3] & index[5] & index[7] & index[10] & index[11]) | (index[1] & index[2] & index[3] & index[4] & index[6] & index[7] & index[8] & index[11]) | (~index[0] & ~index[1] & ~index[2] & ~index[3] & ~index[5] & index[6] & ~index[8] & ~index[9] & ~index[10] & ~index[11]) | (~index[0] & index[1] & ~index[2] & ~index[3] & ~index[4] & ~index[5] & ~index[6] & ~index[7] & ~index[10]) | (~index[0] & ~index[1] & index[2] & index[6] & index[7] & index[8] & ~index[9] & index[10]) | (~index[0] & index[1] & index[2] & index[4] & ~index[6] & ~index[7] & ~index[8] & ~index[9] & index[10]) | (~index[0] & ~index[1] & index[2] & index[3] & ~index[4] & ~index[5] & index[6] & ~index[8] & ~index[9] & index[10]) | (index[0] & index[1] & ~index[2] & ~index[3] & index[4] & index[7] & index[8] & index[9] & ~index[11]) | (~index[2] & ~index[3] & ~index[4] & ~index[5] & ~index[6] & index[7] & index[8] & ~index[9] & index[10] & ~index[11]) | (index[0] & index[2] & ~index[4] & index[6] & index[7] & index[8] & ~index[9] & index[11]) | (index[0] & index[1] & ~index[3] & ~index[4] & index[6] & ~index[7] & ~index[9] & index[10]) | (~index[0] & ~index[2] & index[3] & index[4] & ~index[6] & index[8] & ~index[9] & index[11]) | (index[0] & ~index[1] & ~index[2] & ~index[3] & index[4] & ~index[7] & ~index[8] & ~index[9] & index[10]) | (~index[0] & ~index[1] & index[2] & index[4] & index[6] & ~index[7] & ~index[8] & index[9] & index[10]) | (index[0] & ~index[1] & ~index[2] & ~index[3] & ~index[4] & ~index[5] & index[6] & index[7] & ~index[10] & ~index[11]) | (~index[0] & index[1] & ~index[3] & ~index[4] & ~index[7] & ~index[8] & ~index[10] & ~index[11]) | (~index[0] & index[1] & index[2] & index[3] & index[4] & index[6] & ~index[7] & index[8] & index[10]) | (index[0] & index[2] & ~index[3] & ~index[4] & ~index[5] & index[6] & index[9] & ~index[10] & ~index[11]) | (~index[0] & index[1] & ~index[2] & index[4] & index[5] & index[7]) | (~index[0] & index[2] & index[3] & index[4] & ~index[6] & index[7] & ~index[8] & index[10]) | (index[0] & index[2] & index[3] & ~index[4] & index[7] & ~index[8] & index[9] & index[11]) | (~index[0] & ~index[2] & index[3] & index[5] & index[9] & ~index[10]) | (index[0] & ~index[1] & index[2] & ~index[3] & index[4] & ~index[6] & index[7] & ~index[8] & index[10]) | (~index[0] & index[1] & index[3] & index[4] & index[6] & index[7] & index[11]) | (index[0] & ~index[1] & index[2] & index[3] & ~index[4] & ~index[7] & ~index[8] & ~index[9] & index[11]) | (index[0] & ~index[1] & index[2] & ~index[3] & index[4] & index[6] & index[7] & ~index[9] & index[11]) | (~index[0] & index[2] & index[3] & index[4] & index[6] & index[9] & index[11]) | (~index[0] & ~index[1] & ~index[3] & index[5] & index[6] & index[7] & ~index[9] & index[10]) | (~index[1] & index[2] & ~index[3] & index[5] & index[6] & index[8] & ~index[10]) | (~index[0] & ~index[1] & index[2] & ~index[3] & ~index[4] & ~index[6] & index[7] & index[8] & index[11]) | (~index[0] & index[1] & ~index[2] & index[3] & ~index[4] & ~index[6] & index[7] & index[8] & ~index[11]) | (index[0] & index[1] & ~index[2] & index[3] & ~index[4] & ~index[6] & ~index[8] & ~index[9] & index[10]) | (index[0] & ~index[1] & ~index[2] & index[3] & index[4] & ~index[7] & index[9] & index[11]) | (index[0] & ~index[1] & index[2] & index[5] & ~index[7] & ~index[9] & index[10]) | (index[0] & index[1] & ~index[3] & ~index[4] & ~index[5] & ~index[7] & index[9] & ~index[10] & index[11]) | (~index[0] & index[1] & ~index[3] & ~index[4] & ~index[5] & ~index[6] & ~index[7] & index[8] & index[9] & ~index[11]) | (index[0] & ~index[1] & ~index[2] & ~index[5] & index[6] & index[7] & index[8] & index[9] & ~index[10]) | (index[0] & index[1] & index[3] & index[4] & ~index[6] & ~index[8] & ~index[10] & ~index[11]) | (~index[0] & index[1] & ~index[2] & index[3] & ~index[5] & ~index[6] & ~index[7] & index[8] & index[11]) | (~index[1] & index[2] & index[5] & ~index[7] & ~index[8] & ~index[9] & index[10]) | (~index[0] & index[2] & index[4] & index[6] & index[7] & index[9] & ~index[10] & index[11]) | (index[0] & index[1] & ~index[3] & ~index[6] & ~index[8] & ~index[9] & ~index[10] & ~index[11]) | (~index[0] & ~index[2] & index[3] & ~index[4] & ~index[5] & index[6] & index[7] & ~index[9] & ~index[10] & ~index[11]) | (~index[1] & ~index[2] & index[4] & ~index[6] & ~index[7] & ~index[8] & index[9] & index[11]) | (~index[0] & ~index[1] & ~index[2] & index[3] & ~index[4] & ~index[6] & ~index[7] & ~index[9] & ~index[10] & ~index[11]) | (index[1] & ~index[2] & index[4] & ~index[6] & index[7] & index[8] & ~index[10] & index[11]) | (~index[0] & ~index[2] & index[3] & index[4] & index[7] & ~index[9] & index[11]) | (~index[0] & index[1] & ~index[2] & index[3] & index[4] & ~index[6] & ~index[7] & ~index[9] & index[10]) | (~index[0] & index[2] & index[4] & index[5] & index[6]) | (~index[0] & index[1] & ~index[2] & ~index[3] & index[4] & ~index[6] & index[8] & ~index[9] & index[10]) | (~index[0] & ~index[3] & index[5] & ~index[6] & ~index[8] & ~index[9] & index[11]) | (index[0] & ~index[1] & index[2] & index[3] & ~index[4] & ~index[6] & index[7] & index[11]) | (~index[0] & index[1] & ~index[2] & ~index[3] & index[4] & ~index[6] & ~index[8] & ~index[9] & index[11]) | (~index[0] & ~index[2] & index[3] & index[6] & ~index[7] & index[8] & ~index[9] & index[10]) | (~index[0] & ~index[1] & ~index[2] & index[4] & index[5] & ~index[6] & ~index[7]) | (index[0] & ~index[1] & ~index[2] & ~index[4] & index[6] & ~index[7] & index[9] & ~index[10] & index[11]) | (~index[0] & index[1] & index[2] & index[3] & ~index[4] & index[6] & index[9] & ~index[10]) | (~index[0] & index[2] & ~index[3] & index[4] & ~index[6] & index[8] & index[9] & index[10] & ~index[11]) | (index[1] & ~index[2] & index[3] & index[4] & index[6] & ~index[7] & index[8] & index[9] & ~index[10]) | (index[0] & ~index[1] & index[2] & index[3] & ~index[4] & index[6] & index[8] & index[9] & index[10] & ~index[11]) | (~index[1] & index[2] & ~index[3] & ~index[4] & ~index[5] & ~index[6] & ~index[7] & index[9] & index[10] & ~index[11]) | (index[0] & ~index[1] & ~index[2] & ~index[3] & ~index[5] & index[7] & index[10] & index[11]) | (~index[0] & index[1] & index[2] & ~index[3] & index[6] & index[10] & index[11]) | (~index[0] & index[1] & index[2] & index[3] & index[4] & index[7] & ~index[8] & index[9] & index[10]) | (~index[0] & ~index[1] & index[2] & index[3] & ~index[4] & ~index[6] & ~index[7] & index[8] & ~index[9] & index[11]) | (~index[1] & ~index[2] & ~index[3] & index[4] & ~index[6] & ~index[7] & ~index[9] & ~index[10] & ~index[11]) | (~index[0] & index[2] & ~index[3] & ~index[4] & ~index[5] & ~index[6] & index[7] & index[8] & index[9] & ~index[10]) | (~index[0] & index[1] & index[2] & ~index[3] & index[4] & ~index[7] & index[8] & ~index[9] & ~index[10] & ~index[11]) | (~index[1] & ~index[2] & index[3] & ~index[4] & ~index[5] & index[6] & index[7] & ~index[8] & ~index[9] & index[10]) | (~index[1] & index[2] & ~index[3] & index[6] & index[7] & index[8] & ~index[9] & index[10]) | (index[0] & index[2] & index[3] & ~index[4] & index[6] & index[7] & ~index[9] & ~index[10] & ~index[11]) | (index[0] & index[1] & index[2] & index[3] & index[4] & index[6] & ~index[7] & ~index[8] & index[10]) | (index[0] & ~index[1] & ~index[2] & index[3] & index[4] & ~index[7] & ~index[8] & index[11]) | (index[0] & ~index[2] & index[3] & ~index[4] & index[6] & ~index[7] & ~index[8] & index[9] & index[10]) | (~index[0] & ~index[1] & index[2] & index[3] & index[4] & ~index[6] & index[9] & index[10]) | (index[0] & ~index[1] & ~index[3] & index[4] & index[6] & ~index[8] & ~index[9] & index[10]) | (index[0] & ~index[1] & ~index[2] & index[3] & index[4] & index[6] & index[9] & index[11]) | (index[0] & ~index[1] & index[2] & ~index[3] & index[5] & ~index[6] & ~index[8] & ~index[9] & index[10]) | (~index[0] & index[1] & index[2] & index[3] & index[5] & ~index[6] & ~index[7]) | (index[0] & ~index[1] & index[2] & ~index[4] & ~index[6] & ~index[7] & index[10] & index[11]) | (index[0] & ~index[1] & index[2] & index[3] & ~index[4] & ~index[6] & ~index[8] & ~index[9] & ~index[10]) | (index[0] & ~index[1] & index[2] & index[3] & ~index[6] & index[7] & index[8] & ~index[9] & index[10]) | (~index[0] & ~index[1] & ~index[2] & index[3] & ~index[5] & index[6] & ~index[7] & ~index[8] & ~index[9] & index[11]) | (index[0] & ~index[1] & ~index[3] & ~index[4] & index[7] & index[8] & ~index[9] & ~index[10] & ~index[11]) | (index[0] & index[2] & index[4] & ~index[6] & ~index[7] & index[8] & index[9] & ~index[10]) | (~index[0] & ~index[1] & index[2] & ~index[3] & ~index[4] & index[6] & ~index[7] & index[9] & index[11]) | (index[0] & ~index[1] & ~index[3] & ~index[4] & index[5] & ~index[6] & ~index[7] & index[10] & index[11]) | (~index[0] & index[1] & ~index[2] & index[3] & index[6] & ~index[7] & ~index[8] & index[9] & index[10]) | (~index[0] & ~index[1] & index[2] & ~index[3] & ~index[5] & index[6] & ~index[7] & ~index[8] & ~index[9] & index[11]) | (index[0] & ~index[1] & ~index[2] & ~index[3] & index[5] & index[6] & ~index[7] & index[11]) | (~index[0] & ~index[1] & ~index[2] & ~index[4] & ~index[6] & index[7] & ~index[8] & ~index[9] & ~index[10] & index[11]) | (index[1] & ~index[2] & index[3] & ~index[4] & ~index[5] & ~index[7] & index[10] & index[11]) | (index[0] & index[1] & index[2] & index[4] & ~index[6] & index[7] & index[8] & ~index[10] & ~index[11]) | (index[0] & index[1] & index[2] & index[3] & index[4] & index[9] & ~index[10]) | (~index[0] & ~index[2] & ~index[3] & ~index[4] & ~index[5] & ~index[6] & ~index[7] & index[8] & ~index[9] & ~index[10] & index[11]) | (~index[0] & ~index[1] & ~index[2] & ~index[3] & ~index[5] & index[6] & ~index[7] & index[8] & index[9] & ~index[10] & ~index[11]) | (index[0] & ~index[2] & ~index[3] & index[4] & index[6] & index[7] & index[9] & ~index[10] & ~index[11]) | (index[0] & ~index[1] & ~index[2] & ~index[3] & ~index[5] & index[6] & ~index[7] & index[8] & index[10] & ~index[11]) | (~index[1] & index[2] & index[3] & index[4] & index[6] & index[7] & index[8] & index[9] & ~index[10]) | (~index[0] & ~index[1] & ~index[2] & index[3] & ~index[4] & index[7] & index[10] & index[11]) | (index[0] & ~index[1] & ~index[2] & index[3] & index[6] & index[7] & index[8] & ~index[9] & index[10]) | (~index[0] & index[1] & index[2] & ~index[3] & ~index[4] & ~index[5] & index[6] & index[7] & ~index[9] & ~index[10] & ~index[11]) | (index[0] & index[1] & index[5] & ~index[6] & index[7] & ~index[10]) | (index[0] & ~index[1] & index[2] & index[3] & ~index[6] & index[7] & index[10] & index[11]) | (~index[0] & index[1] & index[2] & index[6] & index[7] & index[9] & index[11]) | (~index[0] & index[1] & ~index[3] & index[4] & ~index[6] & index[7] & index[8] & ~index[9] & index[10]) | (~index[0] & index[1] & ~index[2] & ~index[3] & ~index[4] & ~index[5] & index[6] & index[7] & index[10] & ~index[11]) | (index[0] & index[2] & index[4] & ~index[6] & ~index[7] & ~index[8] & ~index[9] & index[11]) | (index[0] & ~index[1] & ~index[2] & ~index[3] & ~index[4] & ~index[6] & index[7] & index[8] & ~index[9]) | (index[1] & index[2] & ~index[3] & ~index[4] & ~index[5] & ~index[6] & index[8] & ~index[10] & index[11]) | (index[0] & index[2] & ~index[3] & ~index[4] & index[6] & ~index[7] & ~index[8] & ~index[9] & index[10]) | (index[0] & ~index[1] & ~index[2] & index[3] & index[4] & ~index[6] & index[7] & ~index[8] & ~index[9] & index[10]) | (~index[0] & index[1] & index[2] & ~index[3] & ~index[4] & ~index[5] & index[7] & ~index[8] & index[9] & index[10]) | (index[0] & ~index[1] & ~index[3] & index[4] & index[6] & ~index[7] & index[8] & index[9] & index[10] & ~index[11]) | (index[0] & ~index[1] & ~index[2] & ~index[3] & ~index[4] & ~index[5] & ~index[6] & index[8] & index[9] & ~index[10]) | (index[0] & ~index[1] & index[2] & index[4] & index[7] & index[8] & ~index[9] & index[10]) | (index[0] & ~index[2] & ~index[3] & ~index[4] & index[6] & index[9] & ~index[10] & index[11]) | (~index[0] & ~index[1] & index[2] & ~index[3] & index[4] & ~index[6] & ~index[8] & index[9] & ~index[10] & ~index[11]) | (~index[0] & index[1] & ~index[2] & index[4] & ~index[5] & ~index[6] & ~index[7] & index[10] & index[11]) | (index[1] & ~index[2] & ~index[3] & index[4] & ~index[6] & index[8] & index[9] & ~index[10]) | (~index[0] & ~index[1] & ~index[2] & ~index[3] & index[4] & ~index[6] & ~index[7] & ~index[9] & ~index[11]) | (index[0] & ~index[1] & ~index[2] & ~index[3] & index[4] & ~index[8] & index[9] & ~index[10] & ~index[11]) | (index[0] & index[2] & index[3] & index[4] & ~index[7] & index[8] & ~index[9] & index[11]) | (index[0] & ~index[1] & index[2] & ~index[3] & index[6] & index[8] & index[9] & ~index[10]) | (index[0] & index[1] & ~index[2] & index[3] & ~index[4] & ~index[6] & index[9] & index[11]) | (~index[0] & index[1] & index[2] & index[3] & index[4] & index[6] & ~index[8] & ~index[10] & ~index[11]) | (~index[0] & index[1] & ~index[2] & ~index[4] & ~index[5] & ~index[7] & ~index[8] & index[9] & index[10]) | (~index[0] & ~index[1] & ~index[2] & ~index[3] & index[5] & ~index[7] & index[8] & index[10] & ~index[11]) | (index[0] & ~index[1] & ~index[2] & index[3] & index[4] & index[6] & index[7] & index[8] & ~index[10] & ~index[11]) | (~index[0] & index[1] & ~index[2] & index[3] & index[4] & index[6] & index[7] & index[8] & index[10]) | (~index[0] & index[1] & ~index[2] & index[3] & ~index[4] & ~index[6] & index[7] & ~index[9] & ~index[11]) | (index[0] & ~index[2] & ~index[3] & ~index[5] & index[6] & index[7] & ~index[8] & ~index[9] & index[10]) | (~index[0] & ~index[2] & ~index[3] & ~index[4] & ~index[5] & index[6] & index[7] & ~index[8] & index[9] & index[10] & ~index[11]) | (index[1] & index[3] & index[4] & index[7] & ~index[8] & ~index[9] & ~index[10] & ~index[11]) | (~index[0] & ~index[1] & index[2] & index[4] & index[5] & index[7]) | (index[0] & ~index[2] & index[3] & ~index[4] & ~index[7] & ~index[8] & ~index[10] & ~index[11]) | (~index[0] & ~index[1] & index[2] & index[3] & index[4] & ~index[6] & index[7] & index[8] & index[11]) | (~index[0] & index[2] & index[3] & index[4] & index[7] & ~index[8] & ~index[9] & ~index[10] & ~index[11]) | (index[1] & index[2] & ~index[3] & index[5] & index[6] & index[9] & index[11]) | (index[0] & ~index[2] & ~index[3] & index[5] & index[6] & ~index[7] & index[9] & index[11]) | (~index[0] & ~index[1] & ~index[2] & ~index[3] & index[4] & ~index[7] & ~index[8] & index[9] & index[10]) | (~index[0] & index[1] & index[2] & index[5] & index[6] & index[7] & index[8] & index[10]) | (~index[0] & index[1] & index[2] & ~index[3] & ~index[4] & ~index[5] & ~index[7] & index[8] & ~index[9] & index[10]) | (index[0] & ~index[2] & index[5] & ~index[7] & ~index[8] & index[9] & index[10]) | (~index[0] & index[1] & index[2] & index[4] & ~index[6] & ~index[7] & index[9] & ~index[10] & index[11]) | (index[1] & index[2] & index[3] & ~index[6] & index[7] & index[8] & index[9] & ~index[10]) | (~index[0] & ~index[1] & index[2] & index[3] & ~index[4] & ~index[6] & ~index[8] & index[9] & ~index[11]) | (index[1] & ~index[2] & ~index[3] & ~index[4] & ~index[5] & ~index[6] & ~index[7] & index[9] & index[10] & ~index[11]) | (~index[0] & index[2] & ~index[3] & index[6] & ~index[7] & index[8] & ~index[9] & index[10]) | (~index[0] & index[1] & ~index[2] & index[3] & index[4] & index[7] & ~index[9] & ~index[10]) | (index[1] & index[2] & index[3] & index[4] & ~index[6] & ~index[7] & index[11]) | (index[0] & index[1] & ~index[2] & ~index[3] & index[6] & ~index[7] & index[8] & ~index[10] & index[11]) | (index[0] & index[1] & ~index[2] & ~index[4] & ~index[5] & index[6] & ~index[7] & index[8] & index[11]) | (~index[0] & index[1] & ~index[2] & ~index[4] & ~index[6] & index[7] & index[8] & ~index[9] & ~index[11]) | (~index[0] & ~index[1] & index[2] & ~index[3] & ~index[4] & index[6] & ~index[7] & index[8] & ~index[9] & ~index[11]) | (~index[0] & ~index[1] & ~index[2] & index[3] & index[4] & ~index[6] & index[7] & index[8] & ~index[9] & index[10]) | (index[0] & ~index[1] & index[2] & index[3] & index[4] & ~index[6] & ~index[7] & ~index[8] & index[10]) | (~index[0] & ~index[1] & ~index[2] & ~index[3] & index[4] & ~index[6] & index[7] & index[8] & ~index[10] & ~index[11]) | (index[0] & index[1] & ~index[2] & ~index[3] & ~index[6] & index[7] & index[8] & index[9] & ~index[10]) | (~index[0] & ~index[1] & ~index[2] & ~index[3] & ~index[4] & ~index[5] & ~index[6] & index[8] & index[9] & index[10] & index[11]) | (~index[0] & index[1] & ~index[2] & ~index[3] & ~index[4] & index[5] & ~index[6] & ~index[7] & index[9] & index[11]) | (~index[2] & ~index[3] & ~index[4] & ~index[5] & index[6] & ~index[7] & ~index[8] & index[9] & ~index[10] & index[11]) | (~index[0] & ~index[1] & ~index[2] & index[3] & ~index[6] & index[7] & ~index[8] & ~index[9] & ~index[10]) | (index[0] & index[1] & index[3] & ~index[4] & index[6] & index[7] & ~index[9] & index[11]) | (index[0] & index[3] & index[5] & ~index[7] & ~index[11]) | (~index[1] & ~index[2] & ~index[3] & ~index[5] & index[6] & index[7] & index[8] & index[9] & index[10] & index[11]) | (index[0] & ~index[1] & ~index[2] & ~index[3] & ~index[5] & ~index[6] & index[7] & ~index[8] & ~index[9] & index[11]) | (~index[0] & ~index[1] & ~index[2] & ~index[4] & index[6] & index[7] & ~index[8] & index[9] & ~index[10]) | (index[0] & ~index[2] & index[3] & ~index[4] & index[6] & index[8] & ~index[10] & index[11]) | (~index[0] & ~index[1] & ~index[3] & index[4] & index[6] & ~index[8] & index[9] & index[10]) | (~index[0] & ~index[1] & ~index[3] & index[4] & index[6] & ~index[7] & ~index[9] & index[11]) | (~index[1] & ~index[3] & ~index[4] & index[6] & index[7] & ~index[8] & index[9] & ~index[10] & ~index[11]) | (index[0] & index[2] & index[3] & index[4] & ~index[8] & index[9] & ~index[10] & ~index[11]) | (~index[0] & index[1] & ~index[3] & ~index[4] & ~index[6] & ~index[8] & index[9] & ~index[10] & ~index[11]) | (index[0] & index[1] & ~index[2] & ~index[3] & index[5] & index[6] & index[7] & ~index[8]) | (index[1] & ~index[2] & ~index[3] & index[5] & ~index[7] & ~index[9] & index[10]) | (index[1] & index[2] & index[3] & index[6] & ~index[7] & index[8] & ~index[9] & ~index[10] & ~index[11]) | (~index[0] & index[1] & ~index[3] & ~index[5] & ~index[6] & ~index[7] & index[8] & index[9] & index[10] & ~index[11]) | (~index[0] & index[2] & index[3] & ~index[4] & index[6] & ~index[7] & index[8] & index[9] & ~index[10]) | (~index[0] & index[1] & index[2] & ~index[3] & index[4] & index[6] & index[7] & index[8] & index[9] & index[10]) | (~index[0] & ~index[1] & index[2] & index[3] & index[4] & ~index[6] & ~index[7] & index[8] & index[10]) | (index[0] & index[1] & index[2] & index[5] & ~index[6] & index[9] & ~index[11]) | (index[0] & index[3] & ~index[4] & ~index[5] & ~index[6] & ~index[7] & index[10] & index[11]) | (index[0] & index[1] & ~index[3] & index[5] & index[6] & ~index[9] & index[10]) | (~index[0] & index[1] & index[2] & ~index[4] & ~index[6] & ~index[8] & ~index[9] & index[11]) | (index[0] & index[1] & ~index[2] & index[3] & ~index[4] & ~index[5] & index[6] & index[8] & index[9] & ~index[11]) | (index[0] & index[1] & index[2] & index[3] & index[4] & ~index[6] & ~index[8] & index[11]) | (index[0] & ~index[2] & index[3] & index[4] & index[6] & ~index[7] & ~index[8] & ~index[9] & index[10]) | (index[0] & ~index[1] & index[2] & ~index[4] & ~index[6] & ~index[7] & ~index[9] & ~index[10] & ~index[11]) | (index[0] & ~index[3] & index[4] & ~index[5] & ~index[6] & ~index[7] & index[10] & index[11]) | (index[0] & index[2] & index[3] & index[4] & index[6] & index[7] & index[8] & index[9] & ~index[11]) | (index[0] & index[1] & index[2] & index[3] & ~index[4] & ~index[7] & ~index[8] & ~index[9] & ~index[11]) | (~index[0] & index[1] & index[2] & ~index[3] & index[5] & ~index[6] & index[7] & ~index[8] & ~index[9]) | (index[1] & index[3] & index[4] & index[6] & index[7] & index[10] & index[11]) | (~index[0] & ~index[1] & ~index[3] & ~index[6] & ~index[7] & ~index[8] & index[9] & ~index[10] & index[11]) | (index[0] & index[2] & ~index[3] & index[4] & ~index[5] & ~index[6] & index[10] & index[11]) | (~index[0] & ~index[1] & index[2] & ~index[3] & ~index[4] & ~index[5] & index[7] & index[8] & ~index[9] & index[10]) | (index[0] & index[1] & index[2] & ~index[3] & ~index[5] & index[6] & index[7] & ~index[8] & index[9] & index[10]) | (index[0] & ~index[2] & ~index[4] & ~index[5] & ~index[6] & index[7] & index[10] & index[11]) | (~index[0] & ~index[1] & index[4] & index[6] & ~index[7] & ~index[8] & ~index[9] & index[11]) | (~index[0] & index[1] & ~index[2] & ~index[3] & index[4] & ~index[6] & index[7] & ~index[10] & index[11]) | (index[0] & ~index[1] & index[2] & index[5] & index[7] & index[8] & ~index[10]) | (index[0] & ~index[1] & index[2] & index[3] & ~index[4] & ~index[5] & ~index[7] & index[10] & index[11]) | (~index[0] & ~index[1] & ~index[2] & ~index[3] & ~index[6] & ~index[7] & index[8] & ~index[9] & index[10] & ~index[11]) | (index[0] & ~index[1] & index[5] & index[6] & index[7] & ~index[8] & index[11]) | (~index[0] & index[1] & index[3] & ~index[4] & index[6] & ~index[8] & index[9] & ~index[10] & ~index[11]) | (index[0] & index[2] & index[4] & index[6] & index[7] & index[8] & index[9] & ~index[10]) | (~index[0] & ~index[1] & ~index[2] & ~index[4] & index[6] & ~index[7] & index[8] & ~index[9] & ~index[10] & index[11]) | (~index[0] & index[2] & ~index[3] & ~index[4] & index[6] & index[10] & index[11]) | (~index[0] & index[1] & index[2] & index[3] & ~index[4] & index[6] & index[7] & index[8] & index[9]) | (~index[0] & ~index[1] & ~index[2] & index[4] & index[6] & index[7] & index[9] & index[10] & ~index[11]) | (~index[0] & index[1] & ~index[2] & ~index[3] & ~index[4] & ~index[5] & ~index[6] & ~index[7] & ~index[8]) | (index[0] & index[1] & index[2] & ~index[4] & ~index[5] & index[6] & ~index[8] & ~index[9] & ~index[10] & ~index[11]) | (index[0] & index[1] & index[2] & index[3] & ~index[4] & index[6] & index[8] & ~index[9] & ~index[11]) | (index[0] & index[1] & index[3] & ~index[4] & ~index[5] & ~index[6] & ~index[7] & index[8] & index[9]) | (index[0] & ~index[2] & ~index[3] & ~index[4] & ~index[6] & index[7] & ~index[9] & ~index[10] & ~index[11]) | (index[0] & index[2] & ~index[3] & ~index[4] & ~index[5] & index[7] & index[8] & index[9] & index[10] & ~index[11]) | (~index[0] & index[1] & ~index[2] & ~index[4] & ~index[5] & index[6] & ~index[8] & index[9] & index[10]) | (index[1] & index[2] & ~index[3] & index[4] & index[6] & ~index[7] & ~index[8] & ~index[9] & index[11]) | (~index[0] & index[3] & index[4] & ~index[6] & index[7] & ~index[8] & index[9] & index[10]) | (index[0] & ~index[1] & index[3] & index[5] & index[6] & index[7] & ~index[9]) | (~index[0] & index[1] & ~index[4] & ~index[5] & index[6] & ~index[7] & ~index[8] & index[9] & index[10]) | (~index[0] & index[1] & index[2] & index[3] & ~index[4] & ~index[6] & index[8] & ~index[9] & index[10]) | (~index[0] & ~index[1] & ~index[2] & index[3] & index[4] & ~index[6] & index[7] & ~index[8] & index[9]) | (index[0] & ~index[1] & index[2] & ~index[3] & index[4] & index[7] & index[8] & ~index[10] & index[11]) | (~index[0] & index[1] & ~index[2] & index[3] & index[4] & index[7] & index[8] & index[11]) | (~index[0] & index[1] & ~index[2] & ~index[3] & index[4] & index[6] & ~index[7] & ~index[8] & ~index[9] & index[10]) | (~index[0] & ~index[1] & ~index[2] & index[4] & index[6] & ~index[7] & ~index[8] & ~index[9] & ~index[10]) | (~index[0] & index[1] & ~index[2] & index[5] & index[6] & index[7] & index[9] & ~index[10]) | (~index[0] & ~index[1] & index[2] & ~index[3] & index[4] & index[6] & index[7] & index[8] & ~index[9] & ~index[11]) | (~index[0] & index[1] & index[4] & index[6] & index[7] & ~index[8] & ~index[9] & ~index[10] & ~index[11]) | (~index[0] & ~index[1] & ~index[2] & index[3] & index[4] & index[6] & ~index[7] & index[8] & index[9]) | (index[0] & ~index[1] & ~index[2] & ~index[4] & ~index[6] & index[7] & index[8] & ~index[9] & index[10]);

assign val[2] = (index[0] & ~index[2] & ~index[4] & index[6] & ~index[7] & index[8] & ~index[9] & index[10]) | (index[1] & ~index[2] & ~index[3] & index[4] & ~index[6] & ~index[8] & index[9] & index[10]) | (index[0] & ~index[1] & index[2] & ~index[3] & ~index[4] & ~index[5] & index[7] & ~index[8] & index[11]) | (~index[1] & ~index[2] & index[3] & ~index[4] & ~index[5] & ~index[6] & ~index[7] & index[8] & index[10] & ~index[11]) | (index[1] & index[2] & index[3] & index[4] & index[6] & index[7] & ~index[10] & index[11]) | (~index[0] & index[1] & index[2] & index[3] & ~index[6] & index[7] & index[9] & index[10] & ~index[11]) | (~index[1] & ~index[2] & index[3] & index[5] & ~index[10]) | (index[1] & index[2] & index[3] & ~index[4] & index[7] & index[9] & ~index[10] & index[11]) | (~index[0] & ~index[1] & ~index[4] & ~index[5] & ~index[6] & index[7] & index[9] & ~index[10] & ~index[11]) | (index[0] & index[2] & ~index[3] & index[4] & ~index[6] & ~index[7] & index[8] & ~index[9] & ~index[10]) | (index[0] & index[1] & ~index[2] & ~index[4] & ~index[6] & ~index[7] & ~index[9] & ~index[10] & ~index[11]) | (index[1] & ~index[2] & ~index[3] & ~index[4] & ~index[5] & index[6] & index[7] & ~index[8] & ~index[9] & ~index[10]) | (~index[1] & index[2] & ~index[3] & ~index[4] & index[7] & ~index[8] & index[9] & index[11]) | (index[0] & ~index[1] & index[3] & ~index[4] & ~index[6] & ~index[7] & index[8] & index[10] & ~index[11]) | (~index[0] & index[1] & ~index[2] & index[3] & ~index[4] & index[8] & ~index[10] & ~index[11]) | (~index[0] & index[1] & ~index[2] & ~index[4] & ~index[5] & index[6] & index[8] & index[9]) | (~index[0] & ~index[1] & ~index[3] & index[6] & ~index[7] & index[8] & ~index[9] & ~index[10] & ~index[11]) | (index[0] & index[1] & ~index[3] & index[4] & index[7] & index[8] & index[9] & index[10] & ~index[11]) | (index[0] & index[1] & index[2] & index[3] & index[5] & index[11]) | (~index[0] & index[2] & index[3] & ~index[6] & index[7] & index[8] & ~index[9] & index[11]) | (~index[0] & ~index[1] & index[3] & index[4] & index[6] & index[8] & ~index[9] & index[10]) | (~index[0] & index[2] & ~index[3] & index[5] & ~index[6] & index[7] & ~index[8] & index[11]) | (index[1] & index[2] & index[3] & index[6] & index[7] & index[8] & ~index[9] & index[11]) | (index[0] & index[1] & ~index[2] & index[5] & ~index[6] & ~index[8] & ~index[9]) | (~index[0] & ~index[1] & index[2] & index[3] & ~index[4] & index[6] & ~index[8] & ~index[9] & index[11]) | (index[0] & index[1] & index[2] & ~index[3] & ~index[4] & ~index[5] & index[7] & index[9] & index[10]) | (index[0] & ~index[2] & ~index[3] & ~index[4] & ~index[5] & ~index[6] & index[7] & ~index[9] & index[10]) | (index[0] & index[1] & index[2] & index[3] & ~index[6] & ~index[7] & ~index[8] & index[9] & index[11]) | (~index[1] & index[3] & index[4] & index[5]) | (~index[0] & index[1] & index[2] & index[3] & ~index[6] & ~index[7] & ~index[8] & ~index[9]) | (index[1] & ~index[2] & ~index[3] & ~index[4] & ~index[6] & ~index[7] & index[10] & index[11]) | (~index[0] & index[1] & index[4] & index[6] & index[7] & index[8] & ~index[9] & ~index[10] & ~index[11]) | (index[0] & index[1] & ~index[2] & ~index[3] & index[4] & ~index[6] & index[9] & ~index[10] & index[11]) | (index[0] & ~index[1] & index[2] & ~index[3] & ~index[4] & ~index[5] & index[10] & index[11]) | (index[0] & index[1] & ~index[2] & ~index[4] & ~index[5] & index[6] & index[7] & ~index[8] & index[11]) | (~index[0] & ~index[1] & index[2] & ~index[3] & index[4] & index[6] & index[7] & ~index[9] & ~index[11]) | (~index[0] & ~index[1] & ~index[3] & ~index[4] & ~index[5] & ~index[6] & ~index[7] & index[9] & index[10] & ~index[11]) | (index[1] & index[3] & ~index[4] & index[6] & index[7] & index[8] & index[9] & ~index[10]) | (~index[1] & index[2] & ~index[3] & index[6] & ~index[7] & index[8] & ~index[9] & ~index[10] & ~index[11]) | (index[0] & index[1] & ~index[2] & index[3] & index[4] & index[6] & ~index[7] & index[8] & index[10]) | (~index[0] & index[2] & index[3] & ~index[4] & index[6] & ~index[7] & index[8] & ~index[9] & ~index[11]) | (index[0] & index[1] & index[2] & ~index[3] & ~index[4] & ~index[7] & index[8] & ~index[9] & index[11]) | (index[0] & index[1] & ~index[2] & index[4] & index[6] & ~index[7] & index[8] & index[9] & index[10]) | (~index[0] & ~index[1] & index[2] & index[3] & index[4] & index[6] & ~index[7] & index[10]) | (~index[0] & ~index[1] & ~index[3] & ~index[4] & index[5] & ~index[6] & index[7] & index[9] & index[11]) | (index[0] & ~index[1] & index[3] & ~index[4] & ~index[5] & index[6] & ~index[7] & index[10] & index[11]) | (~index[0] & ~index[2] & ~index[3] & index[4] & ~index[5] & index[6] & ~index[7] & index[10] & index[11]) | (index[0] & index[2] & index[5] & index[6] & ~index[7] & ~index[9]) | (~index[0] & index[2] & ~index[3] & ~index[4] & ~index[5] & ~index[6] & ~index[7] & index[8] & index[10]) | (~index[0] & ~index[1] & ~index[2] & index[3] & ~index[4] & index[6] & ~index[7] & index[8] & ~index[9]) | (~index[0] & index[1] & ~index[2] & ~index[4] & index[6] & ~index[7] & ~index[8] & ~index[9] & index[10]) | (~index[1] & index[3] & index[4] & ~index[6] & ~index[7] & ~index[9] & ~index[10] & ~index[11]) | (~index[0] & ~index[1] & ~index[3] & index[4] & ~index[6] & index[7] & index[8] & ~index[9] & ~index[11]) | (index[0] & ~index[1] & ~index[2] & index[4] & index[6] & ~index[7] & ~index[8] & ~index[9] & index[11]) | (index[0] & index[1] & index[2] & index[5] & ~index[7] & ~index[9]) | (~index[1] & index[2] & ~index[3] & ~index[4] & ~index[5] & index[6] & index[7] & index[9] & ~index[10]) | (~index[0] & index[1] & ~index[2] & ~index[3] & ~index[7] & ~index[8] & ~index[9] & index[10]) | (index[0] & ~index[1] & index[2] & ~index[3] & index[4] & ~index[7] & ~index[8] & index[9] & index[10]) | (~index[0] & ~index[1] & ~index[2] & index[5] & ~index[7] & ~index[8] & index[10]) | (~index[0] & ~index[2] & ~index[3] & index[4] & ~index[6] & ~index[8] & index[9] & index[10]) | (index[0] & index[1] & index[2] & ~index[4] & ~index[6] & ~index[7] & index[8] & ~index[10] & index[11]) | (~index[0] & index[1] & index[2] & index[3] & index[4] & index[8] & ~index[9] & ~index[10]) | (index[0] & index[1] & index[2] & ~index[4] & index[6] & ~index[7] & ~index[8] & ~index[9] & ~index[11]) | (index[0] & index[1] & index[2] & index[3] & ~index[7] & ~index[8] & ~index[9] & index[10]) | (~index[0] & index[2] & ~index[4] & ~index[5] & ~index[6] & ~index[7] & index[10] & index[11]) | (~index[0] & ~index[1] & ~index[2] & index[3] & ~index[4] & ~index[6] & index[7] & ~index[8] & index[9]) | (index[0] & index[2] & index[3] & ~index[4] & ~index[7] & ~index[8] & ~index[10] & ~index[11]) | (~index[1] & index[2] & index[3] & index[4] & ~index[8] & ~index[9] & ~index[10] & ~index[11]) | (index[1] & ~index[2] & ~index[3] & index[4] & ~index[7] & ~index[8] & ~index[9] & index[10]) | (~index[1] & index[2] & index[3] & index[4] & ~index[6] & ~index[7] & ~index[8] & index[9] & index[10]) | (~index[0] & index[1] & ~index[2] & ~index[3] & ~index[4] & ~index[5] & index[6] & index[9] & index[11]) | (~index[0] & index[1] & ~index[2] & ~index[4] & ~index[5] & index[6] & index[7] & index[9] & index[10]) | (~index[2] & index[4] & ~index[6] & ~index[8] & ~index[9] & ~index[10] & ~index[11]) | (index[0] & index[1] & index[3] & index[4] & index[6] & index[7] & ~index[8] & ~index[9] & ~index[10]) | (index[0] & index[1] & index[2] & ~index[3] & index[6] & index[8] & ~index[9] & index[10]) | (~index[0] & ~index[1] & index[2] & index[4] & index[7] & index[8] & index[10] & ~index[11]) | (index[1] & ~index[2] & index[3] & ~index[4] & index[6] & index[7] & index[8] & ~index[10]) | (~index[0] & index[3] & ~index[4] & ~index[6] & index[7] & ~index[8] & index[9] & ~index[10]) | (~index[0] & ~index[1] & ~index[2] & index[4] & index[6] & index[7] & index[8] & index[9] & ~index[10]) | (~index[0] & index[2] & index[5] & index[7] & index[8] & ~index[9] & index[10]) | (index[1] & ~index[2] & index[3] & index[5] & index[7] & index[9] & index[11]) | (~index[0] & ~index[1] & index[2] & index[3] & ~index[4] & ~index[5] & index[6] & index[8] & ~index[10] & ~index[11]) | (~index[0] & ~index[1] & index[2] & index[3] & index[6] & index[7] & ~index[8] & ~index[9]) | (~index[0] & index[1] & ~index[3] & ~index[4] & ~index[5] & ~index[6] & ~index[9] & index[10]) | (index[0] & ~index[1] & ~index[2] & ~index[3] & ~index[4] & ~index[5] & index[6] & ~index[8] & index[10]) | (index[0] & ~index[1] & index[2] & ~index[6] & ~index[7] & index[8] & index[9] & ~index[10]) | (index[1] & index[2] & index[4] & ~index[6] & ~index[9] & ~index[10] & ~index[11]) | (~index[0] & index[1] & index[2] & ~index[4] & ~index[5] & index[7] & ~index[8] & ~index[9] & index[10]) | (index[0] & ~index[1] & index[2] & index[4] & ~index[6] & index[8] & ~index[10] & ~index[11]) | (~index[0] & index[2] & index[3] & index[4] & ~index[7] & ~index[9] & ~index[10] & ~index[11]) | (index[0] & ~index[1] & index[2] & index[5] & ~index[6] & index[9] & ~index[10]) | (~index[0] & index[2] & ~index[3] & index[4] & ~index[6] & index[7] & index[8] & index[9] & ~index[11]) | (index[0] & index[1] & ~index[2] & ~index[3] & ~index[7] & index[8] & ~index[9] & ~index[10] & ~index[11]) | (index[0] & index[1] & index[3] & index[4] & ~index[6] & index[7] & index[8] & ~index[10] & index[11]) | (~index[1] & index[2] & index[6] & index[7] & index[8] & ~index[9] & index[10]) | (~index[0] & index[1] & ~index[2] & ~index[3] & index[4] & ~index[6] & ~index[8] & ~index[9]) | (index[0] & ~index[2] & index[3] & ~index[4] & ~index[5] & index[6] & index[7] & ~index[8] & ~index[9] & index[10]) | (~index[0] & ~index[2] & ~index[3] & index[4] & index[7] & ~index[8] & index[9] & index[10]) | (index[0] & ~index[1] & ~index[2] & ~index[5] & index[6] & ~index[7] & ~index[8] & ~index[9] & index[10]) | (~index[1] & ~index[2] & index[3] & ~index[4] & ~index[6] & ~index[8] & ~index[10] & ~index[11]) | (~index[0] & ~index[1] & ~index[3] & ~index[4] & ~index[5] & index[7] & ~index[8] & index[9] & index[10] & ~index[11]) | (~index[0] & index[1] & ~index[3] & ~index[4] & ~index[5] & ~index[7] & index[9] & index[11]) | (index[0] & ~index[1] & ~index[2] & index[3] & index[5] & ~index[6] & index[11]) | (index[0] & index[2] & ~index[3] & ~index[5] & index[6] & index[7] & index[10] & index[11]) | (~index[0] & index[2] & index[3] & ~index[4] & ~index[5] & ~index[6] & ~index[8] & ~index[9] & index[10]) | (index[1] & index[2] & index[3] & index[4] & ~index[7] & index[8] & ~index[10] & ~index[11]) | (~index[1] & ~index[2] & ~index[3] & index[4] & ~index[6] & ~index[7] & index[8] & ~index[9] & ~index[10]) | (~index[1] & index[3] & ~index[4] & ~index[5] & ~index[7] & index[8] & ~index[9] & index[10]) | (index[1] & index[2] & ~index[3] & index[4] & index[6] & ~index[7] & ~index[8] & ~index[10]) | (~index[0] & ~index[1] & index[2] & ~index[3] & index[4] & ~index[6] & index[9] & ~index[10] & ~index[11]) | (index[0] & ~index[1] & ~index[2] & ~index[4] & ~index[7] & ~index[8] & index[9] & index[10]) | (~index[0] & ~index[1] & index[2] & ~index[3] & ~index[4] & ~index[5] & ~index[7] & index[9] & index[10] & ~index[11]) | (index[0] & index[1] & index[2] & index[5] & index[6] & ~index[8] & ~index[11]) | (index[1] & ~index[2] & ~index[3] & ~index[4] & ~index[5] & index[6] & index[8] & index[9] & ~index[11]) | (~index[0] & ~index[1] & ~index[3] & ~index[4] & ~index[5] & index[6] & ~index[7] & ~index[9] & ~index[10] & ~index[11]) | (index[1] & index[2] & index[3] & ~index[4] & index[6] & ~index[7] & ~index[8] & ~index[9] & index[11]) | (~index[0] & ~index[1] & ~index[3] & index[5] & index[6] & ~index[7] & index[8] & index[10]) | (~index[0] & index[1] & ~index[2] & ~index[4] & ~index[5] & ~index[6] & ~index[7] & index[8] & index[11]) | (~index[0] & index[2] & ~index[3] & index[4] & index[6] & index[7] & ~index[8] & ~index[9] & ~index[11]) | (~index[1] & index[2] & ~index[3] & ~index[5] & index[7] & index[8] & ~index[9] & index[10]) | (~index[0] & index[1] & index[3] & index[4] & index[6] & ~index[7] & index[8] & ~index[9] & index[11]) | (~index[0] & index[1] & ~index[2] & ~index[3] & ~index[4] & ~index[5] & ~index[6] & index[7] & ~index[9]) | (~index[1] & index[2] & index[3] & ~index[4] & ~index[6] & index[8] & ~index[10] & index[11]) | (index[0] & ~index[1] & ~index[2] & ~index[3] & ~index[4] & ~index[5] & ~index[6] & index[11]) | (index[0] & ~index[1] & index[5] & index[6] & ~index[7] & index[9] & ~index[10]) | (index[1] & ~index[2] & index[4] & ~index[6] & index[7] & ~index[8] & index[9] & index[11]) | (~index[0] & ~index[2] & ~index[3] & index[4] & ~index[7] & ~index[8] & ~index[10] & ~index[11]) | (index[0] & index[1] & index[2] & index[3] & ~index[4] & ~index[6] & index[7] & index[8] & ~index[11]) | (~index[0] & ~index[2] & ~index[3] & ~index[4] & ~index[5] & index[7] & index[8] & index[9] & index[10] & ~index[11]) | (index[1] & ~index[2] & index[3] & index[4] & ~index[7] & index[8] & index[9] & index[10] & ~index[11]) | (index[0] & index[1] & index[2] & index[3] & index[4] & index[6] & ~index[7] & ~index[8] & index[10]) | (index[1] & index[2] & ~index[3] & ~index[4] & ~index[5] & ~index[6] & index[8] & ~index[9] & index[11]) | (index[0] & index[1] & ~index[2] & index[5] & ~index[6] & ~index[8] & index[11]) | (index[0] & index[1] & ~index[2] & ~index[4] & ~index[6] & index[7] & ~index[8] & ~index[9] & index[11]) | (~index[0] & ~index[1] & ~index[2] & index[3] & ~index[6] & ~index[7] & ~index[8] & index[11]) | (index[1] & ~index[2] & ~index[3] & index[4] & ~index[7] & index[8] & index[9] & ~index[10]) | (index[0] & ~index[1] & ~index[2] & ~index[3] & ~index[5] & ~index[6] & ~index[7] & index[8] & index[11]) | (~index[0] & index[1] & ~index[2] & index[3] & index[4] & index[6] & ~index[8] & index[9] & ~index[10]) | (~index[0] & ~index[1] & index[2] & index[4] & index[7] & ~index[9] & index[10]) | (index[0] & index[1] & index[2] & ~index[3] & ~index[4] & ~index[6] & index[8] & index[9] & index[10] & ~index[11]) | (index[2] & ~index[3] & index[5] & index[6] & index[7] & ~index[8] & index[9]) | (~index[0] & ~index[1] & index[4] & index[6] & index[7] & ~index[8] & ~index[9] & ~index[10] & ~index[11]) | (index[0] & index[2] & ~index[3] & ~index[4] & ~index[5] & ~index[6] & index[7] & index[8] & index[10]) | (index[0] & ~index[1] & index[2] & index[5] & ~index[7] & index[8] & ~index[11]) | (~index[0] & ~index[1] & index[2] & ~index[3] & index[6] & ~index[7] & index[8] & ~index[9] & ~index[10]) | (~index[1] & ~index[2] & ~index[3] & ~index[4] & ~index[5] & index[6] & ~index[9] & index[10] & ~index[11]) | (index[2] & ~index[3] & ~index[4] & ~index[5] & index[6] & index[7] & index[10] & index[11]) | (index[0] & ~index[1] & ~index[2] & index[3] & index[4] & ~index[7] & index[10] & index[11]) | (~index[0] & ~index[1] & index[2] & ~index[3] & index[4] & ~index[6] & index[8] & index[9] & ~index[11]) | (~index[0] & index[2] & index[6] & ~index[7] & index[8] & ~index[9] & ~index[10] & ~index[11]) | (~index[0] & index[1] & ~index[2] & ~index[3] & ~index[4] & ~index[5] & index[6] & ~index[7] & index[11]) | (~index[0] & index[2] & ~index[3] & index[4] & ~index[7] & ~index[8] & ~index[9] & index[11]) | (~index[1] & index[2] & index[3] & index[4] & index[6] & ~index[8] & index[9] & index[11]) | (~index[0] & ~index[1] & ~index[2] & ~index[4] & ~index[5] & index[7] & ~index[8] & ~index[9] & index[10] & ~index[11]) | (index[0] & ~index[1] & index[2] & ~index[3] & ~index[6] & index[7] & index[10] & index[11]) | (index[0] & index[1] & index[2] & ~index[3] & index[4] & ~index[6] & ~index[8] & ~index[9]) | (index[0] & ~index[1] & index[2] & ~index[3] & ~index[4] & ~index[5] & index[6] & index[8] & index[11]) | (~index[0] & index[1] & ~index[2] & ~index[3] & index[4] & index[7] & ~index[9] & index[11]) | (index[0] & ~index[1] & ~index[2] & ~index[3] & ~index[4] & ~index[5] & index[6] & ~index[7] & ~index[8] & ~index[9]) | (~index[0] & ~index[1] & index[3] & ~index[4] & index[6] & index[7] & ~index[9] & index[11]) | (~index[2] & ~index[3] & index[4] & ~index[6] & index[7] & ~index[8] & index[9] & index[11]) | (index[0] & index[1] & ~index[2] & index[5] & index[7] & index[9] & ~index[10]) | (index[2] & index[4] & index[5] & ~index[6] & ~index[7]) | (~index[0] & ~index[1] & index[2] & index[3] & ~index[5] & index[6] & ~index[7] & index[9] & index[11]) | (~index[2] & index[3] & ~index[6] & ~index[8] & ~index[9] & ~index[10] & ~index[11]) | (index[0] & ~index[1] & ~index[2] & ~index[3] & index[4] & index[6] & index[7] & ~index[9] & index[11]) | (~index[0] & ~index[1] & index[2] & index[3] & ~index[4] & ~index[5] & index[7] & ~index[9] & ~index[10]) | (~index[0] & ~index[1] & ~index[2] & index[5] & index[6] & index[9] & index[11]) | (index[1] & index[2] & index[3] & ~index[4] & ~index[6] & index[7] & ~index[8] & index[9] & ~index[10]) | (index[0] & ~index[1] & ~index[2] & ~index[3] & index[4] & index[6] & ~index[7] & index[9] & ~index[10]) | (index[0] & index[2] & index[3] & index[4] & ~index[7] & index[8] & ~index[10] & ~index[11]) | (~index[0] & index[3] & index[4] & index[6] & index[7] & index[8] & ~index[9] & index[10]) | (~index[0] & ~index[1] & index[2] & ~index[4] & ~index[5] & index[6] & index[7] & index[8] & index[11]) | (index[2] & index[3] & ~index[4] & ~index[5] & ~index[6] & index[7] & ~index[8] & ~index[9] & index[10]) | (index[1] & ~index[3] & ~index[4] & ~index[5] & index[6] & index[7] & ~index[8] & ~index[9] & index[11]) | (index[0] & ~index[2] & index[3] & ~index[4] & index[6] & index[7] & index[8] & ~index[10]) | (index[1] & index[2] & index[4] & ~index[6] & ~index[7] & ~index[8] & ~index[9]) | (~index[0] & index[1] & ~index[2] & ~index[3] & ~index[5] & index[6] & index[10] & index[11]) | (~index[1] & ~index[2] & index[3] & ~index[4] & index[6] & ~index[7] & index[8] & ~index[9] & ~index[11]) | (index[0] & index[3] & ~index[4] & ~index[6] & index[7] & ~index[8] & ~index[9] & index[11]) | (~index[0] & index[2] & index[3] & index[4] & index[6] & ~index[7] & index[8] & index[9] & index[10]) | (~index[1] & ~index[3] & ~index[4] & index[5] & index[6] & ~index[7] & index[9] & index[11]) | (~index[0] & index[1] & ~index[2] & ~index[3] & ~index[4] & index[6] & index[8] & index[9] & index[10]) | (index[0] & ~index[1] & ~index[2] & index[3] & index[4] & ~index[6] & ~index[7] & index[9] & index[11]) | (index[0] & ~index[2] & ~index[3] & ~index[4] & ~index[5] & index[6] & ~index[7] & index[9] & ~index[11]) | (index[0] & index[1] & ~index[2] & index[3] & index[5] & index[7] & index[9]) | (~index[0] & ~index[1] & ~index[2] & index[3] & index[5] & index[6] & index[8]) | (index[1] & ~index[2] & ~index[4] & ~index[5] & index[6] & index[8] & index[9] & ~index[10]) | (index[0] & ~index[1] & index[5] & ~index[6] & ~index[8] & index[9] & index[10]) | (index[0] & ~index[1] & index[2] & index[3] & index[5] & index[8] & ~index[11]) | (index[0] & index[1] & ~index[2] & ~index[4] & ~index[5] & index[6] & ~index[8] & ~index[9] & index[11]) | (index[0] & index[1] & index[5] & ~index[6] & index[8] & index[9] & ~index[11]) | (~index[0] & index[1] & index[5] & index[6] & ~index[7] & ~index[11]) | (index[0] & ~index[1] & ~index[2] & ~index[3] & ~index[6] & index[7] & ~index[9] & index[10]) | (~index[0] & ~index[1] & ~index[2] & index[3] & ~index[4] & ~index[8] & ~index[9] & ~index[10] & ~index[11]) | (~index[0] & ~index[1] & index[2] & ~index[3] & index[5] & ~index[9] & index[11]) | (index[0] & index[1] & ~index[2] & index[3] & index[6] & index[7] & index[8] & index[9] & ~index[10]) | (~index[0] & index[1] & index[3] & index[4] & ~index[6] & ~index[7] & index[9] & ~index[11]) | (index[0] & ~index[1] & index[2] & ~index[3] & ~index[4] & ~index[6] & index[7] & ~index[9] & ~index[10] & ~index[11]) | (~index[0] & index[1] & ~index[2] & ~index[4] & ~index[6] & index[7] & index[8] & ~index[9] & ~index[11]) | (~index[0] & index[1] & ~index[2] & ~index[3] & ~index[4] & index[6] & ~index[7] & index[10]) | (~index[0] & ~index[1] & index[2] & index[3] & ~index[4] & index[6] & index[7] & ~index[8] & ~index[11]) | (index[0] & index[1] & ~index[2] & ~index[3] & ~index[6] & index[7] & index[8] & index[9] & ~index[10]) | (index[0] & ~index[1] & index[2] & ~index[3] & index[4] & ~index[6] & ~index[7] & ~index[11]) | (~index[1] & index[2] & index[3] & index[4] & ~index[6] & index[7] & index[9] & index[11]) | (~index[1] & index[3] & ~index[4] & index[6] & ~index[7] & ~index[8] & index[9] & index[10]) | (~index[0] & ~index[1] & index[3] & index[4] & index[6] & index[7] & index[8] & index[9] & ~index[11]) | (index[0] & index[1] & index[2] & index[3] & index[4] & index[6] & ~index[9] & index[11]) | (~index[1] & ~index[2] & ~index[3] & ~index[4] & index[6] & index[7] & index[8] & ~index[9] & ~index[11]) | (~index[0] & ~index[1] & ~index[3] & ~index[4] & ~index[6] & ~index[7] & ~index[9] & ~index[10] & index[11]) | (index[0] & index[1] & ~index[2] & index[3] & ~index[7] & ~index[8] & ~index[10] & ~index[11]) | (~index[0] & index[1] & ~index[2] & ~index[3] & index[4] & ~index[6] & ~index[7] & index[8]) | (index[1] & ~index[2] & ~index[4] & ~index[5] & index[6] & index[7] & index[8] & ~index[10] & ~index[11]) | (~index[1] & ~index[2] & index[5] & index[7] & ~index[9] & ~index[10] & ~index[11]) | (~index[0] & ~index[1] & ~index[2] & ~index[3] & index[5] & index[6] & ~index[8] & index[9]) | (~index[0] & index[1] & ~index[2] & ~index[5] & ~index[6] & ~index[7] & index[10] & index[11]) | (index[0] & ~index[1] & index[5] & ~index[7] & index[8] & ~index[9] & index[10]) | (~index[0] & ~index[1] & index[3] & ~index[4] & ~index[6] & index[7] & ~index[10] & ~index[11]) | (~index[0] & ~index[1] & ~index[2] & index[5] & ~index[7] & ~index[8] & index[9]) | (~index[0] & index[1] & ~index[2] & ~index[3] & index[4] & index[7] & ~index[8] & index[10]) | (index[0] & index[5] & ~index[6] & index[7] & index[9] & ~index[10]) | (index[0] & ~index[1] & index[2] & index[3] & index[4] & ~index[6] & index[7] & index[9] & index[10]) | (~index[0] & index[1] & index[2] & ~index[4] & ~index[6] & ~index[7] & index[10] & index[11]) | (~index[1] & ~index[3] & index[4] & ~index[6] & index[7] & index[8] & index[9] & ~index[10]) | (index[0] & ~index[1] & ~index[2] & index[6] & index[7] & index[8] & ~index[9] & ~index[10] & ~index[11]) | (~index[0] & index[2] & ~index[3] & ~index[4] & ~index[5] & index[6] & ~index[8] & index[9] & ~index[11]) | (index[0] & ~index[1] & ~index[3] & ~index[4] & ~index[5] & index[7] & index[9] & index[11]) | (index[0] & index[1] & index[2] & ~index[4] & index[6] & index[7] & ~index[8] & index[9] & index[10]) | (index[0] & index[1] & index[5] & index[6] & index[7] & index[8] & index[11]) | (index[0] & ~index[1] & index[2] & ~index[3] & index[5] & index[7] & ~index[8] & index[10]) | (index[0] & index[1] & index[2] & ~index[4] & ~index[5] & ~index[6] & ~index[7] & ~index[8] & index[9] & index[11]) | (index[1] & index[2] & index[3] & ~index[4] & index[6] & ~index[7] & index[8] & index[9] & index[10] & ~index[11]) | (index[0] & ~index[3] & ~index[4] & ~index[5] & ~index[6] & index[7] & index[8] & ~index[9] & ~index[11]) | (index[0] & index[1] & index[2] & ~index[4] & index[6] & ~index[8] & ~index[9] & ~index[10] & ~index[11]) | (~index[0] & ~index[1] & index[2] & ~index[3] & ~index[5] & index[6] & index[7] & index[9] & index[11]) | (index[0] & index[1] & ~index[2] & index[3] & ~index[4] & index[7] & index[11]) | (~index[0] & index[1] & ~index[3] & index[4] & index[6] & index[7] & index[8] & ~index[10] & ~index[11]) | (index[0] & ~index[2] & index[3] & ~index[4] & ~index[6] & index[7] & index[11]) | (index[0] & ~index[1] & index[2] & index[3] & ~index[4] & ~index[6] & ~index[9] & index[11]) | (index[0] & index[1] & index[2] & index[3] & ~index[4] & index[6] & ~index[9] & ~index[10] & ~index[11]) | (index[0] & index[1] & ~index[2] & index[3] & index[4] & index[6] & index[7] & index[9] & index[10] & ~index[11]) | (index[1] & index[2] & index[3] & ~index[4] & ~index[5] & ~index[6] & index[7] & index[9] & index[11]) | (index[0] & ~index[1] & ~index[2] & index[4] & index[6] & ~index[8] & index[9] & ~index[10] & ~index[11]) | (index[0] & index[1] & ~index[3] & ~index[4] & ~index[6] & ~index[8] & index[9] & ~index[10] & ~index[11]) | (index[0] & ~index[3] & ~index[4] & ~index[5] & index[6] & ~index[7] & index[8] & index[9] & ~index[10]) | (~index[0] & ~index[1] & index[2] & index[5] & index[6] & index[7] & ~index[8] & index[10]) | (~index[1] & index[2] & index[3] & ~index[4] & ~index[5] & index[6] & ~index[8] & index[9] & index[10]) | (index[0] & index[1] & index[5] & index[6] & index[7] & ~index[8] & index[9]) | (index[0] & ~index[2] & index[3] & ~index[4] & index[6] & ~index[7] & ~index[8] & index[9]) | (~index[0] & index[1] & ~index[3] & index[5] & ~index[8] & ~index[10] & ~index[11]) | (~index[2] & ~index[3] & index[4] & index[6] & index[7] & index[8] & ~index[10] & index[11]) | (~index[0] & ~index[1] & index[2] & ~index[5] & index[6] & ~index[7] & ~index[8] & index[9] & index[10]) | (index[0] & ~index[2] & ~index[3] & ~index[5] & ~index[6] & ~index[7] & ~index[9] & ~index[10] & ~index[11]) | (index[0] & ~index[1] & ~index[2] & ~index[3] & index[7] & index[8] & ~index[10] & index[11]) | (~index[0] & ~index[2] & ~index[3] & index[4] & index[5] & ~index[6]) | (~index[0] & ~index[1] & index[2] & index[3] & ~index[6] & ~index[9] & ~index[10] & ~index[11]) | (~index[0] & index[1] & ~index[2] & ~index[3] & ~index[4] & ~index[5] & index[10] & index[11]) | (~index[0] & index[1] & ~index[2] & ~index[3] & ~index[4] & ~index[5] & ~index[7] & ~index[8] & index[9]) | (index[0] & index[1] & ~index[2] & index[3] & ~index[4] & ~index[6] & ~index[8] & index[9] & index[10]) | (~index[0] & ~index[1] & index[2] & ~index[3] & index[4] & index[8] & ~index[9] & index[10]) | (index[0] & index[1] & index[3] & ~index[4] & ~index[6] & ~index[7] & ~index[8] & index[9]) | (index[0] & ~index[1] & ~index[2] & index[3] & index[4] & ~index[6] & ~index[7] & index[8] & index[9]) | (~index[1] & ~index[2] & index[3] & ~index[4] & ~index[5] & index[6] & index[7] & index[8] & index[9] & index[10] & ~index[11]) | (index[0] & ~index[2] & index[3] & ~index[4] & ~index[7] & index[8] & ~index[9] & index[10]) | (~index[0] & ~index[2] & ~index[3] & ~index[4] & ~index[5] & index[6] & index[7] & ~index[8] & ~index[9] & ~index[10] & index[11]) | (~index[0] & ~index[1] & ~index[3] & ~index[4] & ~index[6] & ~index[7] & ~index[8] & index[10] & ~index[11]) | (index[1] & ~index[3] & index[4] & ~index[6] & index[7] & ~index[8] & ~index[9] & ~index[10]) | (~index[1] & index[2] & ~index[3] & index[4] & index[7] & ~index[9] & index[10]) | (~index[0] & ~index[1] & index[2] & ~index[4] & index[6] & index[7] & index[8] & ~index[9]) | (~index[1] & index[3] & index[4] & index[6] & index[7] & index[8] & ~index[9] & index[10]) | (index[0] & index[2] & ~index[3] & index[4] & index[6] & index[7] & index[8] & index[9] & ~index[10]) | (index[0] & index[2] & index[5] & ~index[6] & index[9] & ~index[11]) | (index[0] & index[2] & ~index[3] & index[4] & ~index[6] & index[7] & ~index[8] & ~index[9] & index[11]) | (index[1] & index[2] & ~index[3] & index[4] & index[6] & ~index[7] & index[9] & index[11]) | (index[0] & index[1] & index[2] & index[3] & index[4] & index[7] & index[8] & ~index[9]) | (index[0] & ~index[1] & index[2] & index[4] & ~index[7] & ~index[9] & ~index[10] & ~index[11]) | (index[0] & ~index[1] & ~index[2] & ~index[4] & ~index[6] & index[7] & index[8] & ~index[9] & index[10]) | (~index[0] & index[2] & ~index[3] & index[4] & ~index[6] & ~index[7] & ~index[8] & index[11]);

assign val[3] = (index[0] & index[2] & index[3] & ~index[4] & ~index[5] & index[6] & ~index[7] & index[10] & index[11]) | (~index[0] & index[2] & index[3] & index[4] & ~index[6] & ~index[7] & ~index[8] & index[11]) | (~index[0] & ~index[2] & index[3] & index[4] & ~index[6] & ~index[7] & ~index[8] & index[9] & index[10]) | (~index[0] & ~index[1] & ~index[2] & ~index[3] & index[4] & index[7] & index[8] & ~index[9] & index[10]) | (index[0] & ~index[1] & index[3] & ~index[4] & ~index[6] & index[7] & index[8] & ~index[9] & index[11]) | (~index[0] & ~index[1] & ~index[2] & ~index[3] & index[4] & ~index[6] & ~index[7] & ~index[8] & ~index[9] & index[11]) | (~index[0] & ~index[1] & index[3] & index[6] & ~index[7] & index[8] & ~index[9] & index[10]) | (index[0] & index[5] & index[7] & ~index[8] & index[9] & index[11]) | (index[0] & index[1] & index[2] & index[5] & index[7] & ~index[8] & index[9]) | (index[0] & index[1] & ~index[2] & index[3] & ~index[4] & index[6] & ~index[8] & index[9] & index[10]) | (index[0] & index[1] & index[2] & ~index[3] & index[4] & ~index[6] & ~index[7] & index[8] & index[9] & index[10] & ~index[11]) | (index[0] & index[1] & ~index[2] & index[4] & index[6] & ~index[7] & index[8] & index[9] & ~index[10]) | (~index[1] & ~index[2] & ~index[3] & ~index[4] & ~index[5] & index[6] & ~index[7] & index[8] & index[10] & ~index[11]) | (index[0] & ~index[1] & index[2] & ~index[3] & ~index[4] & ~index[5] & ~index[6] & ~index[7] & index[8] & index[11]) | (~index[0] & ~index[1] & ~index[2] & ~index[3] & ~index[4] & ~index[5] & index[6] & index[7] & ~index[9] & ~index[10] & index[11]) | (index[0] & index[1] & ~index[2] & ~index[3] & ~index[6] & ~index[7] & ~index[9] & ~index[10] & ~index[11]) | (~index[1] & ~index[2] & index[3] & index[4] & ~index[6] & ~index[7] & index[10] & index[11]) | (index[0] & index[1] & ~index[3] & index[4] & index[6] & ~index[7] & ~index[8] & ~index[9] & index[11]) | (index[0] & index[1] & index[2] & ~index[4] & ~index[5] & ~index[6] & index[7] & ~index[8] & ~index[9] & index[10]) | (~index[0] & index[1] & ~index[3] & ~index[4] & ~index[5] & index[6] & ~index[7] & index[9] & index[11]) | (index[0] & index[1] & ~index[2] & index[3] & ~index[4] & index[9] & ~index[10] & index[11]) | (index[1] & ~index[2] & index[3] & ~index[4] & ~index[5] & ~index[6] & ~index[7] & index[8] & index[11]) | (index[0] & index[2] & index[3] & index[6] & ~index[7] & ~index[8] & ~index[9] & index[10]) | (~index[0] & ~index[1] & index[2] & ~index[3] & ~index[4] & index[5] & ~index[6] & index[7] & index[11]) | (~index[1] & index[2] & ~index[3] & index[4] & ~index[6] & index[7] & index[8] & index[9] & ~index[10]) | (index[0] & index[1] & ~index[3] & index[4] & ~index[6] & ~index[7] & index[9] & ~index[10] & index[11]) | (index[0] & index[1] & ~index[2] & index[3] & index[4] & index[6] & index[7] & ~index[8]) | (~index[0] & index[1] & index[2] & index[4] & index[6] & ~index[7] & index[8] & index[9] & index[10]) | (~index[0] & index[1] & index[2] & index[3] & ~index[6] & ~index[7] & ~index[8] & ~index[9]) | (index[0] & ~index[1] & index[2] & index[3] & ~index[4] & ~index[6] & index[7] & index[8] & ~index[9] & ~index[10]) | (index[0] & index[1] & ~index[2] & ~index[4] & ~index[5] & index[6] & index[7] & ~index[8] & index[11]) | (index[0] & ~index[1] & ~index[2] & ~index[3] & index[4] & ~index[7] & index[8] & ~index[9] & index[11]) | (index[0] & index[1] & ~index[2] & index[3] & ~index[6] & index[7] & index[10] & index[11]) | (index[0] & ~index[1] & index[2] & index[3] & ~index[4] & index[6] & ~index[7] & index[8] & ~index[10]) | (index[0] & ~index[1] & ~index[3] & index[6] & index[7] & ~index[8] & index[9] & index[10]) | (~index[0] & index[1] & index[2] & index[4] & index[7] & ~index[8] & ~index[9] & index[10]) | (~index[0] & ~index[2] & index[3] & index[5] & index[7] & ~index[9] & ~index[10]) | (index[0] & index[1] & ~index[3] & index[6] & index[7] & index[8] & ~index[9] & index[10]) | (index[0] & index[1] & ~index[2] & ~index[3] & index[4] & ~index[6] & ~index[8] & index[9] & index[10]) | (index[0] & index[2] & ~index[3] & index[4] & ~index[7] & ~index[8] & ~index[9] & index[10]) | (index[0] & ~index[1] & index[2] & ~index[3] & ~index[4] & ~index[5] & index[7] & index[8] & index[9] & ~index[10]) | (index[0] & ~index[1] & index[3] & ~index[6] & ~index[7] & index[8] & index[9] & ~index[10]) | (index[0] & index[1] & ~index[2] & ~index[3] & index[4] & ~index[6] & index[7] & index[8] & index[9] & ~index[11]) | (index[0] & index[1] & index[2] & ~index[3] & index[4] & index[6] & ~index[7] & ~index[8] & index[9]) | (index[0] & index[1] & index[2] & ~index[3] & index[4] & index[6] & index[7] & index[8] & ~index[10] & ~index[11]) | (index[0] & index[1] & ~index[4] & ~index[7] & ~index[8] & ~index[10] & ~index[11]) | (index[0] & index[1] & index[2] & index[3] & ~index[6] & ~index[7] & ~index[8] & index[9]) | (~index[0] & ~index[1] & index[2] & index[6] & index[7] & index[8] & ~index[9] & index[10]) | (index[0] & index[3] & index[4] & index[6] & index[7] & ~index[8] & index[9]) | (~index[0] & ~index[1] & index[2] & ~index[3] & ~index[6] & ~index[7] & index[8] & ~index[9] & index[10]) | (~index[1] & index[2] & ~index[3] & index[5] & ~index[8] & ~index[9] & index[10]) | (index[0] & index[1] & index[2] & index[3] & index[6] & ~index[8] & index[9] & ~index[10]) | (index[1] & index[3] & index[4] & index[6] & ~index[7] & index[8] & ~index[10] & index[11]) | (index[0] & index[1] & index[5] & ~index[7] & ~index[8] & ~index[9] & index[10]) | (~index[0] & ~index[1] & index[2] & ~index[3] & ~index[4] & index[6] & ~index[8] & ~index[9] & index[10]) | (~index[0] & index[1] & ~index[2] & index[3] & index[4] & ~index[6] & index[8] & index[9] & ~index[10]) | (index[0] & ~index[1] & index[2] & ~index[3] & ~index[4] & ~index[6] & index[7] & index[9] & ~index[10] & index[11]) | (index[0] & index[1] & ~index[2] & index[3] & index[4] & index[7] & index[8] & index[11]) | (index[0] & ~index[2] & index[4] & ~index[6] & ~index[7] & ~index[9] & ~index[10] & ~index[11]) | (~index[0] & ~index[1] & index[2] & ~index[3] & index[6] & ~index[8] & index[9] & ~index[10] & ~index[11]) | (index[0] & ~index[2] & ~index[3] & ~index[4] & ~index[6] & ~index[8] & ~index[9] & index[11]) | (~index[0] & ~index[1] & ~index[3] & ~index[4] & ~index[5] & index[6] & ~index[7] & index[9] & index[10] & ~index[11]) | (index[0] & ~index[1] & ~index[2] & index[3] & index[4] & index[7] & index[8] & index[10] & ~index[11]) | (~index[0] & ~index[1] & ~index[2] & ~index[3] & index[4] & index[7] & index[8] & index[9] & ~index[10]) | (~index[0] & index[1] & index[2] & index[4] & ~index[6] & index[8] & ~index[9] & ~index[10]) | (~index[0] & ~index[1] & index[2] & ~index[3] & ~index[5] & ~index[7] & ~index[8] & index[9] & index[10]) | (index[0] & ~index[2] & index[3] & index[4] & index[7] & ~index[8] & index[9] & index[10]) | (index[0] & index[1] & index[3] & ~index[4] & ~index[6] & ~index[7] & index[8] & ~index[10] & index[11]) | (~index[0] & ~index[1] & ~index[2] & ~index[3] & index[4] & ~index[7] & ~index[9] & ~index[10] & ~index[11]) | (~index[0] & index[1] & index[2] & index[4] & index[6] & index[7] & ~index[10] & index[11]) | (index[0] & index[1] & ~index[2] & index[3] & index[6] & index[7] & ~index[10] & index[11]) | (~index[0] & ~index[1] & index[2] & ~index[4] & ~index[5] & index[6] & index[7] & ~index[8] & ~index[9] & index[11]) | (~index[0] & index[2] & index[3] & ~index[4] & ~index[5] & index[6] & index[7] & index[8] & index[9] & ~index[10]) | (~index[0] & index[1] & index[2] & index[3] & ~index[7] & ~index[9] & ~index[10] & ~index[11]) | (~index[0] & ~index[1] & index[2] & ~index[3] & ~index[4] & ~index[5] & ~index[6] & index[7] & ~index[8] & index[10]) | (~index[0] & index[1] & index[3] & index[4] & ~index[6] & index[7] & ~index[8] & ~index[9] & index[10]) | (~index[0] & index[1] & ~index[2] & index[3] & ~index[5] & index[6] & ~index[7] & ~index[8] & ~index[9] & ~index[10]) | (index[0] & ~index[1] & index[2] & ~index[3] & index[4] & ~index[6] & ~index[7] & index[8] & ~index[10]) | (index[0] & ~index[1] & ~index[2] & ~index[3] & ~index[4] & index[7] & index[8] & ~index[9] & ~index[10] & ~index[11]) | (~index[0] & index[1] & index[2] & ~index[5] & ~index[6] & ~index[7] & ~index[8] & ~index[9] & index[10]) | (index[1] & index[2] & ~index[3] & index[4] & ~index[6] & ~index[8] & ~index[10] & ~index[11]) | (index[0] & ~index[1] & ~index[3] & ~index[4] & ~index[5] & ~index[6] & index[8] & ~index[9] & index[10]) | (~index[0] & ~index[1] & index[2] & ~index[4] & index[6] & ~index[7] & index[8] & ~index[9] & ~index[10] & ~index[11]) | (~index[0] & index[1] & index[2] & ~index[3] & ~index[4] & ~index[5] & index[6] & ~index[8] & index[9] & index[10]) | (~index[0] & ~index[1] & index[5] & index[6] & index[8] & ~index[9]) | (~index[0] & ~index[1] & index[3] & ~index[4] & index[6] & ~index[7] & index[8] & ~index[9]) | (index[0] & index[1] & ~index[2] & index[3] & index[4] & ~index[7] & index[8] & index[9] & index[10] & ~index[11]) | (~index[0] & ~index[1] & ~index[2] & ~index[3] & index[5] & ~index[6] & index[7] & index[8] & index[9]) | (~index[0] & index[1] & ~index[2] & ~index[6] & ~index[8] & ~index[9] & ~index[10] & ~index[11]) | (index[0] & ~index[1] & ~index[2] & ~index[3] & ~index[4] & ~index[7] & index[8] & index[9] & index[10] & ~index[11]) | (~index[0] & index[1] & index[5] & index[6] & index[8] & ~index[10] & ~index[11]) | (index[0] & ~index[2] & ~index[4] & index[6] & index[7] & index[9] & ~index[10] & index[11]) | (index[0] & ~index[2] & index[3] & ~index[4] & ~index[5] & index[7] & index[8] & index[9] & ~index[10]) | (~index[0] & ~index[1] & index[2] & index[3] & ~index[4] & ~index[5] & ~index[6] & index[7] & index[9] & index[11]) | (~index[0] & index[1] & ~index[2] & ~index[3] & ~index[4] & ~index[5] & ~index[6] & index[8] & ~index[9] & index[10]) | (~index[0] & ~index[1] & index[2] & ~index[3] & ~index[6] & ~index[8] & ~index[9] & ~index[10] & ~index[11]) | (index[1] & ~index[2] & index[3] & index[5] & ~index[6] & index[7] & ~index[9]) | (index[0] & index[1] & ~index[3] & ~index[4] & ~index[5] & ~index[6] & index[7] & ~index[8] & index[9] & ~index[11]) | (index[0] & index[1] & ~index[3] & ~index[4] & index[6] & index[8] & ~index[9] & index[10]) | (~index[0] & index[1] & ~index[2] & ~index[3] & ~index[4] & ~index[5] & ~index[6] & ~index[7] & ~index[8] & index[9]) | (~index[0] & index[1] & ~index[3] & ~index[4] & ~index[5] & ~index[6] & index[7] & ~index[8] & ~index[9] & index[11]) | (~index[0] & index[1] & ~index[2] & ~index[3] & ~index[4] & ~index[5] & ~index[6] & index[7] & ~index[9]) | (~index[0] & ~index[2] & ~index[3] & ~index[4] & index[6] & index[7] & index[8] & index[9] & index[10] & ~index[11]) | (~index[0] & ~index[1] & ~index[2] & index[3] & index[4] & index[6] & ~index[7] & index[8] & index[9] & ~index[10]) | (index[0] & ~index[1] & index[2] & index[3] & index[4] & ~index[7] & ~index[9] & index[11]) | (index[0] & ~index[1] & index[2] & ~index[3] & index[4] & ~index[5] & index[6] & index[10] & index[11]) | (index[1] & ~index[2] & index[3] & ~index[4] & index[6] & index[7] & index[8] & ~index[9] & ~index[11]) | (~index[1] & index[2] & index[3] & index[5] & ~index[8] & index[9]) | (index[2] & index[3] & index[4] & ~index[6] & index[7] & ~index[8] & ~index[9] & index[10]) | (index[0] & ~index[2] & index[3] & index[5] & index[7] & index[8] & index[10]) | (~index[0] & index[2] & index[3] & index[4] & index[6] & ~index[7] & index[10] & index[11]) | (index[0] & ~index[1] & index[2] & index[3] & index[4] & index[7] & ~index[8] & index[11]) | (~index[0] & ~index[1] & index[2] & index[5] & index[6] & ~index[7] & index[9] & index[11]) | (index[0] & index[1] & index[3] & index[4] & index[6] & index[8] & ~index[9] & index[11]) | (~index[0] & index[1] & ~index[2] & ~index[3] & index[4] & index[7] & index[11]) | (index[0] & ~index[1] & ~index[2] & index[3] & ~index[6] & ~index[7] & ~index[10] & ~index[11]) | (~index[0] & ~index[1] & index[2] & index[3] & index[4] & ~index[6] & index[9] & ~index[10] & ~index[11]) | (~index[0] & index[1] & ~index[3] & ~index[4] & ~index[5] & index[6] & index[10] & index[11]) | (index[0] & ~index[1] & ~index[2] & index[4] & ~index[5] & index[6] & index[7] & index[9] & index[10] & ~index[11]) | (index[0] & ~index[1] & index[2] & ~index[3] & index[4] & ~index[5] & index[7] & index[10] & index[11]) | (index[0] & index[1] & index[3] & index[5] & index[7] & index[11]) | (~index[0] & index[1] & ~index[2] & ~index[3] & index[7] & index[8] & index[9] & index[10] & ~index[11]) | (index[0] & index[1] & ~index[2] & index[3] & index[4] & index[7] & ~index[9] & index[11]) | (index[0] & index[1] & index[2] & ~index[3] & ~index[5] & index[6] & index[7] & ~index[8] & ~index[9] & ~index[10] & ~index[11]) | (index[0] & ~index[1] & ~index[2] & index[3] & ~index[4] & ~index[5] & index[6] & ~index[7] & ~index[8] & ~index[9] & index[11]) | (index[0] & index[1] & index[2] & ~index[3] & ~index[4] & ~index[5] & ~index[6] & ~index[7] & index[9] & ~index[10]) | (~index[0] & ~index[2] & ~index[3] & index[5] & index[6] & ~index[7] & ~index[9] & index[11]) | (~index[0] & ~index[1] & ~index[2] & index[3] & ~index[4] & ~index[5] & index[7] & ~index[8] & ~index[9] & ~index[11]) | (~index[0] & index[1] & index[2] & ~index[5] & index[6] & ~index[7] & index[10] & index[11]) | (~index[0] & ~index[1] & index[2] & index[4] & ~index[6] & ~index[7] & index[9] & index[10] & ~index[11]) | (~index[1] & ~index[2] & index[3] & ~index[4] & ~index[5] & index[6] & ~index[7] & index[10] & index[11]) | (index[0] & ~index[1] & ~index[2] & ~index[3] & ~index[4] & ~index[6] & index[7] & index[8] & index[10]) | (index[0] & ~index[1] & ~index[2] & ~index[3] & ~index[4] & ~index[5] & ~index[6] & ~index[7] & ~index[10] & index[11]) | (index[0] & ~index[1] & index[2] & index[3] & index[4] & ~index[6] & ~index[7] & ~index[9] & index[10]) | (~index[0] & ~index[1] & ~index[2] & index[4] & index[6] & index[7] & index[8] & ~index[10] & index[11]) | (index[0] & index[1] & index[2] & index[3] & index[4] & ~index[8] & ~index[10] & ~index[11]) | (index[1] & index[2] & index[4] & index[5] & ~index[7]) | (index[0] & ~index[1] & index[2] & ~index[3] & ~index[6] & index[7] & index[8] & ~index[9] & index[10]) | (~index[0] & index[1] & index[2] & index[4] & ~index[5] & ~index[6] & index[7] & index[8] & index[11]) | (index[0] & ~index[1] & index[2] & index[5] & index[8] & index[9] & index[10] & ~index[11]) | (~index[0] & index[1] & index[2] & index[3] & ~index[4] & ~index[6] & ~index[8] & index[9] & ~index[10] & ~index[11]) | (index[0] & ~index[1] & ~index[3] & index[4] & ~index[6] & ~index[7] & ~index[8] & ~index[9] & index[10]) | (~index[0] & ~index[2] & index[3] & ~index[4] & ~index[6] & index[7] & index[8] & ~index[9] & index[10]) | (index[0] & ~index[1] & ~index[2] & index[3] & index[4] & ~index[7] & index[10] & index[11]) | (~index[0] & index[1] & ~index[2] & ~index[3] & ~index[4] & ~index[5] & index[8] & ~index[10] & index[11]) | (index[0] & index[1] & ~index[2] & index[3] & ~index[4] & ~index[5] & index[7] & index[8] & ~index[10] & ~index[11]) | (index[0] & index[1] & ~index[2] & index[5] & index[8] & index[9] & index[10] & ~index[11]) | (index[1] & ~index[2] & ~index[3] & index[4] & ~index[6] & index[7] & ~index[8] & ~index[9] & ~index[10]) | (index[0] & ~index[1] & ~index[2] & ~index[3] & ~index[4] & ~index[5] & index[7] & index[8] & index[9] & index[10]) | (index[0] & ~index[2] & ~index[3] & ~index[6] & index[7] & index[8] & index[9] & index[10] & ~index[11]) | (index[0] & ~index[1] & ~index[3] & index[4] & index[6] & index[7] & ~index[9] & ~index[10] & ~index[11]) | (index[0] & ~index[2] & index[3] & index[4] & index[6] & index[7] & ~index[8] & index[10]) | (index[0] & ~index[1] & ~index[2] & ~index[3] & index[4] & index[6] & ~index[8] & index[9] & index[10]) | (~index[0] & index[1] & ~index[2] & ~index[3] & index[4] & ~index[7] & index[9] & ~index[10]) | (~index[0] & ~index[2] & index[3] & ~index[4] & ~index[6] & ~index[7] & index[9] & ~index[10] & index[11]) | (~index[0] & index[1] & ~index[2] & ~index[3] & ~index[4] & index[5] & ~index[7] & index[8] & index[11]) | (index[0] & ~index[1] & ~index[2] & ~index[3] & ~index[4] & index[6] & ~index[7] & index[8] & index[10]) | (~index[0] & index[1] & index[5] & index[6] & ~index[7] & index[8] & ~index[11]) | (~index[0] & ~index[1] & index[2] & index[3] & index[4] & index[7] & index[8] & index[9] & ~index[10]) | (~index[0] & ~index[1] & index[2] & ~index[3] & ~index[4] & index[7] & ~index[9] & index[10]) | (~index[0] & ~index[2] & ~index[3] & ~index[5] & ~index[6] & index[7] & ~index[8] & index[9] & ~index[10] & index[11]) | (~index[0] & ~index[1] & index[2] & index[4] & index[7] & ~index[8] & ~index[9] & ~index[10] & ~index[11]) | (~index[0] & ~index[1] & ~index[2] & ~index[3] & ~index[4] & index[5] & index[7] & index[9] & ~index[11]) | (~index[0] & index[1] & ~index[2] & ~index[3] & ~index[4] & ~index[5] & index[6] & index[7] & index[9] & index[10]) | (index[0] & index[1] & ~index[2] & index[3] & ~index[6] & ~index[7] & ~index[9] & index[11]) | (index[0] & ~index[1] & index[2] & index[5] & ~index[6] & index[7] & ~index[9] & index[10]) | (~index[0] & ~index[1] & ~index[2] & index[3] & index[4] & ~index[7] & index[8] & ~index[9] & index[10]) | (index[0] & ~index[2] & ~index[3] & ~index[4] & ~index[6] & ~index[8] & index[9] & ~index[10] & ~index[11]) | (~index[0] & ~index[1] & index[2] & index[3] & index[6] & index[7] & ~index[9] & index[11]) | (~index[0] & ~index[1] & ~index[2] & ~index[3] & index[4] & ~index[5] & index[6] & ~index[7] & index[10] & index[11]) | (~index[0] & ~index[1] & ~index[3] & index[5] & ~index[6] & ~index[7] & ~index[9] & ~index[11]) | (~index[0] & index[1] & ~index[2] & index[5] & ~index[7] & index[8] & ~index[9]) | (~index[0] & index[2] & index[4] & index[5] & ~index[7]) | (~index[0] & index[1] & ~index[2] & index[3] & ~index[4] & index[6] & ~index[7] & index[8] & index[9] & ~index[11]) | (~index[0] & index[1] & ~index[2] & index[4] & index[7] & index[9] & ~index[10] & index[11]) | (index[0] & index[1] & ~index[2] & index[3] & index[4] & ~index[6] & index[7] & index[8] & index[10]) | (index[0] & ~index[1] & index[2] & ~index[3] & index[4] & ~index[8] & ~index[9] & index[10]) | (index[0] & ~index[1] & ~index[2] & index[3] & ~index[4] & ~index[6] & index[9] & ~index[10] & ~index[11]) | (index[0] & ~index[1] & ~index[2] & index[5] & ~index[7] & index[9] & ~index[11]) | (index[0] & ~index[1] & ~index[2] & index[5] & index[6] & index[7] & ~index[8] & ~index[9]) | (~index[0] & ~index[1] & ~index[2] & ~index[3] & index[4] & index[6] & index[7] & ~index[8] & index[10]) | (~index[0] & index[1] & index[2] & ~index[3] & ~index[5] & ~index[6] & ~index[7] & index[8] & ~index[9] & ~index[10]) | (~index[0] & index[1] & ~index[2] & ~index[3] & index[4] & index[6] & index[7] & index[8] & index[10]) | (index[0] & ~index[1] & index[2] & index[4] & index[6] & index[7] & index[10] & index[11]) | (index[0] & index[1] & ~index[2] & ~index[3] & ~index[4] & ~index[8] & index[9] & ~index[10] & ~index[11]) | (index[0] & ~index[1] & ~index[2] & index[3] & index[4] & ~index[6] & ~index[7] & index[9] & index[11]) | (~index[0] & ~index[1] & index[2] & ~index[3] & index[4] & index[6] & ~index[7] & ~index[10] & index[11]) | (index[0] & ~index[1] & index[2] & index[4] & index[6] & index[8] & ~index[9] & ~index[10] & ~index[11]) | (index[0] & ~index[1] & ~index[2] & ~index[4] & index[6] & index[7] & ~index[8] & ~index[9] & index[10]) | (index[0] & index[1] & index[4] & ~index[6] & index[7] & ~index[9] & ~index[10] & ~index[11]) | (index[0] & ~index[2] & ~index[3] & ~index[4] & ~index[7] & ~index[8] & ~index[10] & ~index[11]) | (index[0] & index[1] & index[2] & index[3] & ~index[5] & ~index[6] & index[7] & ~index[8] & ~index[9] & ~index[11]) | (index[0] & index[1] & ~index[2] & index[3] & index[4] & ~index[6] & ~index[7] & ~index[8] & ~index[9]) | (index[0] & ~index[1] & index[2] & index[3] & index[4] & index[6] & ~index[7] & ~index[8] & ~index[11]) | (index[0] & index[1] & ~index[2] & ~index[4] & index[6] & index[8] & ~index[9] & index[10]) | (index[1] & index[2] & index[3] & index[6] & index[7] & index[9] & ~index[10] & index[11]) | (index[0] & index[2] & index[5] & ~index[6] & index[8] & ~index[10]) | (index[0] & index[1] & index[2] & ~index[3] & ~index[4] & ~index[5] & ~index[6] & index[7] & index[8] & index[11]) | (~index[0] & ~index[1] & index[2] & index[4] & index[6] & ~index[8] & index[9] & index[11]) | (~index[1] & ~index[2] & index[3] & ~index[4] & ~index[6] & index[7] & index[8] & index[9] & ~index[10]) | (~index[0] & index[2] & ~index[3] & ~index[4] & ~index[5] & ~index[7] & index[8] & index[9] & index[10] & ~index[11]) | (index[0] & index[1] & index[2] & ~index[3] & ~index[4] & index[6] & index[7] & ~index[9] & index[10]) | (index[0] & ~index[1] & ~index[2] & index[4] & index[5] & ~index[6] & ~index[7]) | (~index[0] & index[1] & ~index[2] & ~index[3] & index[4] & ~index[5] & ~index[6] & index[9] & index[11]) | (index[0] & ~index[1] & ~index[3] & index[5] & index[7] & ~index[9] & ~index[11]) | (index[0] & ~index[1] & index[2] & index[5] & ~index[7] & ~index[9] & index[11]) | (index[0] & ~index[1] & ~index[2] & ~index[3] & index[4] & index[6] & ~index[8] & index[9] & index[11]) | (index[1] & index[2] & index[3] & index[4] & ~index[7] & ~index[9] & ~index[10] & ~index[11]) | (~index[0] & index[2] & ~index[3] & ~index[4] & ~index[6] & index[7] & ~index[8] & ~index[9] & index[10]) | (~index[1] & ~index[2] & index[5] & index[7] & ~index[9] & ~index[10] & ~index[11]) | (~index[1] & index[2] & index[3] & ~index[4] & ~index[5] & ~index[6] & index[7] & index[10] & index[11]) | (~index[0] & ~index[1] & index[3] & index[4] & ~index[6] & index[7] & index[8] & index[11]) | (~index[0] & ~index[1] & ~index[2] & index[5] & ~index[6] & ~index[7] & ~index[8] & index[11]) | (index[0] & ~index[1] & index[2] & ~index[3] & ~index[4] & ~index[5] & index[8] & ~index[9] & index[11]) | (~index[1] & index[2] & ~index[3] & index[5] & index[7] & index[8] & index[10] & ~index[11]) | (index[0] & index[1] & index[2] & ~index[4] & ~index[6] & ~index[7] & index[8] & ~index[9] & index[10]) | (index[0] & index[1] & ~index[2] & ~index[4] & ~index[5] & index[6] & index[7] & index[8] & ~index[9] & ~index[11]) | (index[0] & index[2] & index[3] & ~index[6] & index[7] & index[8] & index[9] & index[10] & ~index[11]) | (index[0] & index[1] & ~index[2] & index[4] & ~index[6] & ~index[7] & index[8] & ~index[9] & ~index[10]) | (~index[0] & ~index[1] & index[2] & index[5] & index[8] & ~index[9]) | (~index[0] & ~index[1] & ~index[3] & ~index[4] & ~index[6] & index[7] & ~index[8] & ~index[9] & index[10] & ~index[11]) | (index[0] & ~index[1] & ~index[2] & ~index[4] & ~index[5] & index[6] & ~index[7] & index[8] & index[9] & index[10]) | (~index[0] & ~index[1] & index[3] & index[4] & ~index[6] & index[7] & index[8] & ~index[9] & ~index[10]) | (index[0] & index[1] & ~index[2] & index[3] & index[5] & index[6] & index[9] & index[10]) | (index[0] & index[5] & index[6] & index[9] & ~index[10] & index[11]) | (~index[0] & ~index[1] & ~index[2] & ~index[3] & ~index[5] & ~index[6] & ~index[7] & index[8] & index[9] & ~index[11]) | (index[0] & index[2] & index[3] & ~index[5] & ~index[6] & index[7] & ~index[8] & ~index[9] & index[10]) | (~index[0] & index[1] & ~index[2] & ~index[3] & index[4] & index[6] & ~index[7] & ~index[9] & ~index[11]) | (~index[0] & index[1] & index[2] & index[3] & index[4] & ~index[6] & index[8] & ~index[9]) | (index[0] & index[1] & ~index[2] & index[3] & index[6] & ~index[7] & index[8] & index[9] & ~index[10]) | (index[1] & index[2] & index[4] & index[6] & ~index[7] & index[8] & ~index[9] & ~index[10]) | (~index[0] & ~index[1] & index[2] & index[3] & ~index[4] & index[6] & index[7] & ~index[8] & index[9] & index[10]) | (~index[0] & ~index[1] & index[2] & index[3] & ~index[4] & ~index[7] & index[8] & ~index[9] & ~index[10]) | (index[1] & ~index[2] & index[3] & ~index[4] & ~index[5] & index[6] & index[7] & ~index[8] & index[9] & index[10]) | (~index[0] & index[1] & index[2] & index[3] & index[4] & ~index[6] & index[7] & index[10]) | (~index[0] & index[1] & ~index[2] & index[4] & index[6] & ~index[7] & index[8] & ~index[9] & ~index[11]) | (~index[0] & index[1] & index[2] & index[3] & index[5] & ~index[6]) | (~index[1] & index[3] & ~index[4] & ~index[5] & index[6] & index[7] & ~index[8] & ~index[9] & index[10]) | (index[0] & ~index[1] & index[2] & index[3] & ~index[6] & ~index[8] & ~index[9] & index[11]) | (index[0] & index[1] & index[3] & ~index[4] & ~index[6] & index[7] & index[8] & index[9] & ~index[11]) | (~index[0] & ~index[1] & ~index[2] & index[3] & ~index[4] & index[6] & ~index[8] & ~index[10] & ~index[11]) | (index[0] & index[1] & index[2] & ~index[3] & ~index[4] & ~index[6] & index[7] & index[8] & ~index[9] & ~index[10]) | (~index[0] & ~index[1] & index[2] & ~index[3] & ~index[4] & ~index[5] & ~index[6] & ~index[7] & ~index[8] & index[9]) | (~index[1] & ~index[2] & index[3] & index[4] & index[6] & index[7] & ~index[8] & index[9] & ~index[10]) | (~index[0] & index[1] & index[2] & index[3] & ~index[4] & index[6] & index[7] & index[8] & index[9] & ~index[11]) | (~index[1] & index[2] & index[3] & ~index[4] & index[6] & ~index[7] & index[8] & ~index[9]) | (~index[0] & ~index[2] & index[3] & index[4] & index[6] & ~index[7] & ~index[8] & ~index[9] & index[11]) | (index[1] & index[2] & index[3] & ~index[4] & ~index[6] & ~index[7] & ~index[8] & index[10]) | (~index[0] & index[1] & index[4] & index[5] & index[6]) | (~index[0] & index[1] & ~index[3] & index[4] & index[6] & ~index[7] & index[8] & ~index[10] & ~index[11]) | (~index[0] & index[1] & index[2] & index[3] & index[4] & index[7] & index[8] & index[11]) | (index[0] & index[1] & index[2] & index[4] & ~index[7] & ~index[8] & index[11]) | (~index[0] & index[1] & ~index[3] & index[4] & ~index[6] & index[7] & ~index[8] & index[9]) | (index[0] & ~index[1] & ~index[2] & index[3] & ~index[4] & ~index[7] & ~index[8] & index[10]) | (index[0] & ~index[1] & ~index[2] & ~index[4] & ~index[6] & index[7] & index[8] & ~index[9] & index[10]) | (index[0] & ~index[2] & ~index[3] & ~index[4] & ~index[5] & ~index[6] & ~index[7] & ~index[8] & ~index[9]);

assign val[4] = (index[0] & index[1] & index[3] & index[4] & ~index[6] & ~index[7] & ~index[9] & index[11]) | (~index[0] & index[1] & ~index[2] & ~index[3] & ~index[4] & ~index[5] & index[7] & ~index[8] & index[9] & index[11]) | (index[0] & ~index[1] & ~index[2] & ~index[3] & ~index[6] & index[7] & index[8] & ~index[10] & index[11]) | (~index[0] & index[1] & index[3] & index[4] & ~index[6] & index[7] & index[8] & index[9] & ~index[10]) | (index[0] & ~index[1] & index[2] & index[3] & ~index[4] & ~index[8] & ~index[9] & ~index[10] & ~index[11]) | (index[0] & ~index[1] & ~index[2] & ~index[3] & ~index[4] & ~index[5] & index[6] & index[9] & ~index[10] & ~index[11]) | (~index[0] & ~index[2] & ~index[3] & index[4] & ~index[6] & ~index[7] & index[8] & ~index[9] & index[11]) | (index[0] & ~index[1] & index[2] & ~index[3] & ~index[4] & ~index[5] & ~index[6] & index[7] & ~index[8] & ~index[9]) | (~index[0] & ~index[1] & index[2] & index[3] & index[4] & ~index[6] & index[8] & ~index[9] & index[10]) | (~index[0] & index[1] & ~index[3] & ~index[4] & ~index[5] & ~index[6] & ~index[7] & index[10] & index[11]) | (~index[0] & ~index[1] & index[2] & index[3] & ~index[4] & ~index[6] & index[7] & ~index[8] & index[10]) | (~index[0] & index[1] & index[2] & index[3] & ~index[4] & ~index[5] & ~index[6] & ~index[7] & index[9] & index[11]) | (~index[0] & index[1] & ~index[2] & ~index[3] & index[4] & ~index[6] & ~index[7] & ~index[8] & index[9] & index[10]) | (~index[1] & index[2] & ~index[3] & index[4] & ~index[6] & index[7] & ~index[8] & ~index[9] & index[11]) | (index[0] & ~index[1] & index[2] & index[3] & ~index[4] & ~index[7] & index[8] & index[9] & index[10] & ~index[11]) | (index[0] & ~index[2] & ~index[3] & index[4] & index[6] & index[7] & ~index[8] & ~index[9] & index[11]) | (~index[0] & ~index[1] & ~index[2] & ~index[4] & ~index[6] & index[7] & ~index[8] & index[9] & ~index[10] & ~index[11]) | (index[0] & index[1] & index[3] & index[6] & ~index[8] & index[9] & ~index[10] & ~index[11]) | (~index[0] & index[1] & ~index[2] & ~index[3] & index[5] & ~index[6] & index[7] & ~index[8] & index[9] & index[10]) | (~index[0] & ~index[1] & index[2] & index[3] & ~index[4] & ~index[6] & index[7] & index[8] & ~index[10] & ~index[11]) | (~index[0] & ~index[1] & ~index[2] & ~index[3] & ~index[5] & ~index[6] & ~index[7] & index[8] & ~index[9] & index[10] & ~index[11]) | (index[0] & ~index[1] & ~index[2] & ~index[3] & ~index[4] & ~index[5] & index[8] & index[9] & ~index[10]) | (index[0] & ~index[1] & index[3] & index[4] & ~index[7] & ~index[8] & ~index[9] & index[11]) | (~index[0] & ~index[1] & ~index[2] & ~index[3] & index[5] & index[6] & index[8] & index[10] & ~index[11]) | (~index[0] & index[1] & ~index[2] & index[3] & index[4] & index[6] & index[7] & ~index[8] & index[11]) | (index[0] & ~index[1] & index[3] & ~index[4] & index[5] & ~index[6] & ~index[7]) | (index[0] & ~index[1] & ~index[3] & index[4] & index[6] & ~index[7] & index[8] & ~index[9] & index[11]) | (index[0] & index[1] & ~index[5] & index[6] & ~index[7] & index[10] & index[11]) | (~index[0] & index[1] & index[2] & index[3] & ~index[4] & index[6] & ~index[7] & ~index[9] & index[11]) | (~index[0] & ~index[1] & ~index[2] & ~index[3] & ~index[4] & ~index[5] & index[6] & ~index[7] & ~index[9] & ~index[10] & ~index[11]) | (~index[0] & ~index[1] & index[2] & ~index[4] & ~index[5] & index[6] & index[7] & ~index[8] & ~index[9] & ~index[10] & ~index[11]) | (~index[0] & ~index[1] & ~index[2] & ~index[4] & ~index[5] & ~index[6] & ~index[7] & ~index[8] & index[9] & index[10] & ~index[11]) | (index[1] & ~index[2] & ~index[3] & ~index[4] & ~index[5] & ~index[6] & index[7] & index[10] & index[11]) | (~index[0] & ~index[1] & index[3] & index[5] & ~index[6] & index[7] & ~index[9] & index[10]) | (index[0] & index[1] & index[2] & ~index[3] & ~index[4] & index[6] & index[8] & ~index[10] & index[11]) | (~index[0] & ~index[1] & ~index[2] & index[3] & index[4] & ~index[8] & ~index[9] & ~index[10] & ~index[11]) | (~index[0] & ~index[1] & ~index[2] & index[3] & ~index[4] & ~index[6] & ~index[7] & ~index[10] & ~index[11]) | (index[0] & ~index[1] & index[3] & ~index[4] & ~index[6] & ~index[7] & index[8] & ~index[10] & index[11]) | (index[0] & index[1] & index[2] & ~index[3] & index[5] & ~index[6] & index[7] & index[11]) | (~index[0] & ~index[1] & ~index[2] & index[3] & ~index[5] & index[6] & ~index[7] & index[10] & index[11]) | (~index[0] & ~index[1] & ~index[2] & ~index[3] & index[5] & index[6] & index[7] & index[8] & index[9]) | (~index[0] & index[1] & index[2] & ~index[3] & index[5] & index[6] & index[7] & index[9]) | (index[0] & ~index[1] & index[2] & ~index[3] & index[4] & ~index[7] & ~index[8] & index[9] & index[10]) | (index[0] & ~index[1] & index[2] & ~index[3] & ~index[4] & index[6] & index[8] & ~index[9] & ~index[10] & ~index[11]) | (index[0] & index[1] & ~index[2] & ~index[4] & ~index[6] & index[7] & index[8] & index[9] & index[10] & ~index[11]) | (~index[1] & ~index[2] & index[3] & ~index[4] & index[6] & ~index[7] & index[8] & index[9] & index[10] & ~index[11]) | (~index[0] & index[2] & ~index[3] & index[4] & index[6] & index[7] & index[8] & index[9] & index[10]) | (index[0] & ~index[2] & ~index[3] & index[5] & index[6] & index[7] & ~index[9] & index[10]) | (index[0] & index[1] & ~index[2] & index[3] & ~index[5] & ~index[6] & ~index[8] & ~index[9] & ~index[10]) | (~index[1] & ~index[2] & ~index[4] & ~index[5] & ~index[6] & ~index[7] & index[8] & index[9] & index[10] & index[11]) | (~index[0] & index[1] & index[2] & ~index[3] & ~index[4] & index[6] & index[7] & ~index[8] & index[9] & ~index[10]) | (index[0] & index[1] & ~index[2] & index[3] & ~index[4] & ~index[6] & ~index[7] & index[8] & index[9] & ~index[10]) | (~index[1] & index[2] & ~index[3] & ~index[4] & ~index[6] & ~index[7] & ~index[9] & ~index[10] & ~index[11]) | (index[0] & index[1] & ~index[2] & ~index[3] & index[4] & ~index[5] & index[6] & index[8] & index[11]) | (index[0] & index[1] & ~index[2] & index[3] & index[4] & index[6] & ~index[7] & ~index[9] & index[10]) | (~index[1] & index[2] & index[3] & ~index[4] & ~index[6] & ~index[7] & index[9] & index[10] & ~index[11]) | (~index[0] & ~index[1] & ~index[2] & index[3] & index[4] & index[6] & index[7] & ~index[8] & index[9] & index[10]) | (index[0] & ~index[1] & index[2] & ~index[3] & index[4] & ~index[6] & ~index[8] & ~index[9] & index[11]) | (~index[0] & index[1] & index[2] & ~index[3] & ~index[5] & index[7] & ~index[8] & ~index[9] & index[11]) | (index[0] & ~index[1] & index[2] & index[5] & ~index[7] & ~index[9] & index[10]) | (index[0] & index[1] & ~index[3] & ~index[4] & ~index[5] & ~index[6] & index[7] & ~index[9] & index[10]) | (~index[0] & ~index[1] & index[2] & ~index[3] & ~index[4] & ~index[5] & index[6] & ~index[7] & index[11]) | (index[0] & ~index[1] & ~index[2] & index[5] & ~index[6] & index[8] & ~index[9] & index[11]) | (~index[0] & index[1] & index[2] & ~index[3] & index[4] & index[7] & ~index[10] & index[11]) | (index[0] & ~index[1] & index[3] & ~index[4] & ~index[5] & index[6] & index[7] & ~index[8] & index[9] & index[10]) | (index[0] & index[1] & ~index[2] & index[4] & ~index[6] & index[7] & index[9] & ~index[10] & index[11]) | (index[0] & index[1] & ~index[2] & index[4] & index[6] & index[7] & index[9] & ~index[10] & ~index[11]) | (index[0] & ~index[1] & index[2] & index[3] & ~index[4] & ~index[5] & ~index[6] & index[7] & index[9] & index[11]) | (~index[0] & ~index[2] & ~index[3] & index[5] & ~index[6] & ~index[8] & ~index[9] & index[11]) | (index[0] & index[3] & index[4] & ~index[6] & index[7] & index[8] & index[10] & ~index[11]) | (~index[1] & index[2] & index[3] & index[4] & ~index[6] & index[7] & index[9] & index[10] & ~index[11]) | (index[0] & index[1] & index[2] & ~index[4] & ~index[5] & index[6] & index[7] & index[8] & index[9] & ~index[10]) | (index[0] & ~index[1] & ~index[2] & ~index[3] & index[4] & index[6] & index[10] & index[11]) | (~index[0] & index[1] & index[2] & index[3] & index[4] & index[6] & index[7] & ~index[8] & index[9]) | (~index[0] & ~index[1] & ~index[2] & ~index[3] & index[4] & ~index[6] & ~index[7] & index[8] & index[9] & ~index[11]) | (~index[1] & ~index[2] & index[3] & ~index[4] & index[6] & index[7] & index[8] & ~index[9] & ~index[10] & ~index[11]) | (~index[0] & ~index[1] & ~index[2] & index[3] & ~index[5] & ~index[6] & index[7] & ~index[8] & ~index[9] & index[11]) | (~index[0] & index[2] & ~index[3] & ~index[4] & ~index[6] & ~index[7] & ~index[10] & ~index[11]) | (~index[1] & ~index[2] & ~index[3] & index[4] & ~index[6] & ~index[7] & ~index[8] & index[9] & index[11]) | (~index[0] & ~index[1] & index[2] & ~index[3] & ~index[4] & index[7] & index[9] & ~index[10] & index[11]) | (index[0] & ~index[1] & ~index[2] & ~index[3] & ~index[5] & ~index[6] & index[7] & index[8] & index[9] & ~index[10]) | (index[0] & index[2] & ~index[3] & index[4] & index[6] & index[7] & ~index[8] & index[9] & index[10]) | (index[0] & index[1] & ~index[2] & index[3] & ~index[6] & ~index[7] & ~index[8] & ~index[9]) | (~index[0] & ~index[1] & ~index[2] & index[3] & index[4] & ~index[6] & index[7] & ~index[8] & index[11]) | (~index[0] & index[1] & index[2] & index[4] & ~index[6] & index[8] & index[9] & index[10] & ~index[11]) | (~index[0] & ~index[1] & index[2] & ~index[3] & ~index[4] & ~index[5] & ~index[6] & ~index[7] & ~index[8] & ~index[9]) | (index[0] & index[1] & index[2] & index[3] & ~index[4] & index[7] & ~index[8] & index[9] & index[10]) | (index[0] & index[1] & index[2] & index[3] & ~index[4] & index[6] & ~index[8] & ~index[9] & index[11]) | (~index[0] & index[1] & ~index[2] & index[5] & ~index[6] & ~index[7] & ~index[8] & index[11]) | (index[0] & ~index[1] & index[3] & ~index[4] & index[7] & index[9] & ~index[10] & index[11]) | (index[0] & ~index[1] & index[2] & ~index[3] & ~index[4] & ~index[5] & index[6] & index[7] & index[8] & index[9] & index[10] & ~index[11]) | (index[0] & ~index[1] & index[2] & index[3] & ~index[4] & ~index[6] & ~index[7] & index[8] & index[10] & ~index[11]) | (~index[1] & ~index[2] & ~index[3] & ~index[4] & index[6] & index[7] & index[8] & ~index[9] & index[10] & ~index[11]) | (~index[0] & ~index[1] & index[2] & index[3] & index[4] & ~index[6] & ~index[7] & index[9] & index[11]) | (index[0] & index[1] & ~index[2] & ~index[3] & ~index[4] & index[5] & ~index[7] & index[10] & index[11]) | (~index[0] & index[1] & ~index[2] & index[3] & ~index[5] & ~index[6] & index[7] & ~index[8] & index[9] & index[10]) | (~index[0] & ~index[1] & index[2] & ~index[3] & index[6] & ~index[7] & index[8] & ~index[9] & index[10]) | (index[0] & index[2] & index[4] & ~index[5] & ~index[6] & ~index[7] & index[10] & index[11]) | (index[0] & ~index[1] & index[2] & index[3] & index[7] & ~index[8] & ~index[9] & ~index[10] & ~index[11]) | (index[0] & index[1] & index[2] & index[3] & ~index[6] & index[7] & index[8] & ~index[9] & ~index[10]) | (~index[0] & ~index[1] & ~index[3] & ~index[4] & ~index[5] & ~index[6] & index[7] & index[8] & ~index[9] & ~index[10] & index[11]) | (~index[0] & ~index[1] & ~index[2] & index[3] & ~index[4] & index[7] & index[10] & index[11]) | (index[0] & index[1] & index[2] & index[3] & index[4] & ~index[7] & ~index[8] & index[9] & index[10]) | (index[0] & ~index[1] & index[2] & ~index[4] & index[5] & ~index[7] & index[9] & index[11]) | (index[0] & index[1] & ~index[3] & index[4] & ~index[5] & ~index[7] & index[10] & index[11]) | (index[0] & index[1] & ~index[2] & ~index[3] & index[5] & index[6] & ~index[8] & ~index[11]) | (index[1] & index[2] & index[4] & index[6] & index[7] & index[10] & index[11]) | (~index[0] & ~index[1] & index[2] & ~index[3] & ~index[4] & ~index[5] & index[8] & ~index[10] & index[11]) | (~index[0] & ~index[1] & index[2] & index[5] & index[6] & index[7] & ~index[8] & index[11]) | (index[0] & ~index[1] & index[2] & ~index[4] & index[6] & ~index[7] & ~index[8] & ~index[9] & index[10]) | (~index[0] & ~index[1] & index[2] & ~index[3] & ~index[4] & ~index[5] & ~index[6] & index[7] & index[8] & index[11]) | (~index[0] & index[1] & index[2] & ~index[3] & index[4] & ~index[6] & index[7] & index[9] & index[10] & ~index[11]) | (index[0] & ~index[1] & ~index[2] & index[3] & ~index[4] & index[6] & index[8] & ~index[10] & index[11]) | (~index[0] & index[1] & ~index[3] & index[4] & ~index[6] & index[7] & index[8] & ~index[9] & index[10]) | (index[0] & index[1] & ~index[2] & ~index[3] & index[4] & index[7] & index[8] & ~index[10] & index[11]) | (~index[0] & ~index[1] & index[2] & ~index[3] & ~index[4] & ~index[5] & index[6] & index[7] & ~index[8] & index[10]) | (index[0] & ~index[1] & index[3] & ~index[4] & ~index[5] & index[6] & index[7] & ~index[9] & ~index[10] & ~index[11]) | (~index[0] & index[1] & index[2] & index[3] & ~index[4] & index[6] & ~index[7] & ~index[8] & index[9] & index[10]) | (index[0] & ~index[1] & index[2] & index[3] & ~index[4] & ~index[6] & index[8] & index[9] & index[10] & ~index[11]) | (~index[0] & ~index[1] & index[2] & ~index[3] & ~index[4] & ~index[5] & index[6] & ~index[7] & ~index[8] & ~index[10]) | (index[0] & ~index[1] & index[2] & ~index[4] & ~index[5] & index[6] & index[7] & ~index[8] & ~index[9] & index[11]) | (index[0] & index[1] & index[2] & ~index[3] & ~index[4] & ~index[5] & index[6] & ~index[7] & index[8] & index[9] & index[10]) | (index[0] & ~index[1] & ~index[2] & index[3] & index[4] & ~index[7] & index[8] & index[9] & index[10] & ~index[11]) | (index[2] & index[3] & index[4] & index[6] & index[7] & index[9] & index[11]) | (index[1] & index[2] & index[3] & index[6] & index[7] & index[10] & index[11]) | (~index[1] & index[2] & ~index[3] & ~index[4] & index[5] & ~index[6] & ~index[7] & index[10] & index[11]) | (~index[0] & ~index[1] & ~index[2] & ~index[3] & ~index[4] & ~index[5] & ~index[6] & index[7] & ~index[10] & ~index[11]) | (~index[1] & index[2] & ~index[3] & index[5] & index[6] & index[9] & ~index[10]) | (~index[1] & index[2] & index[5] & ~index[6] & index[7] & ~index[8] & index[9]) | (index[0] & index[1] & index[2] & index[3] & ~index[4] & index[6] & ~index[7] & ~index[8] & index[11]) | (index[0] & index[1] & index[2] & ~index[3] & ~index[4] & ~index[6] & index[7] & index[9] & ~index[10] & index[11]) | (index[0] & ~index[2] & ~index[3] & ~index[4] & ~index[5] & index[6] & index[8] & index[9] & ~index[10]) | (~index[0] & index[1] & index[2] & ~index[4] & ~index[5] & index[6] & index[7] & ~index[8] & ~index[9] & index[10]) | (~index[1] & index[2] & index[3] & index[5] & index[6] & ~index[9]) | (index[0] & ~index[1] & ~index[2] & index[3] & index[4] & index[6] & index[7] & index[8] & ~index[10] & ~index[11]) | (index[0] & index[2] & index[5] & index[6] & index[8] & ~index[9]) | (~index[0] & index[1] & index[2] & index[3] & ~index[4] & ~index[5] & index[7] & ~index[8] & ~index[9] & index[10]) | (~index[0] & index[1] & index[2] & index[3] & ~index[4] & ~index[6] & ~index[7] & index[8] & ~index[9] & index[10]) | (~index[1] & ~index[2] & ~index[3] & ~index[4] & ~index[5] & index[6] & index[8] & index[9] & ~index[10] & ~index[11]) | (index[0] & ~index[1] & index[3] & index[4] & index[6] & ~index[7] & ~index[8] & index[11]) | (index[0] & ~index[1] & index[2] & index[3] & index[4] & index[6] & index[7] & index[8] & index[9]) | (index[1] & index[2] & index[4] & ~index[5] & ~index[6] & ~index[7] & index[10] & index[11]) | (~index[0] & index[2] & ~index[3] & index[4] & index[6] & index[7] & index[8] & ~index[9] & ~index[10] & ~index[11]) | (~index[0] & ~index[1] & index[2] & index[3] & ~index[4] & index[6] & index[7] & ~index[8] & ~index[10] & ~index[11]) | (index[0] & index[1] & ~index[2] & ~index[3] & ~index[4] & index[6] & ~index[7] & index[9] & index[11]) | (index[0] & ~index[3] & ~index[4] & ~index[5] & index[6] & ~index[7] & index[10] & index[11]) | (index[0] & index[1] & index[2] & ~index[3] & index[4] & index[6] & ~index[7] & ~index[9] & index[10]) | (~index[0] & index[1] & ~index[2] & index[3] & index[4] & ~index[6] & index[7] & index[8] & index[11]) | (~index[0] & index[1] & index[2] & index[3] & index[4] & ~index[6] & ~index[7] & index[9] & index[10]) | (index[0] & ~index[1] & ~index[2] & index[4] & index[6] & ~index[7] & ~index[8] & ~index[9] & index[10]) | (index[0] & index[1] & ~index[2] & ~index[3] & ~index[4] & index[6] & ~index[8] & ~index[9] & index[10]) | (index[0] & ~index[1] & ~index[2] & index[3] & ~index[4] & index[6] & ~index[7] & index[8] & index[10] & ~index[11]) | (~index[0] & index[1] & ~index[2] & ~index[4] & index[6] & ~index[7] & index[8] & ~index[9] & ~index[11]) | (~index[0] & index[1] & ~index[2] & index[3] & index[4] & index[6] & ~index[7] & ~index[8] & index[9]) | (~index[0] & index[3] & ~index[4] & ~index[5] & index[6] & ~index[7] & index[10] & index[11]) | (~index[0] & index[1] & ~index[2] & ~index[3] & index[6] & index[8] & ~index[9] & index[10]) | (index[0] & ~index[1] & ~index[2] & ~index[3] & ~index[5] & ~index[6] & index[7] & ~index[8] & index[10]) | (~index[1] & ~index[2] & ~index[3] & index[4] & ~index[6] & index[7] & ~index[8] & index[9] & index[10]) | (index[0] & index[1] & index[2] & ~index[3] & ~index[4] & ~index[5] & ~index[7] & ~index[8] & ~index[9] & index[11]) | (~index[0] & ~index[1] & ~index[3] & index[4] & ~index[6] & ~index[7] & index[8] & ~index[9] & index[11]) | (~index[0] & index[1] & index[2] & ~index[3] & index[5] & index[6] & index[9] & index[11]) | (index[0] & index[1] & index[2] & index[3] & ~index[5] & ~index[7] & index[10] & index[11]) | (~index[0] & index[1] & index[2] & ~index[3] & index[4] & ~index[8] & ~index[9] & index[11]) | (~index[0] & ~index[1] & ~index[2] & ~index[4] & ~index[6] & ~index[7] & ~index[8] & ~index[9] & ~index[10] & index[11]) | (index[0] & index[1] & ~index[2] & index[3] & index[4] & index[6] & index[9] & index[11]) | (~index[0] & index[1] & ~index[2] & index[3] & index[4] & index[7] & ~index[8] & ~index[9] & index[10]) | (index[0] & index[1] & ~index[2] & ~index[3] & index[5] & index[6] & index[7] & ~index[8]) | (index[1] & index[2] & index[3] & index[4] & ~index[7] & index[8] & index[9] & ~index[10]) | (index[0] & ~index[1] & index[2] & index[3] & ~index[4] & index[6] & index[7] & ~index[9] & ~index[10]) | (index[0] & index[1] & index[2] & index[3] & index[4] & ~index[6] & index[7] & ~index[10]) | (~index[0] & ~index[1] & ~index[2] & index[3] & ~index[5] & ~index[6] & ~index[7] & ~index[8] & index[10]) | (~index[0] & ~index[1] & index[2] & ~index[3] & index[4] & index[7] & ~index[8] & ~index[9] & index[10]) | (~index[0] & ~index[1] & ~index[2] & index[5] & index[6] & index[7] & index[8] & index[11]) | (index[0] & index[2] & index[3] & index[4] & ~index[6] & index[7] & ~index[8] & index[9] & index[10]) | (~index[0] & ~index[1] & index[2] & ~index[3] & ~index[6] & ~index[8] & index[9] & ~index[10] & ~index[11]) | (index[0] & index[1] & index[2] & ~index[3] & ~index[5] & ~index[6] & index[7] & ~index[8] & ~index[9] & index[10]) | (~index[0] & index[1] & index[2] & ~index[3] & index[4] & index[6] & ~index[7] & index[9] & ~index[11]) | (index[0] & index[2] & ~index[3] & ~index[4] & ~index[6] & ~index[7] & ~index[8] & index[9] & index[10]) | (~index[0] & ~index[1] & ~index[2] & ~index[3] & index[4] & index[6] & index[7] & index[8] & index[10]) | (~index[0] & ~index[2] & ~index[3] & ~index[4] & ~index[5] & index[6] & ~index[7] & ~index[8] & ~index[9] & index[10] & ~index[11]) | (index[0] & index[1] & index[3] & ~index[4] & index[6] & ~index[7] & ~index[8] & ~index[9] & index[11]) | (index[0] & index[1] & ~index[2] & ~index[3] & index[6] & index[7] & ~index[8] & ~index[9] & index[10]) | (index[1] & ~index[2] & index[3] & ~index[4] & ~index[5] & ~index[6] & index[7] & ~index[8] & ~index[9] & index[11]) | (index[0] & ~index[1] & ~index[2] & ~index[3] & ~index[5] & index[6] & ~index[7] & ~index[8] & index[9] & index[10]) | (index[1] & ~index[2] & ~index[3] & index[4] & ~index[5] & index[6] & ~index[7] & index[8] & index[9] & index[10]) | (~index[0] & ~index[1] & ~index[2] & index[4] & ~index[6] & ~index[7] & index[8] & ~index[10] & index[11]) | (index[0] & ~index[1] & ~index[4] & ~index[6] & ~index[8] & ~index[9] & ~index[10] & ~index[11]) | (~index[0] & ~index[2] & index[3] & index[4] & ~index[6] & ~index[7] & index[8] & ~index[9] & index[10]) | (index[0] & ~index[1] & ~index[2] & index[3] & index[5] & index[6] & ~index[8] & index[9]) | (~index[0] & index[1] & index[3] & index[6] & index[7] & index[10] & index[11]) | (index[0] & index[1] & ~index[2] & ~index[4] & index[6] & index[7] & ~index[8] & ~index[9] & index[10]) | (~index[0] & index[1] & index[2] & index[4] & index[6] & ~index[7] & index[8] & ~index[9] & index[10]) | (index[0] & ~index[1] & index[2] & index[3] & index[4] & index[6] & index[7] & ~index[9] & index[10]) | (~index[0] & index[1] & ~index[2] & ~index[3] & index[4] & index[6] & index[7] & ~index[8] & index[10]) | (index[0] & index[1] & index[2] & ~index[3] & index[4] & ~index[6] & index[7] & index[8] & index[9]) | (~index[0] & index[1] & ~index[3] & ~index[4] & ~index[7] & index[8] & ~index[9] & ~index[10] & ~index[11]) | (~index[0] & ~index[1] & index[2] & index[4] & ~index[6] & index[7] & index[8] & ~index[9] & index[10]) | (~index[0] & ~index[1] & ~index[2] & ~index[4] & ~index[5] & index[6] & index[8] & index[9] & index[10] & index[11]) | (~index[0] & index[1] & ~index[2] & index[3] & ~index[6] & index[7] & index[8] & ~index[9] & ~index[10] & ~index[11]) | (~index[0] & index[1] & index[2] & ~index[6] & index[7] & index[8] & index[9] & index[10] & ~index[11]) | (index[0] & index[1] & ~index[2] & ~index[4] & ~index[6] & ~index[7] & index[8] & ~index[9] & index[10]) | (index[0] & index[1] & ~index[3] & ~index[4] & ~index[6] & ~index[7] & ~index[8] & index[9] & index[10]) | (index[0] & ~index[1] & ~index[2] & index[4] & index[6] & index[7] & index[9] & index[11]) | (~index[0] & index[1] & index[2] & index[3] & index[4] & index[6] & index[7] & ~index[8] & ~index[10] & ~index[11]) | (~index[0] & index[1] & ~index[2] & ~index[3] & index[4] & ~index[6] & index[7] & index[9] & ~index[10] & ~index[11]) | (index[0] & index[1] & index[2] & index[3] & ~index[4] & index[6] & ~index[7] & index[8] & ~index[9] & index[10]) | (~index[0] & ~index[1] & ~index[2] & ~index[3] & index[4] & index[6] & ~index[7] & ~index[8] & ~index[9] & index[11]) | (~index[0] & index[1] & ~index[3] & ~index[4] & ~index[5] & index[6] & ~index[7] & index[8] & index[9] & ~index[11]) | (~index[0] & index[1] & index[2] & ~index[3] & index[6] & index[7] & index[8] & ~index[9] & ~index[10] & ~index[11]) | (index[0] & ~index[1] & index[2] & ~index[3] & ~index[4] & ~index[5] & index[6] & ~index[8] & ~index[9] & index[10]) | (~index[0] & ~index[1] & index[2] & ~index[3] & index[4] & ~index[8] & index[9] & ~index[10] & ~index[11]) | (index[1] & index[5] & index[6] & index[7] & index[9] & index[11]) | (~index[0] & ~index[1] & index[5] & index[7] & index[9] & ~index[10] & index[11]) | (index[0] & index[1] & ~index[2] & ~index[3] & index[4] & ~index[6] & ~index[7] & index[8] & index[9] & ~index[10]) | (~index[0] & index[1] & index[2] & ~index[3] & ~index[6] & index[7] & index[8] & index[10] & ~index[11]) | (index[0] & index[1] & ~index[2] & ~index[3] & ~index[4] & ~index[5] & ~index[6] & index[8] & index[10] & ~index[11]) | (~index[0] & index[1] & ~index[2] & index[4] & ~index[5] & ~index[6] & index[7] & index[10] & index[11]) | (~index[0] & ~index[1] & ~index[2] & ~index[3] & ~index[4] & ~index[5] & ~index[6] & index[7] & index[9] & ~index[11]) | (~index[0] & index[1] & ~index[2] & ~index[3] & ~index[4] & ~index[5] & index[6] & index[7] & index[8] & ~index[10] & index[11]) | (index[1] & ~index[2] & index[3] & index[4] & index[6] & index[7] & index[8] & index[9] & index[10]);

assign val[5] = (index[0] & ~index[2] & ~index[4] & index[6] & index[7] & index[8] & index[9] & ~index[11]) | (~index[0] & index[1] & ~index[3] & ~index[5] & ~index[6] & index[7] & ~index[8]) | (index[0] & index[1] & ~index[2] & ~index[3] & ~index[6] & index[11]) | (index[0] & ~index[2] & index[3] & index[6] & ~index[7] & ~index[11]) | (index[1] & ~index[2] & ~index[3] & ~index[4] & ~index[6] & index[8] & index[10]) | (index[0] & ~index[1] & ~index[3] & index[5] & ~index[6] & index[10]) | (~index[1] & ~index[4] & index[6] & ~index[7] & index[8] & index[9] & index[10] & index[11]) | (~index[0] & index[1] & index[3] & ~index[4] & ~index[9] & ~index[10] & ~index[11]) | (~index[1] & ~index[2] & ~index[3] & index[4] & index[6] & ~index[9]) | (index[2] & ~index[3] & ~index[4] & ~index[5] & index[6] & ~index[8] & index[9]) | (~index[0] & index[1] & ~index[3] & ~index[5] & index[7] & index[8] & ~index[10] & ~index[11]) | (~index[0] & index[1] & index[2] & index[4] & ~index[9] & ~index[11]) | (index[0] & ~index[1] & ~index[3] & ~index[4] & ~index[6] & ~index[8]) | (index[0] & ~index[1] & ~index[2] & ~index[4] & index[5] & index[9]) | (index[0] & ~index[1] & ~index[6] & index[9] & ~index[10] & ~index[11]) | (index[1] & ~index[2] & ~index[3] & ~index[4] & index[6] & ~index[9] & index[11]) | (index[1] & index[2] & ~index[3] & ~index[5] & ~index[6] & index[8] & ~index[9]) | (index[1] & ~index[2] & ~index[3] & ~index[5] & index[7] & index[9] & ~index[11]) | (~index[1] & ~index[2] & index[4] & ~index[7] & index[8] & index[11]) | (~index[0] & index[1] & ~index[2] & index[3] & ~index[4] & ~index[6] & index[8]) | (~index[1] & index[2] & index[3] & index[4] & index[9] & index[11]) | (~index[0] & ~index[1] & index[2] & index[6] & ~index[7] & index[9]) | (index[2] & ~index[3] & index[4] & index[6] & ~index[7] & index[8] & ~index[10]) | (~index[0] & index[2] & ~index[3] & index[4] & index[8] & ~index[10]) | (index[1] & index[3] & ~index[4] & ~index[6] & ~index[8] & ~index[10]) | (index[0] & ~index[1] & ~index[2] & index[3] & index[7] & index[11]) | (~index[1] & ~index[3] & index[4] & ~index[8] & index[9] & index[10]) | (~index[0] & ~index[1] & ~index[2] & ~index[5] & index[6] & ~index[8] & ~index[9] & ~index[10] & ~index[11]) | (index[0] & ~index[2] & ~index[3] & ~index[6] & ~index[7] & index[11]) | (index[2] & ~index[3] & index[5] & ~index[8] & ~index[9] & ~index[11]) | (~index[0] & ~index[2] & index[3] & ~index[5] & ~index[6] & index[7] & ~index[9] & ~index[11]) | (~index[1] & index[3] & ~index[7] & index[10] & index[11]) | (index[3] & ~index[4] & ~index[5] & index[6] & index[8] & index[10]) | (~index[0] & ~index[1] & index[3] & ~index[4] & index[6] & index[11]) | (~index[0] & ~index[2] & index[5] & index[6] & index[7] & ~index[9]) | (index[0] & ~index[1] & index[3] & ~index[4] & index[7] & ~index[10] & ~index[11]) | (index[2] & ~index[3] & ~index[4] & ~index[7] & index[10] & index[11]) | (~index[0] & index[1] & ~index[2] & ~index[3] & index[7] & ~index[8] & ~index[9]) | (~index[0] & index[3] & ~index[5] & index[6] & index[7] & index[10]) | (index[0] & ~index[1] & ~index[4] & index[6] & index[7] & index[8] & ~index[11]) | (index[1] & ~index[2] & ~index[4] & ~index[5] & index[6] & index[9] & index[10] & ~index[11]) | (~index[1] & ~index[2] & index[3] & index[6] & ~index[8] & ~index[10] & ~index[11]) | (index[2] & ~index[5] & index[6] & ~index[7] & ~index[8] & index[9]) | (index[0] & index[1] & ~index[3] & ~index[5] & index[6] & ~index[8] & ~index[10]) | (~index[1] & ~index[2] & index[5] & index[9] & index[11]) | (~index[1] & index[2] & index[3] & index[6] & index[10]) | (index[0] & index[2] & ~index[5] & index[7] & ~index[8] & ~index[9] & index[10]) | (~index[1] & index[3] & ~index[5] & index[6] & ~index[9] & index[10]) | (~index[1] & ~index[2] & index[4] & ~index[9] & index[10]) | (index[0] & ~index[4] & ~index[5] & ~index[6] & index[9] & ~index[10] & ~index[11]) | (index[1] & ~index[3] & index[4] & ~index[5] & index[7] & index[11]) | (~index[0] & index[2] & index[8] & ~index[9] & ~index[10] & ~index[11]) | (~index[0] & ~index[1] & index[4] & index[6] & index[7] & index[8] & ~index[10] & ~index[11]) | (~index[0] & index[1] & index[2] & ~index[3] & ~index[8] & index[10]) | (index[0] & ~index[2] & index[3] & index[4] & ~index[7] & ~index[9]) | (~index[0] & ~index[1] & ~index[3] & index[4] & ~index[10] & index[11]) | (index[0] & ~index[4] & ~index[6] & index[7] & ~index[8] & ~index[9] & index[11]) | (index[0] & ~index[2] & index[3] & index[6] & index[8] & index[9]) | (~index[0] & index[3] & ~index[4] & ~index[5] & index[9] & index[11]) | (index[1] & index[3] & ~index[7] & ~index[9] & ~index[10] & ~index[11]) | (index[0] & ~index[2] & index[3] & ~index[4] & index[6] & index[7] & index[8]) | (~index[0] & ~index[1] & ~index[2] & index[5] & ~index[8] & index[10]) | (~index[1] & ~index[3] & ~index[6] & ~index[7] & ~index[8] & ~index[9] & ~index[10] & index[11]) | (~index[0] & index[2] & ~index[3] & ~index[5] & index[6] & index[8] & index[11]) | (index[0] & index[4] & ~index[5] & index[7] & index[8] & index[9] & index[10]) | (index[0] & ~index[1] & ~index[2] & index[8] & index[9] & ~index[10]) | (~index[0] & ~index[1] & index[3] & ~index[4] & index[7] & ~index[8] & index[10]) | (index[0] & index[2] & index[6] & ~index[8] & ~index[10] & ~index[11]) | (index[0] & ~index[2] & index[4] & ~index[7] & ~index[9] & ~index[11]) | (~index[1] & index[3] & index[6] & ~index[7] & ~index[8] & ~index[9]) | (index[1] & ~index[2] & ~index[5] & ~index[6] & ~index[7] & index[8] & index[11]) | (~index[0] & index[2] & ~index[4] & ~index[5] & index[6] & index[7] & index[10]) | (index[0] & ~index[4] & ~index[5] & index[6] & ~index[7] & index[8] & index[10]) | (index[0] & ~index[1] & index[8] & ~index[9] & index[10]) | (index[1] & ~index[2] & ~index[3] & ~index[4] & ~index[5] & index[6] & index[8] & ~index[11]) | (index[0] & index[2] & ~index[5] & ~index[6] & index[7] & index[8] & index[11]) | (index[2] & ~index[4] & ~index[5] & index[6] & index[9] & index[11]) | (index[0] & ~index[2] & index[3] & ~index[5] & ~index[8] & ~index[9] & ~index[10]) | (~index[0] & ~index[3] & index[4] & index[6] & index[8] & index[11]) | (~index[0] & index[2] & ~index[5] & index[6] & ~index[8] & index[10]) | (~index[1] & index[2] & ~index[3] & index[4] & index[9] & index[10] & ~index[11]) | (index[0] & ~index[1] & ~index[3] & ~index[6] & ~index[8] & index[9]) | (index[0] & ~index[2] & ~index[4] & ~index[5] & index[7] & index[8] & ~index[11]) | (index[2] & ~index[4] & ~index[5] & index[6] & ~index[7] & index[8] & index[11]) | (index[0] & ~index[1] & index[2] & ~index[3] & ~index[9] & index[11]) | (index[0] & index[2] & ~index[3] & index[6] & ~index[9] & ~index[10] & ~index[11]) | (index[0] & index[1] & index[4] & index[7] & ~index[8] & ~index[9]) | (index[0] & ~index[2] & index[4] & ~index[8] & ~index[9] & ~index[11]) | (~index[1] & index[2] & ~index[4] & ~index[5] & ~index[8] & index[10]) | (index[1] & index[2] & ~index[3] & index[4] & ~index[6] & ~index[9]) | (~index[1] & index[2] & index[3] & index[4] & ~index[6] & index[7] & ~index[8] & index[9]) | (~index[0] & index[3] & ~index[5] & index[6] & ~index[7] & ~index[8] & ~index[10]) | (~index[0] & index[1] & index[3] & index[4] & index[8] & index[9] & ~index[11]) | (index[1] & index[2] & ~index[3] & index[4] & ~index[7] & index[10]) | (~index[0] & index[2] & ~index[4] & ~index[6] & index[10] & index[11]) | (~index[0] & ~index[1] & ~index[2] & ~index[3] & index[4] & ~index[7] & index[10]) | (index[1] & ~index[2] & index[3] & index[5] & index[6] & index[7] & index[10]) | (~index[1] & ~index[2] & index[4] & ~index[7] & ~index[8] & ~index[11]) | (index[0] & ~index[2] & ~index[5] & ~index[7] & ~index[8] & ~index[9]) | (index[2] & ~index[6] & ~index[7] & index[8] & ~index[9] & index[10]) | (index[0] & index[1] & ~index[5] & index[10] & index[11]) | (index[1] & index[4] & index[7] & index[8] & index[9] & ~index[10]) | (index[1] & ~index[4] & ~index[5] & index[6] & ~index[7] & index[9] & index[10]) | (~index[0] & ~index[1] & index[2] & ~index[3] & ~index[5] & index[6] & index[9]) | (index[1] & ~index[3] & index[4] & index[6] & ~index[7] & ~index[9] & ~index[11]) | (index[0] & ~index[2] & index[3] & ~index[4] & index[8] & ~index[10] & ~index[11]) | (index[1] & index[4] & ~index[8] & ~index[9] & index[10]) | (~index[0] & ~index[1] & index[2] & ~index[4] & ~index[5] & index[7] & index[8] & index[9]) | (~index[0] & ~index[1] & ~index[3] & index[5] & index[8] & ~index[10] & ~index[11]) | (index[0] & index[3] & ~index[4] & ~index[5] & index[6] & index[8] & index[9]) | (~index[1] & ~index[2] & index[3] & ~index[5] & index[8] & ~index[9] & index[10]) | (~index[1] & index[3] & ~index[5] & index[6] & index[7] & index[8] & index[9]) | (index[0] & index[1] & index[3] & ~index[5] & ~index[6] & ~index[8] & ~index[11]) | (~index[0] & index[2] & index[5] & ~index[7] & ~index[8]) | (~index[1] & ~index[2] & index[4] & index[10] & index[11]) | (index[0] & ~index[1] & index[3] & index[4] & index[7] & index[9]) | (index[0] & ~index[2] & ~index[3] & ~index[5] & ~index[9] & index[10]) | (~index[1] & index[2] & ~index[3] & ~index[4] & index[6] & ~index[9]) | (index[2] & ~index[3] & index[5] & index[6] & index[7] & ~index[11]) | (~index[0] & ~index[1] & index[2] & ~index[3] & ~index[4] & ~index[5] & index[10]) | (~index[1] & ~index[2] & index[3] & ~index[4] & ~index[6] & ~index[7] & index[9]) | (~index[0] & index[1] & index[2] & ~index[5] & ~index[6] & ~index[7] & index[8]) | (index[1] & index[3] & ~index[4] & index[7] & index[8] & index[10]) | (~index[0] & index[2] & index[3] & ~index[4] & ~index[7] & ~index[10]) | (~index[0] & ~index[6] & index[7] & ~index[8] & ~index[9] & ~index[10] & ~index[11]) | (index[0] & ~index[2] & ~index[3] & ~index[6] & index[9] & index[10]) | (index[1] & index[2] & ~index[5] & ~index[6] & ~index[7] & index[8] & index[10]) | (index[0] & index[2] & index[3] & index[4] & index[9] & index[10]) | (index[1] & index[2] & index[3] & ~index[4] & index[7] & index[11]) | (~index[1] & ~index[2] & index[5] & ~index[6] & ~index[8]) | (index[1] & ~index[2] & ~index[4] & index[6] & ~index[7] & index[10] & ~index[11]) | (index[1] & index[2] & index[3] & ~index[6] & index[9] & index[10]) | (~index[0] & index[2] & index[5] & index[6] & ~index[7]) | (~index[0] & ~index[1] & ~index[3] & index[5] & index[6] & index[7] & ~index[11]) | (index[1] & ~index[2] & index[4] & index[6] & index[9] & ~index[10]) | (~index[0] & index[1] & ~index[2] & ~index[4] & ~index[5] & ~index[7] & index[10]) | (~index[0] & ~index[1] & index[4] & ~index[6] & ~index[7] & ~index[9]) | (~index[1] & ~index[3] & index[5] & ~index[6] & index[7] & index[8] & index[9]) | (~index[2] & index[4] & index[6] & index[10] & index[11]) | (index[0] & index[1] & ~index[2] & index[3] & ~index[6] & ~index[8]) | (index[0] & ~index[6] & index[7] & ~index[8] & index[9] & ~index[11]) | (index[0] & ~index[1] & ~index[3] & ~index[4] & index[7] & ~index[8] & index[9]) | (index[1] & ~index[2] & ~index[4] & ~index[5] & ~index[6] & ~index[8] & index[11]) | (index[0] & ~index[1] & ~index[2] & ~index[5] & index[6] & ~index[7] & ~index[9]) | (~index[1] & index[2] & ~index[3] & ~index[4] & ~index[7] & index[8] & index[10]) | (~index[0] & ~index[5] & index[6] & ~index[7] & ~index[8] & index[9] & ~index[10] & index[11]) | (index[0] & ~index[2] & ~index[3] & ~index[4] & ~index[5] & index[10] & ~index[11]) | (~index[0] & index[1] & ~index[2] & ~index[3] & ~index[6] & index[7] & ~index[11]) | (index[2] & index[3] & index[4] & ~index[9] & ~index[10] & ~index[11]) | (~index[0] & index[2] & ~index[5] & index[7] & ~index[8] & index[11]) | (~index[0] & index[1] & index[4] & index[7] & ~index[8] & index[10]) | (~index[0] & index[4] & ~index[6] & index[7] & ~index[8] & ~index[9] & ~index[10]) | (index[1] & index[2] & index[3] & ~index[4] & ~index[8] & ~index[10]) | (~index[0] & ~index[3] & index[5] & index[6] & index[7] & ~index[8]) | (index[0] & index[1] & index[4] & ~index[6] & index[9] & index[10]) | (~index[0] & index[1] & ~index[2] & ~index[3] & index[5] & ~index[7] & index[8]) | (index[0] & index[1] & index[2] & index[3] & ~index[5] & ~index[7] & index[9]) | (index[1] & ~index[2] & index[3] & ~index[4] & index[7] & index[8] & ~index[11]) | (~index[1] & ~index[2] & index[5] & ~index[6] & index[9]) | (index[0] & index[1] & ~index[2] & ~index[3] & ~index[6] & ~index[7]) | (~index[1] & index[2] & ~index[4] & ~index[8] & ~index[9] & index[10]) | (index[0] & ~index[5] & index[6] & index[7] & ~index[8] & ~index[9] & index[11]) | (index[0] & index[1] & index[2] & index[4] & index[8] & index[11]) | (index[1] & ~index[2] & index[4] & index[7] & ~index[10] & index[11]) | (~index[1] & ~index[2] & ~index[3] & ~index[4] & index[5] & index[7] & ~index[11]) | (index[0] & index[1] & ~index[4] & ~index[5] & ~index[7] & index[9] & index[11]) | (index[1] & ~index[2] & ~index[3] & index[6] & index[7] & ~index[8] & ~index[10]) | (index[1] & ~index[2] & ~index[5] & ~index[7] & index[9] & index[11]) | (~index[1] & ~index[2] & index[5] & ~index[7] & index[11]) | (index[2] & ~index[3] & ~index[4] & ~index[6] & ~index[7] & ~index[9] & ~index[11]) | (~index[1] & index[2] & ~index[4] & ~index[5] & ~index[7] & index[8] & index[11]) | (index[0] & index[4] & index[7] & index[8] & index[11]) | (~index[0] & index[3] & ~index[4] & ~index[5] & index[8] & index[11]) | (~index[0] & index[1] & index[2] & ~index[6] & index[7] & ~index[9] & ~index[11]) | (~index[0] & ~index[1] & index[4] & ~index[5] & ~index[6] & ~index[7] & index[8]) | (index[1] & ~index[3] & index[4] & ~index[9] & ~index[10] & ~index[11]) | (~index[1] & ~index[2] & index[4] & ~index[6] & index[9] & ~index[10] & ~index[11]) | (index[0] & ~index[1] & ~index[3] & index[6] & index[8] & ~index[9]) | (index[0] & index[2] & index[3] & index[4] & index[7] & ~index[11]) | (~index[1] & index[2] & index[4] & index[7] & index[8] & ~index[9]) | (~index[0] & ~index[2] & ~index[3] & index[4] & index[6] & ~index[8]) | (~index[1] & index[2] & ~index[3] & ~index[4] & ~index[8] & index[11]);

assign val[6] = (~index[0] & ~index[1] & index[5] & index[6] & ~index[7] & index[9]) | (~index[1] & index[2] & ~index[4] & ~index[7] & index[8] & ~index[10] & index[11]) | (index[1] & index[2] & index[3] & ~index[4] & ~index[6] & index[9] & index[11]) | (~index[1] & ~index[3] & ~index[5] & index[6] & ~index[8] & index[9] & index[10] & ~index[11]) | (index[0] & index[1] & ~index[2] & index[8] & index[9] & index[10] & ~index[11]) | (~index[0] & index[1] & index[3] & ~index[4] & index[7] & index[8] & index[9] & ~index[11]) | (~index[1] & ~index[2] & index[3] & index[4] & ~index[7] & index[10] & index[11]) | (~index[1] & index[2] & ~index[3] & ~index[4] & index[7] & index[9] & ~index[10]) | (~index[0] & ~index[2] & ~index[4] & ~index[5] & index[7] & index[8] & ~index[11]) | (index[0] & ~index[1] & index[3] & index[6] & index[7] & index[10] & ~index[11]) | (~index[0] & index[2] & index[3] & index[4] & ~index[6] & index[7] & index[8]) | (~index[0] & ~index[1] & index[2] & ~index[3] & ~index[4] & ~index[10] & index[11]) | (~index[1] & index[2] & index[4] & index[6] & index[7] & ~index[8] & ~index[9] & ~index[11]) | (~index[0] & index[2] & index[6] & ~index[8] & index[9] & index[11]) | (index[1] & index[5] & ~index[6] & index[7] & ~index[9] & index[11]) | (index[1] & index[2] & index[3] & index[7] & ~index[9] & index[11]) | (index[1] & ~index[3] & index[4] & index[7] & index[8] & index[9] & ~index[11]) | (index[0] & index[1] & ~index[2] & ~index[4] & index[7] & index[8] & index[9] & ~index[11]) | (index[0] & ~index[1] & ~index[2] & ~index[3] & index[6] & index[7] & ~index[8]) | (index[0] & index[2] & ~index[3] & index[4] & ~index[6] & ~index[7] & ~index[9]) | (index[0] & index[1] & ~index[2] & ~index[6] & ~index[8] & ~index[9] & ~index[10]) | (~index[0] & ~index[1] & index[4] & index[5]) | (~index[0] & ~index[1] & ~index[2] & index[3] & ~index[6] & index[9] & index[11]) | (~index[0] & ~index[3] & ~index[4] & ~index[6] & index[7] & ~index[8] & index[9] & ~index[11]) | (~index[0] & index[1] & ~index[2] & ~index[3] & index[4] & ~index[6] & index[9]) | (index[0] & index[1] & ~index[3] & index[4] & ~index[5] & ~index[6] & ~index[7]) | (~index[0] & index[4] & index[6] & index[7] & ~index[8] & ~index[9] & ~index[10] & ~index[11]) | (~index[0] & ~index[4] & ~index[5] & index[7] & ~index[8] & ~index[9] & ~index[10] & index[11]) | (index[1] & ~index[2] & index[3] & index[4] & ~index[7] & ~index[9] & index[10]) | (~index[0] & ~index[1] & index[2] & index[6] & index[7] & index[10] & ~index[11]) | (~index[0] & index[1] & index[2] & index[6] & ~index[7] & index[8] & ~index[10]) | (index[0] & ~index[2] & index[6] & ~index[8] & index[9] & index[11]) | (~index[0] & index[1] & ~index[3] & ~index[4] & ~index[6] & index[7] & index[8] & ~index[9]) | (index[0] & index[1] & ~index[2] & index[6] & ~index[7] & index[8] & ~index[9] & ~index[10]) | (index[1] & ~index[2] & index[3] & ~index[4] & index[8] & ~index[10] & ~index[11]) | (index[0] & index[1] & index[2] & index[3] & ~index[8] & index[11]) | (~index[0] & index[1] & ~index[2] & ~index[3] & ~index[4] & ~index[7] & ~index[9]) | (~index[0] & index[3] & index[4] & index[6] & index[7] & ~index[10] & index[11]) | (index[1] & index[2] & index[3] & ~index[6] & ~index[7] & ~index[8]) | (index[0] & index[1] & ~index[2] & ~index[3] & index[5] & index[7] & index[11]) | (~index[0] & ~index[1] & ~index[2] & ~index[3] & ~index[5] & index[8] & ~index[9] & ~index[10]) | (~index[0] & ~index[1] & ~index[2] & ~index[7] & ~index[8] & index[10] & ~index[11]) | (~index[2] & ~index[3] & ~index[4] & ~index[5] & index[10] & ~index[11]) | (index[0] & index[2] & ~index[3] & ~index[4] & ~index[5] & index[6] & index[9] & ~index[10] & ~index[11]) | (~index[0] & ~index[1] & index[4] & ~index[7] & ~index[8] & ~index[9] & ~index[10]) | (index[1] & index[4] & ~index[7] & ~index[8] & ~index[9] & index[10]) | (~index[0] & ~index[2] & index[3] & index[4] & index[6] & ~index[9] & index[11]) | (~index[0] & ~index[1] & ~index[2] & index[4] & ~index[6] & ~index[7] & ~index[10]) | (index[0] & index[2] & index[3] & ~index[4] & ~index[7] & index[8] & index[10] & ~index[11]) | (index[0] & ~index[1] & ~index[5] & ~index[6] & index[7] & ~index[9] & index[10]) | (index[0] & index[2] & ~index[3] & ~index[4] & ~index[5] & index[7] & index[10]) | (index[0] & ~index[1] & index[3] & index[4] & index[8] & index[9] & ~index[11]) | (~index[0] & ~index[1] & index[2] & index[8] & ~index[9] & index[10]) | (~index[0] & index[2] & ~index[4] & ~index[6] & ~index[9] & index[10]) | (index[0] & ~index[1] & ~index[4] & index[8] & ~index[9] & index[11]) | (index[0] & index[3] & index[5] & index[9] & ~index[11]) | (index[0] & index[2] & index[6] & index[7] & index[8] & ~index[9] & index[10]) | (index[0] & ~index[1] & index[2] & index[3] & ~index[7] & ~index[9] & ~index[10]) | (~index[0] & ~index[1] & index[5] & ~index[8] & index[9]) | (index[0] & index[1] & index[3] & ~index[5] & ~index[6] & index[7] & index[11]) | (index[2] & ~index[3] & ~index[4] & index[7] & ~index[8] & index[10]) | (index[0] & index[3] & index[4] & index[6] & index[9] & ~index[10]) | (index[1] & ~index[2] & index[3] & ~index[4] & ~index[6] & index[7] & ~index[8] & ~index[9]) | (~index[1] & ~index[3] & ~index[4] & index[6] & index[8] & ~index[9] & ~index[10]) | (index[0] & index[1] & ~index[2] & index[4] & ~index[6] & index[8] & index[10] & ~index[11]) | (~index[2] & ~index[3] & ~index[5] & ~index[6] & index[7] & index[9] & index[10] & ~index[11]) | (index[0] & index[2] & index[6] & index[7] & ~index[8] & index[9] & index[10]) | (~index[2] & ~index[4] & ~index[5] & index[6] & index[8] & ~index[9] & ~index[11]) | (~index[1] & index[5] & ~index[7] & ~index[9] & index[11]) | (~index[2] & ~index[4] & ~index[6] & index[7] & ~index[8] & ~index[9] & ~index[10] & index[11]) | (index[2] & ~index[3] & index[5] & ~index[6] & ~index[8] & index[10]) | (~index[0] & ~index[1] & ~index[2] & ~index[5] & index[6] & ~index[9] & ~index[10] & index[11]) | (index[0] & index[2] & index[4] & ~index[6] & index[8] & ~index[10] & ~index[11]) | (~index[1] & ~index[4] & ~index[6] & ~index[7] & index[9] & index[10] & ~index[11]) | (index[0] & index[2] & index[6] & ~index[7] & ~index[8] & ~index[9] & index[10]) | (~index[0] & index[1] & ~index[3] & index[4] & ~index[5] & ~index[6] & index[11]) | (~index[0] & index[1] & ~index[3] & ~index[4] & index[6] & index[7] & index[9] & index[11]) | (index[0] & ~index[2] & ~index[3] & index[6] & ~index[8] & index[11]) | (~index[1] & ~index[2] & ~index[3] & ~index[6] & index[7] & index[8] & ~index[11]) | (~index[0] & ~index[1] & index[2] & ~index[4] & index[6] & index[7] & index[10]) | (index[0] & index[2] & index[3] & ~index[4] & ~index[6] & index[11]) | (~index[0] & index[3] & ~index[5] & ~index[6] & ~index[8] & index[9] & index[10]) | (~index[2] & ~index[3] & ~index[4] & ~index[5] & index[7] & index[8] & ~index[11]) | (index[0] & index[1] & ~index[3] & ~index[4] & index[7] & ~index[8] & ~index[9] & ~index[11]) | (index[1] & ~index[2] & index[3] & index[5] & index[6] & index[10]) | (index[1] & index[2] & ~index[4] & ~index[7] & index[8] & ~index[9] & index[10]) | (~index[1] & ~index[2] & ~index[3] & index[4] & ~index[6] & index[7] & ~index[9] & ~index[11]) | (~index[0] & index[1] & ~index[3] & index[6] & index[7] & ~index[8] & ~index[10]) | (~index[1] & index[2] & ~index[3] & ~index[6] & index[9] & ~index[10] & ~index[11]) | (index[1] & ~index[2] & index[6] & index[7] & index[9] & ~index[10] & ~index[11]) | (~index[0] & index[2] & ~index[3] & ~index[5] & ~index[7] & ~index[10] & index[11]) | (index[1] & ~index[2] & ~index[4] & ~index[5] & ~index[8] & index[9] & index[10]) | (~index[0] & index[3] & ~index[4] & ~index[5] & index[7] & index[9] & ~index[10] & ~index[11]) | (~index[0] & index[1] & ~index[2] & ~index[3] & index[8] & index[10] & ~index[11]) | (index[0] & index[2] & ~index[4] & ~index[6] & index[7] & index[9] & index[11]) | (~index[0] & ~index[2] & index[6] & index[7] & index[8] & index[10] & ~index[11]) | (index[1] & ~index[4] & ~index[5] & index[6] & ~index[8] & ~index[9] & index[11]) | (index[1] & ~index[2] & ~index[3] & ~index[5] & index[7] & index[8] & index[10] & ~index[11]) | (~index[1] & ~index[2] & ~index[5] & ~index[6] & ~index[8] & index[9] & ~index[10] & index[11]) | (index[1] & ~index[3] & ~index[5] & ~index[6] & index[8] & index[9] & index[10] & ~index[11]) | (index[2] & ~index[3] & ~index[4] & ~index[5] & ~index[6] & ~index[7] & index[8] & index[9] & ~index[11]) | (~index[1] & index[3] & index[4] & index[6] & index[7] & index[8] & index[9] & ~index[11]) | (~index[1] & ~index[2] & ~index[3] & index[5] & index[6] & ~index[7] & index[9]) | (~index[0] & index[2] & index[6] & ~index[7] & ~index[8] & index[9]) | (~index[0] & ~index[1] & index[3] & ~index[5] & index[6] & ~index[8] & ~index[9]) | (~index[1] & ~index[2] & index[3] & ~index[6] & ~index[7] & ~index[10] & ~index[11]) | (~index[2] & ~index[3] & ~index[4] & index[6] & ~index[7] & index[9] & index[10] & ~index[11]) | (index[1] & index[2] & ~index[3] & index[6] & ~index[8] & ~index[10] & ~index[11]) | (index[0] & ~index[1] & ~index[3] & index[8] & ~index[10] & index[11]) | (~index[1] & ~index[2] & index[3] & ~index[4] & ~index[6] & index[9] & ~index[10]) | (~index[0] & ~index[1] & index[2] & ~index[3] & index[6] & ~index[8] & index[9]) | (index[0] & ~index[1] & ~index[3] & ~index[4] & ~index[5] & index[6] & ~index[8] & index[9]) | (~index[0] & index[1] & ~index[2] & ~index[3] & ~index[6] & ~index[7] & index[8]) | (index[0] & index[1] & ~index[2] & index[3] & index[4] & index[6] & ~index[8] & ~index[11]) | (index[2] & index[3] & index[4] & ~index[6] & index[7] & index[10]) | (~index[0] & ~index[2] & ~index[4] & ~index[5] & index[7] & index[8] & index[9] & index[10]) | (index[0] & ~index[1] & ~index[3] & ~index[5] & ~index[6] & index[7] & index[11]) | (index[1] & index[3] & ~index[4] & ~index[7] & ~index[9] & ~index[10] & ~index[11]) | (~index[0] & ~index[3] & index[5] & index[6] & index[8] & index[9] & ~index[11]) | (index[0] & ~index[2] & ~index[4] & index[6] & ~index[7] & ~index[10] & index[11]) | (~index[1] & index[2] & index[3] & ~index[4] & index[7] & ~index[9] & ~index[11]) | (~index[0] & index[2] & index[4] & ~index[5] & ~index[6] & index[7] & index[8] & index[9]) | (~index[0] & index[2] & index[3] & index[4] & index[6] & ~index[7] & index[10]) | (index[1] & ~index[3] & ~index[5] & ~index[6] & ~index[7] & ~index[10] & index[11]) | (~index[0] & ~index[1] & ~index[2] & index[3] & index[7] & ~index[8] & ~index[10]) | (~index[1] & ~index[3] & ~index[4] & index[5] & ~index[6] & index[7] & index[10]) | (~index[2] & index[3] & ~index[4] & index[6] & index[7] & index[8]) | (~index[0] & ~index[1] & ~index[3] & ~index[4] & ~index[7] & index[10] & ~index[11]) | (~index[0] & index[1] & index[3] & ~index[6] & index[7] & index[8] & index[9]) | (index[2] & index[4] & index[6] & ~index[7] & ~index[8] & index[9]) | (~index[0] & index[1] & ~index[2] & index[4] & ~index[5] & ~index[6] & index[9] & index[10]) | (~index[2] & index[4] & index[6] & index[7] & ~index[9] & index[11]) | (~index[0] & index[2] & ~index[4] & ~index[5] & index[6] & index[7] & ~index[8] & ~index[9]) | (index[0] & index[1] & index[5] & index[6] & index[8] & index[11]) | (~index[1] & index[3] & index[4] & ~index[7] & ~index[8] & ~index[9] & index[11]) | (~index[2] & ~index[4] & ~index[5] & ~index[6] & index[8] & index[9] & index[10] & index[11]) | (index[0] & ~index[1] & ~index[3] & ~index[6] & ~index[7] & index[8] & index[11]) | (index[0] & ~index[1] & ~index[2] & ~index[3] & index[7] & ~index[8] & index[9]) | (~index[0] & index[1] & index[2] & index[4] & index[8] & ~index[9] & ~index[10]) | (~index[0] & ~index[1] & index[5] & ~index[6] & index[7] & ~index[11]) | (~index[1] & index[2] & ~index[6] & ~index[7] & index[9] & ~index[11]) | (index[0] & index[1] & ~index[4] & ~index[7] & ~index[8] & ~index[9] & ~index[10]) | (index[0] & ~index[1] & ~index[3] & ~index[5] & index[7] & index[8] & ~index[10]) | (~index[0] & index[2] & index[3] & index[6] & ~index[7] & index[9] & index[10] & ~index[11]) | (index[1] & ~index[2] & index[3] & index[4] & index[7] & ~index[8] & ~index[10]) | (~index[0] & index[1] & ~index[2] & index[4] & index[8] & index[9] & ~index[11]) | (index[0] & ~index[1] & ~index[5] & index[6] & ~index[8] & ~index[9] & index[10]) | (index[1] & index[2] & ~index[3] & index[4] & index[7] & ~index[10] & ~index[11]) | (~index[0] & ~index[1] & ~index[2] & index[3] & ~index[4] & index[7] & ~index[10]) | (index[0] & index[2] & ~index[6] & ~index[7] & index[9] & ~index[11]) | (index[1] & index[2] & index[6] & index[7] & ~index[8] & ~index[10] & ~index[11]) | (index[0] & index[2] & ~index[4] & ~index[5] & ~index[6] & index[7] & index[8] & ~index[9]) | (index[0] & ~index[1] & ~index[3] & index[4] & index[6] & ~index[7] & index[10] & ~index[11]) | (~index[0] & ~index[1] & index[3] & index[4] & index[6] & index[10] & ~index[11]) | (~index[2] & ~index[5] & index[6] & index[7] & index[8] & index[9] & ~index[11]) | (index[0] & ~index[1] & ~index[4] & ~index[5] & index[6] & ~index[8] & index[10]) | (index[0] & ~index[2] & index[3] & ~index[4] & ~index[6] & ~index[7] & index[10]) | (~index[2] & index[4] & index[6] & index[8] & index[9] & ~index[10]) | (index[0] & ~index[2] & index[6] & index[7] & ~index[8] & ~index[9] & index[10]) | (index[0] & ~index[1] & ~index[2] & ~index[3] & index[4] & index[6] & ~index[8]) | (~index[1] & ~index[3] & ~index[4] & index[7] & ~index[8] & index[9] & ~index[10]) | (~index[1] & index[2] & ~index[4] & ~index[6] & index[7] & ~index[8] & ~index[11]) | (~index[0] & index[2] & ~index[3] & ~index[5] & index[6] & ~index[9] & ~index[10] & ~index[11]) | (index[1] & index[4] & index[6] & ~index[8] & index[9] & ~index[10]) | (~index[0] & index[1] & index[2] & index[4] & index[6] & ~index[7] & ~index[11]) | (~index[1] & index[2] & index[3] & index[4] & ~index[6] & index[7] & index[9]) | (~index[0] & ~index[1] & ~index[2] & index[3] & ~index[8] & ~index[9] & ~index[10]) | (index[0] & index[3] & index[4] & index[7] & index[9] & index[10] & ~index[11]) | (~index[0] & index[1] & ~index[2] & index[4] & index[6] & index[7] & ~index[9]) | (~index[0] & index[1] & index[3] & ~index[5] & ~index[6] & ~index[8] & index[10]) | (index[0] & ~index[1] & ~index[3] & ~index[5] & ~index[8] & ~index[9] & index[10]) | (~index[0] & index[1] & ~index[3] & ~index[6] & ~index[7] & index[9] & index[11]) | (~index[0] & index[2] & ~index[3] & index[5] & index[6] & index[10]) | (~index[1] & ~index[2] & ~index[3] & ~index[5] & ~index[6] & index[8] & ~index[9] & ~index[10]) | (index[2] & index[3] & ~index[5] & ~index[6] & index[7] & ~index[8] & index[10]) | (~index[1] & index[3] & ~index[4] & ~index[8] & ~index[9] & ~index[10] & ~index[11]) | (~index[0] & index[2] & ~index[3] & ~index[6] & ~index[8] & ~index[9] & index[11]) | (~index[0] & index[1] & ~index[2] & ~index[4] & ~index[5] & ~index[7] & ~index[8]) | (index[0] & ~index[2] & index[4] & ~index[8] & index[9] & index[11]) | (index[1] & ~index[2] & ~index[4] & ~index[5] & ~index[6] & ~index[7] & index[11]) | (~index[0] & index[1] & ~index[3] & ~index[5] & ~index[6] & index[7] & index[9] & ~index[11]) | (~index[2] & index[4] & index[7] & index[8] & ~index[9] & index[11]) | (~index[0] & index[1] & ~index[2] & ~index[3] & ~index[4] & ~index[9] & index[11]) | (index[0] & index[2] & ~index[6] & index[7] & index[10] & index[11]) | (index[0] & ~index[1] & index[2] & ~index[3] & index[4] & ~index[5] & ~index[7] & index[8]) | (index[0] & ~index[1] & index[2] & index[4] & ~index[7] & ~index[11]) | (index[0] & ~index[1] & ~index[3] & index[6] & index[7] & ~index[9] & index[11]) | (index[2] & index[4] & ~index[6] & index[7] & index[8] & ~index[10] & ~index[11]) | (index[1] & index[2] & index[4] & index[6] & ~index[7] & index[9] & index[11]) | (~index[0] & ~index[1] & index[3] & ~index[5] & index[8] & ~index[9] & index[10]) | (~index[0] & ~index[1] & ~index[2] & ~index[3] & index[5] & index[7] & ~index[11]) | (index[0] & ~index[2] & ~index[4] & ~index[6] & ~index[7] & index[8] & index[10]) | (~index[1] & index[2] & index[3] & ~index[4] & ~index[7] & index[9] & ~index[11]) | (~index[0] & ~index[1] & ~index[2] & ~index[4] & ~index[5] & index[8] & ~index[10] & ~index[11]) | (index[0] & index[2] & index[3] & index[7] & ~index[8] & index[11]) | (index[1] & index[2] & index[3] & ~index[4] & index[7] & index[9] & ~index[10]) | (~index[0] & ~index[3] & index[4] & index[5] & ~index[7]) | (~index[1] & index[5] & ~index[7] & index[8] & index[9] & ~index[11]) | (~index[0] & index[1] & ~index[2] & ~index[3] & ~index[5] & index[6] & index[7] & ~index[11]) | (index[0] & ~index[2] & index[3] & index[6] & index[7] & index[8] & ~index[10]) | (~index[0] & ~index[1] & index[3] & index[4] & ~index[6] & ~index[8] & index[9]) | (~index[0] & index[2] & index[3] & index[4] & ~index[6] & index[8] & ~index[11]) | (index[0] & ~index[1] & ~index[3] & ~index[4] & ~index[5] & index[7] & index[9]) | (index[0] & ~index[2] & index[3] & index[4] & index[6] & ~index[7] & index[8] & index[9]) | (~index[0] & ~index[2] & ~index[3] & ~index[5] & ~index[6] & index[10] & ~index[11]) | (~index[0] & index[3] & ~index[7] & ~index[8] & index[9] & index[10]) | (index[0] & index[1] & index[3] & index[6] & index[7] & index[8] & ~index[10]) | (index[0] & index[2] & ~index[3] & ~index[4] & index[8] & ~index[10] & index[11]) | (index[1] & index[3] & index[4] & index[8] & ~index[10] & index[11]) | (index[0] & ~index[1] & ~index[4] & ~index[6] & index[8] & index[11]) | (~index[0] & index[1] & ~index[2] & ~index[5] & ~index[6] & index[7] & index[9]) | (index[1] & index[2] & index[4] & ~index[6] & ~index[8] & ~index[9]) | (index[2] & index[3] & index[4] & ~index[8] & index[9] & index[10]) | (index[1] & index[2] & ~index[3] & index[4] & ~index[7] & index[11]) | (index[0] & ~index[2] & ~index[3] & index[6] & ~index[7] & ~index[8] & index[9]) | (index[0] & index[1] & ~index[2] & ~index[3] & ~index[4] & ~index[7] & ~index[8]) | (~index[1] & index[2] & ~index[6] & index[8] & ~index[9] & index[10]) | (~index[0] & index[1] & ~index[3] & index[4] & ~index[8] & ~index[9] & ~index[11]) | (~index[1] & index[2] & ~index[4] & index[5] & ~index[7] & index[11]) | (~index[1] & index[2] & ~index[4] & ~index[5] & ~index[6] & index[8] & index[11]) | (index[0] & ~index[1] & index[4] & index[7] & ~index[8] & index[10]) | (~index[0] & index[2] & ~index[6] & index[7] & ~index[9] & index[10]) | (index[0] & index[5] & index[6] & index[7] & ~index[8] & index[10]) | (index[0] & ~index[1] & index[2] & ~index[4] & index[7] & index[10] & ~index[11]) | (index[0] & index[2] & ~index[3] & index[4] & ~index[7] & ~index[9] & index[10]);

assign val[7] = 0;



endmodule
