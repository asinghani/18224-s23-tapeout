module d01_example_adder (
	io_in,
	io_out
);
	wire _00_;
	wire _01_;
	wire _02_;
	wire _03_;
	wire _04_;
	wire _05_;
	wire _06_;
	wire _07_;
	wire _08_;
	wire _09_;
	wire _10_;
	wire _11_;
	wire _12_;
	wire _13_;
	wire _14_;
	wire _15_;
	wire _16_;
	wire _17_;
	wire _18_;
	wire _19_;
	wire _20_;
	wire _21_;
	wire _22_;
	wire _23_;
	wire _24_;
	wire _25_;
	input wire [13:0] io_in;
	output wire [13:0] io_out;
	wire \mchip.clock ;
	wire [11:0] \mchip.io_in ;
	wire [11:0] \mchip.io_out ;
	wire \mchip.reset ;
	assign _00_ = io_in[11] ^ io_in[5];
	assign _01_ = ~(io_in[10] ^ io_in[4]);
	assign _02_ = _00_ & ~_01_;
	assign _03_ = ~(io_in[9] & io_in[3]);
	assign _04_ = io_in[9] ^ io_in[3];
	assign _05_ = ~(io_in[8] & io_in[2]);
	assign _06_ = _04_ & ~_05_;
	assign _07_ = _03_ & ~_06_;
	assign _08_ = ~(io_in[8] ^ io_in[2]);
	assign _09_ = _04_ & ~_08_;
	assign _10_ = ~(io_in[7] & io_in[1]);
	assign _11_ = io_in[7] ^ io_in[1];
	assign _12_ = ~(io_in[6] & io_in[0]);
	assign _13_ = _11_ & ~_12_;
	assign _14_ = _10_ & ~_13_;
	assign _15_ = _09_ & ~_14_;
	assign _16_ = _07_ & ~_15_;
	assign _17_ = _02_ & ~_16_;
	assign _18_ = ~(io_in[10] & io_in[4]);
	assign _19_ = _00_ & ~_18_;
	assign _20_ = io_in[11] & io_in[5];
	assign _21_ = _20_ | _19_;
	assign io_out[6] = _21_ | _17_;
	assign io_out[1] = ~(_12_ ^ _11_);
	assign io_out[2] = _14_ ^ _08_;
	assign _22_ = ~(_14_ | _08_);
	assign _23_ = _22_ | ~_05_;
	assign io_out[3] = _23_ ^ _04_;
	assign io_out[4] = _16_ ^ _01_;
	assign _24_ = ~(_16_ | _01_);
	assign _25_ = _24_ | ~_18_;
	assign io_out[5] = _25_ ^ _00_;
	assign io_out[0] = io_in[6] ^ io_in[0];
	assign io_out[13:7] = 7'h00;
	assign \mchip.clock  = io_in[12];
	assign \mchip.io_in  = io_in[11:0];
	assign \mchip.io_out  = {5'h00, io_out[6:0]};
	assign \mchip.reset  = io_in[13];
endmodule
module d02_example_counter (
	io_in,
	io_out
);
	wire _000_;
	wire _001_;
	wire _002_;
	wire _003_;
	wire _004_;
	wire _005_;
	wire _006_;
	wire _007_;
	wire _008_;
	wire _009_;
	wire _010_;
	wire _011_;
	wire _012_;
	wire _013_;
	wire _014_;
	wire _015_;
	wire _016_;
	wire _017_;
	wire _018_;
	wire _019_;
	wire _020_;
	wire _021_;
	wire _022_;
	wire _023_;
	wire _024_;
	wire _025_;
	wire _026_;
	wire _027_;
	wire _028_;
	wire _029_;
	wire _030_;
	wire _031_;
	wire _032_;
	wire _033_;
	wire _034_;
	wire _035_;
	wire _036_;
	wire _037_;
	wire _038_;
	wire _039_;
	wire _040_;
	wire _041_;
	wire _042_;
	wire _043_;
	wire _044_;
	wire _045_;
	wire _046_;
	wire _047_;
	wire _048_;
	wire _049_;
	wire _050_;
	wire _051_;
	wire _052_;
	wire _053_;
	wire _054_;
	wire _055_;
	wire _056_;
	wire _057_;
	wire _058_;
	wire [11:0] _059_;
	input wire [13:0] io_in;
	output wire [13:0] io_out;
	wire \mchip.clock ;
	wire \mchip.enable ;
	wire [11:0] \mchip.io_in ;
	reg [11:0] \mchip.io_out ;
	wire \mchip.reset ;
	wire \mchip.updown ;
	assign _059_[0] = ~\mchip.io_out [0];
	assign _001_ = ~(io_in[1] & io_in[0]);
	assign _002_ = io_in[1] | ~io_in[0];
	assign _000_ = ~(_002_ & _001_);
	assign _003_ = _001_ ^ \mchip.io_out [1];
	assign _059_[1] = _003_ ^ _059_[0];
	assign _004_ = \mchip.io_out [1] & ~_001_;
	assign _005_ = \mchip.io_out [0] & ~_003_;
	assign _006_ = _005_ | _004_;
	assign _007_ = _001_ ^ \mchip.io_out [2];
	assign _059_[2] = ~(_007_ ^ _006_);
	assign _008_ = \mchip.io_out [2] & ~_001_;
	assign _009_ = _006_ & ~_007_;
	assign _010_ = ~(_009_ | _008_);
	assign _011_ = _001_ ^ \mchip.io_out [3];
	assign _059_[3] = _011_ ^ _010_;
	assign _012_ = _011_ | _007_;
	assign _013_ = _006_ & ~_012_;
	assign _014_ = \mchip.io_out [3] & ~_001_;
	assign _015_ = _008_ & ~_011_;
	assign _016_ = _015_ | _014_;
	assign _017_ = _016_ | _013_;
	assign _018_ = _001_ ^ \mchip.io_out [4];
	assign _059_[4] = ~(_018_ ^ _017_);
	assign _019_ = \mchip.io_out [4] & ~_001_;
	assign _020_ = _017_ & ~_018_;
	assign _021_ = ~(_020_ | _019_);
	assign _022_ = _001_ ^ \mchip.io_out [5];
	assign _059_[5] = _022_ ^ _021_;
	assign _023_ = _022_ | _018_;
	assign _024_ = _017_ & ~_023_;
	assign _025_ = \mchip.io_out [5] & ~_001_;
	assign _026_ = _019_ & ~_022_;
	assign _027_ = _026_ | _025_;
	assign _028_ = _027_ | _024_;
	assign _029_ = _001_ ^ \mchip.io_out [6];
	assign _059_[6] = ~(_029_ ^ _028_);
	assign _030_ = \mchip.io_out [6] & ~_001_;
	assign _031_ = _028_ & ~_029_;
	assign _032_ = ~(_031_ | _030_);
	assign _033_ = _001_ ^ \mchip.io_out [7];
	assign _059_[7] = _033_ ^ _032_;
	assign _034_ = \mchip.io_out [7] & ~_001_;
	assign _035_ = _030_ & ~_033_;
	assign _036_ = _035_ | _034_;
	assign _037_ = _033_ | _029_;
	assign _038_ = _027_ & ~_037_;
	assign _039_ = _038_ | _036_;
	assign _040_ = _037_ | _023_;
	assign _041_ = _017_ & ~_040_;
	assign _042_ = _041_ | _039_;
	assign _043_ = ~(_001_ ^ \mchip.io_out [8]);
	assign _059_[8] = _043_ ^ _042_;
	assign _044_ = \mchip.io_out [8] & ~_001_;
	assign _045_ = _043_ & _042_;
	assign _046_ = _045_ | _044_;
	assign _047_ = ~(_001_ ^ \mchip.io_out [9]);
	assign _059_[9] = _047_ ^ _046_;
	assign _048_ = \mchip.io_out [9] & ~_001_;
	assign _049_ = _047_ & _044_;
	assign _050_ = _049_ | _048_;
	assign _051_ = ~(_047_ & _043_);
	assign _052_ = _042_ & ~_051_;
	assign _053_ = _052_ | _050_;
	assign _054_ = ~(_001_ ^ \mchip.io_out [10]);
	assign _059_[10] = _054_ ^ _053_;
	assign _055_ = \mchip.io_out [10] & ~_001_;
	assign _056_ = _054_ & _053_;
	assign _057_ = _056_ | _055_;
	assign _058_ = ~(_001_ ^ \mchip.io_out [11]);
	assign _059_[11] = _058_ ^ _057_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.io_out [0] <= 1'h0;
		else if (_000_)
			\mchip.io_out [0] <= _059_[0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.io_out [1] <= 1'h0;
		else if (_000_)
			\mchip.io_out [1] <= _059_[1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.io_out [2] <= 1'h0;
		else if (_000_)
			\mchip.io_out [2] <= _059_[2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.io_out [3] <= 1'h0;
		else if (_000_)
			\mchip.io_out [3] <= _059_[3];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.io_out [4] <= 1'h0;
		else if (_000_)
			\mchip.io_out [4] <= _059_[4];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.io_out [5] <= 1'h0;
		else if (_000_)
			\mchip.io_out [5] <= _059_[5];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.io_out [6] <= 1'h0;
		else if (_000_)
			\mchip.io_out [6] <= _059_[6];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.io_out [7] <= 1'h0;
		else if (_000_)
			\mchip.io_out [7] <= _059_[7];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.io_out [8] <= 1'h0;
		else if (_000_)
			\mchip.io_out [8] <= _059_[8];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.io_out [9] <= 1'h0;
		else if (_000_)
			\mchip.io_out [9] <= _059_[9];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.io_out [10] <= 1'h0;
		else if (_000_)
			\mchip.io_out [10] <= _059_[10];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.io_out [11] <= 1'h0;
		else if (_000_)
			\mchip.io_out [11] <= _059_[11];
	assign io_out = {2'h0, \mchip.io_out };
	assign \mchip.clock  = io_in[12];
	assign \mchip.enable  = io_in[0];
	assign \mchip.io_in  = io_in[11:0];
	assign \mchip.reset  = io_in[13];
	assign \mchip.updown  = io_in[1];
endmodule
module d03_example_beepboop (
	io_in,
	io_out
);
	wire _000_;
	wire _001_;
	wire _002_;
	wire _003_;
	wire _004_;
	wire _005_;
	wire _006_;
	wire _007_;
	wire _008_;
	wire _009_;
	wire _010_;
	wire _011_;
	wire _012_;
	wire _013_;
	wire _014_;
	wire _015_;
	wire _016_;
	wire _017_;
	wire _018_;
	wire _019_;
	wire _020_;
	wire _021_;
	wire _022_;
	wire _023_;
	wire _024_;
	wire _025_;
	wire _026_;
	wire _027_;
	wire _028_;
	wire _029_;
	wire _030_;
	wire _031_;
	wire _032_;
	wire _033_;
	wire _034_;
	wire _035_;
	wire _036_;
	wire _037_;
	wire _038_;
	wire _039_;
	wire _040_;
	wire _041_;
	wire _042_;
	wire _043_;
	wire _044_;
	wire _045_;
	wire _046_;
	wire _047_;
	wire _048_;
	wire _049_;
	wire _050_;
	wire _051_;
	wire _052_;
	wire _053_;
	wire _054_;
	wire _055_;
	wire _056_;
	wire _057_;
	wire _058_;
	wire _059_;
	wire _060_;
	wire _061_;
	wire _062_;
	wire _063_;
	wire _064_;
	wire _065_;
	wire _066_;
	wire _067_;
	wire _068_;
	wire _069_;
	wire _070_;
	wire _071_;
	wire _072_;
	wire _073_;
	wire _074_;
	wire _075_;
	wire _076_;
	wire _077_;
	wire _078_;
	wire _079_;
	wire _080_;
	wire _081_;
	wire _082_;
	wire _083_;
	wire _084_;
	wire _085_;
	wire _086_;
	wire _087_;
	wire _088_;
	wire _089_;
	wire _090_;
	wire _091_;
	wire _092_;
	wire _093_;
	wire _094_;
	wire _095_;
	wire _096_;
	wire _097_;
	wire _098_;
	wire _099_;
	wire _100_;
	wire _101_;
	wire _102_;
	wire _103_;
	wire _104_;
	wire _105_;
	wire _106_;
	wire _107_;
	wire _108_;
	wire _109_;
	wire _110_;
	wire _111_;
	wire _112_;
	wire _113_;
	wire _114_;
	wire _115_;
	wire _116_;
	wire _117_;
	wire _118_;
	wire _119_;
	wire _120_;
	wire _121_;
	wire _122_;
	wire _123_;
	wire _124_;
	wire _125_;
	wire _126_;
	wire _127_;
	wire _128_;
	wire _129_;
	wire _130_;
	wire _131_;
	wire _132_;
	wire _133_;
	wire _134_;
	wire _135_;
	wire _136_;
	wire _137_;
	wire _138_;
	wire _139_;
	wire _140_;
	wire _141_;
	wire _142_;
	wire _143_;
	wire _144_;
	wire _145_;
	wire _146_;
	wire _147_;
	wire _148_;
	wire _149_;
	wire _150_;
	wire _151_;
	wire _152_;
	wire _153_;
	wire _154_;
	wire _155_;
	wire _156_;
	wire _157_;
	wire _158_;
	wire _159_;
	wire _160_;
	wire _161_;
	wire _162_;
	wire _163_;
	wire _164_;
	wire _165_;
	wire _166_;
	wire _167_;
	wire _168_;
	wire _169_;
	wire _170_;
	wire _171_;
	wire _172_;
	wire _173_;
	wire _174_;
	wire _175_;
	wire _176_;
	wire _177_;
	wire _178_;
	wire _179_;
	wire _180_;
	wire _181_;
	wire _182_;
	wire _183_;
	wire _184_;
	wire _185_;
	wire _186_;
	wire _187_;
	wire _188_;
	wire _189_;
	wire _190_;
	wire _191_;
	wire _192_;
	wire _193_;
	wire _194_;
	wire _195_;
	wire _196_;
	wire _197_;
	wire _198_;
	wire _199_;
	wire _200_;
	wire _201_;
	wire _202_;
	wire _203_;
	wire _204_;
	wire _205_;
	wire _206_;
	wire _207_;
	wire _208_;
	wire _209_;
	wire _210_;
	wire _211_;
	wire _212_;
	wire _213_;
	wire _214_;
	wire _215_;
	wire _216_;
	wire _217_;
	wire _218_;
	wire _219_;
	wire _220_;
	wire _221_;
	wire _222_;
	wire _223_;
	wire _224_;
	wire _225_;
	wire _226_;
	wire _227_;
	wire _228_;
	wire _229_;
	wire _230_;
	wire _231_;
	wire _232_;
	wire _233_;
	wire _234_;
	wire _235_;
	wire _236_;
	wire _237_;
	wire _238_;
	wire _239_;
	wire _240_;
	wire _241_;
	wire _242_;
	wire _243_;
	wire _244_;
	wire _245_;
	wire _246_;
	wire _247_;
	wire _248_;
	wire _249_;
	wire _250_;
	wire _251_;
	wire _252_;
	wire _253_;
	wire _254_;
	wire _255_;
	wire _256_;
	wire _257_;
	wire _258_;
	wire _259_;
	wire _260_;
	wire _261_;
	wire _262_;
	wire _263_;
	wire _264_;
	wire [15:0] _265_;
	input wire [13:0] io_in;
	output wire [13:0] io_out;
	wire [0:191] \mchip.beepboop ;
	wire \mchip.btn ;
	wire \mchip.chr_out ;
	wire \mchip.chr_out_valid ;
	wire \mchip.clock ;
	reg [15:0] \mchip.counter ;
	wire \mchip.green ;
	wire [11:0] \mchip.io_in ;
	wire [11:0] \mchip.io_out ;
	wire \mchip.no_walk ;
	wire \mchip.red ;
	wire \mchip.reset ;
	wire \mchip.the_beepbooper ;
	wire \mchip.walk ;
	wire \mchip.yellow ;
	assign _215_ = ~(\mchip.counter [15] | \mchip.counter [14]);
	assign _216_ = \mchip.counter [12] | \mchip.counter [13];
	assign _217_ = _215_ & ~_216_;
	assign _218_ = \mchip.counter [10] | \mchip.counter [11];
	assign _219_ = ~(\mchip.counter [8] | \mchip.counter [9]);
	assign _220_ = _219_ & ~_218_;
	assign _221_ = ~(_220_ & _217_);
	assign _222_ = \mchip.counter [6] | \mchip.counter [7];
	assign _223_ = \mchip.counter [4] | \mchip.counter [5];
	assign _116_ = ~(_223_ | _222_);
	assign _224_ = ~(\mchip.counter [2] | \mchip.counter [3]);
	assign _225_ = \mchip.counter [0] | \mchip.counter [1];
	assign _108_ = _224_ & ~_225_;
	assign _226_ = ~(_108_ & _116_);
	assign _002_ = _226_ | _221_;
	assign _227_ = io_in[0] & ~_002_;
	assign _228_ = \mchip.counter [11] & ~\mchip.counter [10];
	assign _229_ = ~(_228_ & _219_);
	assign _230_ = _217_ & ~_229_;
	assign _231_ = \mchip.counter [2] | ~\mchip.counter [3];
	assign _232_ = _231_ | _225_;
	assign _233_ = \mchip.counter [6] | ~\mchip.counter [7];
	assign _234_ = \mchip.counter [5] | ~\mchip.counter [4];
	assign _235_ = ~(_234_ | _233_);
	assign _236_ = _232_ | ~_235_;
	assign _237_ = _230_ & ~_236_;
	assign _238_ = _237_ | _227_;
	assign _239_ = \mchip.counter [11] | ~_217_;
	assign _240_ = ~(_233_ | _223_);
	assign _241_ = \mchip.counter [7] & ~_240_;
	assign _242_ = _232_ & \mchip.counter [3];
	assign _243_ = _235_ & ~_242_;
	assign _244_ = _241_ & ~_243_;
	assign _245_ = _230_ & ~_244_;
	assign _246_ = _239_ & ~_245_;
	assign _247_ = _246_ | io_in[13];
	assign _001_ = _247_ | _238_;
	assign _248_ = _246_ | _237_;
	assign _249_ = _248_ | _227_;
	assign _000_ = _249_ | _002_;
	assign _250_ = \mchip.counter [9] | ~\mchip.counter [8];
	assign _251_ = _250_ | _218_;
	assign _252_ = _217_ & ~_251_;
	assign _253_ = _222_ | \mchip.counter [5];
	assign _254_ = \mchip.counter [4] | ~\mchip.counter [5];
	assign _255_ = ~(_254_ | _222_);
	assign _256_ = ~(\mchip.counter [2] & \mchip.counter [3]);
	assign _257_ = _225_ & ~_256_;
	assign _258_ = _255_ & ~_257_;
	assign _259_ = _253_ & ~_258_;
	assign _260_ = _252_ & ~_259_;
	assign _261_ = _221_ & ~_260_;
	assign _262_ = _256_ | _225_;
	assign _263_ = _262_ | ~_255_;
	assign _264_ = _263_ | ~_252_;
	assign _004_ = ~(_264_ & _261_);
	assign _005_ = \mchip.counter [4] & \mchip.counter [5];
	assign _006_ = _005_ & ~_222_;
	assign _007_ = \mchip.counter [3] | ~\mchip.counter [2];
	assign _008_ = ~(_007_ | _225_);
	assign _009_ = ~(_008_ & _006_);
	assign _010_ = _230_ & ~_009_;
	assign _011_ = _005_ | _222_;
	assign _012_ = \mchip.counter [2] | \mchip.counter [3];
	assign _013_ = _012_ & ~_008_;
	assign _014_ = _006_ & ~_013_;
	assign _015_ = _011_ & ~_014_;
	assign _016_ = _230_ & ~_015_;
	assign _017_ = _239_ & ~_016_;
	assign _018_ = _017_ | _010_;
	assign _019_ = ~(\mchip.counter [8] & \mchip.counter [9]);
	assign _020_ = \mchip.counter [11] | ~\mchip.counter [10];
	assign _021_ = _020_ | _019_;
	assign _022_ = _217_ & ~_021_;
	assign _023_ = \mchip.counter [7] | ~\mchip.counter [6];
	assign _024_ = _023_ | _254_;
	assign _025_ = _024_ | _262_;
	assign _026_ = _022_ & ~_025_;
	assign _027_ = ~_217_;
	assign _028_ = _019_ & ~_020_;
	assign _029_ = _218_ & ~_028_;
	assign _030_ = _029_ | _027_;
	assign _031_ = ~\mchip.counter [5];
	assign _032_ = _031_ & ~_023_;
	assign _033_ = _222_ & ~_032_;
	assign _034_ = ~(_024_ | _257_);
	assign _035_ = _033_ & ~_034_;
	assign _036_ = _022_ & ~_035_;
	assign _037_ = _030_ & ~_036_;
	assign _038_ = _037_ | _026_;
	assign _039_ = \mchip.counter [6] & \mchip.counter [7];
	assign _040_ = _234_ | ~_039_;
	assign _041_ = _040_ | ~_108_;
	assign _042_ = _022_ & ~_041_;
	assign _043_ = ~(\mchip.counter [4] | \mchip.counter [5]);
	assign _044_ = _039_ & ~_043_;
	assign _045_ = _044_ & _041_;
	assign _046_ = _022_ & ~_045_;
	assign _047_ = _030_ & ~_046_;
	assign _048_ = _047_ | _042_;
	assign _049_ = _038_ & ~_048_;
	assign _050_ = \mchip.counter [8] | ~\mchip.counter [9];
	assign _051_ = _050_ | _020_;
	assign _052_ = _217_ & ~_051_;
	assign _053_ = _254_ | _233_;
	assign _054_ = _053_ | ~_008_;
	assign _055_ = _052_ & ~_054_;
	assign _056_ = ~(_020_ | \mchip.counter [9]);
	assign _057_ = _218_ & ~_056_;
	assign _058_ = _057_ | _027_;
	assign _059_ = _031_ & ~_233_;
	assign _060_ = \mchip.counter [7] & ~_059_;
	assign _061_ = ~(_053_ | _013_);
	assign _062_ = _060_ & ~_061_;
	assign _063_ = _052_ & ~_062_;
	assign _064_ = _058_ & ~_063_;
	assign _065_ = _064_ | _055_;
	assign _066_ = _232_ | ~_116_;
	assign _067_ = _022_ & ~_066_;
	assign _068_ = _242_ | ~_116_;
	assign _069_ = _022_ & ~_068_;
	assign _070_ = _030_ & ~_069_;
	assign _071_ = _070_ | _067_;
	assign _072_ = _065_ & ~_071_;
	assign _073_ = _023_ | _223_;
	assign _074_ = _108_ & ~_073_;
	assign _075_ = ~(_074_ & _052_);
	assign _076_ = _222_ & ~_074_;
	assign _077_ = _052_ & ~_076_;
	assign _078_ = _058_ & ~_077_;
	assign _079_ = _075_ & ~_078_;
	assign _080_ = ~(_020_ | _250_);
	assign _081_ = ~(_080_ & _217_);
	assign _082_ = _040_ | _262_;
	assign _083_ = ~(_082_ | _081_);
	assign _084_ = ~(_040_ | _257_);
	assign _085_ = _044_ & ~_084_;
	assign _086_ = _085_ | _081_;
	assign _087_ = _219_ & ~_020_;
	assign _088_ = _218_ & ~_087_;
	assign _089_ = _217_ & ~_088_;
	assign _090_ = _086_ & ~_089_;
	assign _091_ = ~(_090_ | _083_);
	assign _092_ = _079_ & ~_091_;
	assign _093_ = _092_ | _072_;
	assign _094_ = _093_ | _049_;
	assign _095_ = _094_ | _018_;
	assign \mchip.no_walk  = _095_ | _004_;
	assign \mchip.the_beepbooper  = _091_ & _261_;
	assign _096_ = ~(_039_ & _043_);
	assign _097_ = _096_ | _232_;
	assign _098_ = ~(_097_ | _221_);
	assign _099_ = ~(_096_ | _242_);
	assign _100_ = _039_ & ~_099_;
	assign _101_ = _100_ | _221_;
	assign _102_ = _101_ | _098_;
	assign \mchip.red  = _102_ & ~_248_;
	assign \mchip.yellow  = _002_ & ~_102_;
	assign \mchip.green  = _248_ | ~_002_;
	assign _103_ = _108_ & ~_096_;
	assign _104_ = _221_ | ~_103_;
	assign _105_ = _039_ & ~_103_;
	assign _106_ = ~(_105_ | _221_);
	assign _107_ = _104_ & ~_106_;
	assign \mchip.chr_out_valid  = _002_ & ~_107_;
	assign _109_ = _108_ & ~_223_;
	assign _110_ = _109_ ^ \mchip.counter [6];
	assign _111_ = ~_110_;
	assign _112_ = \mchip.counter [0] & \mchip.counter [1];
	assign _113_ = _225_ & ~_112_;
	assign _114_ = ~\mchip.counter [0];
	assign _115_ = ~\mchip.counter [8];
	assign _117_ = _116_ & ~_108_;
	assign _118_ = _117_ | ~_116_;
	assign _119_ = _118_ ^ _115_;
	assign _120_ = _109_ & ~\mchip.counter [6];
	assign _121_ = ~(_120_ ^ \mchip.counter [7]);
	assign _122_ = _110_ & ~_121_;
	assign _123_ = _122_ | _119_;
	assign _124_ = _115_ & ~_118_;
	assign _125_ = _124_ ^ \mchip.counter [9];
	assign _126_ = _125_ ^ _123_;
	assign _127_ = _126_ | _114_;
	assign _128_ = _114_ & ~_126_;
	assign _129_ = _127_ & ~_128_;
	assign _130_ = _113_ & ~_129_;
	assign _131_ = ~_113_;
	assign _132_ = _131_ & ~_129_;
	assign _133_ = ~(_132_ | _130_);
	assign _134_ = ~\mchip.counter [2];
	assign _135_ = _225_ ^ _134_;
	assign _136_ = _126_ | \mchip.counter [0];
	assign _137_ = (_113_ ? _136_ : _127_);
	assign _138_ = _134_ & ~_225_;
	assign _139_ = _138_ ^ \mchip.counter [3];
	assign _140_ = (_135_ ? _133_ : _137_);
	assign _141_ = _108_ ^ \mchip.counter [4];
	assign _142_ = ~_135_;
	assign _143_ = _136_ | _131_;
	assign _144_ = _127_ | _113_;
	assign _145_ = (_135_ ? _144_ : _143_);
	assign _146_ = _144_ | _135_;
	assign _147_ = (_139_ ? _145_ : _146_);
	assign _148_ = (_141_ ? _140_ : _147_);
	assign _149_ = _108_ & ~\mchip.counter [4];
	assign _150_ = _149_ ^ \mchip.counter [5];
	assign _151_ = (_113_ ? _136_ : _129_);
	assign _152_ = _151_ | _135_;
	assign _153_ = (_135_ ? _136_ : _137_);
	assign _154_ = (_139_ ? _152_ : _153_);
	assign _155_ = (_139_ ? _153_ : _145_);
	assign _156_ = (_141_ ? _154_ : _155_);
	assign _157_ = (_150_ ? _148_ : _156_);
	assign _158_ = _111_ & ~_157_;
	assign _159_ = _121_ ^ _110_;
	assign _160_ = (_135_ ? _143_ : _151_);
	assign _161_ = ~(_160_ | _139_);
	assign _162_ = \mchip.counter [0] & ~_126_;
	assign _163_ = (_113_ ? _128_ : _162_);
	assign _164_ = _113_ & ~_127_;
	assign _165_ = (_135_ ? _164_ : _163_);
	assign _166_ = ~(_136_ & _127_);
	assign _167_ = (_113_ ? _128_ : _166_);
	assign _168_ = (_135_ ? _167_ : _163_);
	assign _169_ = (_139_ ? _165_ : _168_);
	assign _170_ = (_141_ ? _161_ : _169_);
	assign _171_ = (_113_ ? _162_ : _128_);
	assign _172_ = (_135_ ? _171_ : _163_);
	assign _173_ = _113_ & ~_136_;
	assign _174_ = (_135_ ? _130_ : _173_);
	assign _175_ = (_139_ ? _172_ : _174_);
	assign _176_ = _142_ & ~_144_;
	assign _177_ = (_135_ ? _132_ : _163_);
	assign _178_ = (_139_ ? _176_ : _177_);
	assign _179_ = (_141_ ? _175_ : _178_);
	assign _180_ = (_150_ ? _170_ : _179_);
	assign _181_ = (_139_ ? _172_ : _163_);
	assign _182_ = _131_ & ~_136_;
	assign _183_ = (_135_ ? _182_ : _163_);
	assign _184_ = (_139_ ? _163_ : _183_);
	assign _185_ = (_141_ ? _181_ : _184_);
	assign _186_ = _131_ & ~_127_;
	assign _187_ = (_135_ ? _186_ : _167_);
	assign _188_ = (_135_ ? _173_ : _128_);
	assign _189_ = (_139_ ? _187_ : _188_);
	assign _190_ = _142_ & ~_151_;
	assign _191_ = (_139_ ? _176_ : _190_);
	assign _192_ = (_141_ ? _189_ : _191_);
	assign _193_ = (_150_ ? _185_ : _192_);
	assign _194_ = (_110_ ? _193_ : _180_);
	assign _195_ = (_159_ ? _158_ : _194_);
	assign _196_ = _122_ ^ _119_;
	assign \mchip.chr_out  = _195_ & ~_196_;
	assign _265_[1] = \mchip.counter [0] ^ \mchip.counter [1];
	assign _265_[2] = _112_ ^ \mchip.counter [2];
	assign _197_ = _112_ & ~_134_;
	assign _265_[3] = _197_ ^ \mchip.counter [3];
	assign _198_ = _112_ & ~_256_;
	assign _265_[4] = _198_ ^ \mchip.counter [4];
	assign _199_ = _198_ & \mchip.counter [4];
	assign _265_[5] = _199_ ^ \mchip.counter [5];
	assign _200_ = _198_ & _005_;
	assign _265_[6] = _200_ ^ \mchip.counter [6];
	assign _201_ = _200_ & \mchip.counter [6];
	assign _265_[7] = _201_ ^ \mchip.counter [7];
	assign _202_ = _039_ & _005_;
	assign _203_ = ~(_202_ & _198_);
	assign _265_[8] = _203_ ^ _115_;
	assign _204_ = \mchip.counter [8] & ~_203_;
	assign _265_[9] = _204_ ^ \mchip.counter [9];
	assign _205_ = ~(_203_ | _019_);
	assign _265_[10] = _205_ ^ \mchip.counter [10];
	assign _206_ = _205_ & \mchip.counter [10];
	assign _265_[11] = _206_ ^ \mchip.counter [11];
	assign _207_ = ~(\mchip.counter [10] & \mchip.counter [11]);
	assign _208_ = _207_ | _019_;
	assign _209_ = ~(_208_ | _203_);
	assign _265_[12] = _209_ ^ \mchip.counter [12];
	assign _210_ = _209_ & \mchip.counter [12];
	assign _265_[13] = _210_ ^ \mchip.counter [13];
	assign _211_ = ~(\mchip.counter [12] & \mchip.counter [13]);
	assign _212_ = _209_ & ~_211_;
	assign _265_[14] = _212_ ^ \mchip.counter [14];
	assign _213_ = _212_ & \mchip.counter [14];
	assign _265_[15] = _213_ ^ \mchip.counter [15];
	assign _214_ = _114_ & ~_248_;
	assign _003_ = _214_ | _227_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.counter [0] <= 1'h0;
		else if (_000_)
			\mchip.counter [0] <= _003_;
	always @(posedge io_in[12])
		if (_001_)
			\mchip.counter [1] <= 1'h0;
		else if (_002_)
			\mchip.counter [1] <= _265_[1];
	always @(posedge io_in[12])
		if (_001_)
			\mchip.counter [2] <= 1'h0;
		else if (_002_)
			\mchip.counter [2] <= _265_[2];
	always @(posedge io_in[12])
		if (_001_)
			\mchip.counter [3] <= 1'h0;
		else if (_002_)
			\mchip.counter [3] <= _265_[3];
	always @(posedge io_in[12])
		if (_001_)
			\mchip.counter [4] <= 1'h0;
		else if (_002_)
			\mchip.counter [4] <= _265_[4];
	always @(posedge io_in[12])
		if (_001_)
			\mchip.counter [5] <= 1'h0;
		else if (_002_)
			\mchip.counter [5] <= _265_[5];
	always @(posedge io_in[12])
		if (_001_)
			\mchip.counter [6] <= 1'h0;
		else if (_002_)
			\mchip.counter [6] <= _265_[6];
	always @(posedge io_in[12])
		if (_001_)
			\mchip.counter [7] <= 1'h0;
		else if (_002_)
			\mchip.counter [7] <= _265_[7];
	always @(posedge io_in[12])
		if (_001_)
			\mchip.counter [8] <= 1'h0;
		else if (_002_)
			\mchip.counter [8] <= _265_[8];
	always @(posedge io_in[12])
		if (_001_)
			\mchip.counter [9] <= 1'h0;
		else if (_002_)
			\mchip.counter [9] <= _265_[9];
	always @(posedge io_in[12])
		if (_001_)
			\mchip.counter [10] <= 1'h0;
		else if (_002_)
			\mchip.counter [10] <= _265_[10];
	always @(posedge io_in[12])
		if (_001_)
			\mchip.counter [11] <= 1'h0;
		else if (_002_)
			\mchip.counter [11] <= _265_[11];
	always @(posedge io_in[12])
		if (_001_)
			\mchip.counter [12] <= 1'h0;
		else if (_002_)
			\mchip.counter [12] <= _265_[12];
	always @(posedge io_in[12])
		if (_001_)
			\mchip.counter [13] <= 1'h0;
		else if (_002_)
			\mchip.counter [13] <= _265_[13];
	always @(posedge io_in[12])
		if (_001_)
			\mchip.counter [14] <= 1'h0;
		else if (_002_)
			\mchip.counter [14] <= _265_[14];
	always @(posedge io_in[12])
		if (_001_)
			\mchip.counter [15] <= 1'h0;
		else if (_002_)
			\mchip.counter [15] <= _265_[15];
	assign _265_[0] = 1'h0;
	assign io_out = {6'h00, \mchip.chr_out_valid , \mchip.chr_out , \mchip.the_beepbooper , \mchip.no_walk , \mchip.the_beepbooper , \mchip.green , \mchip.yellow , \mchip.red };
	assign \mchip.beepboop  = 192'h4265657020426f6f702054726166666963204c6967687400;
	assign \mchip.btn  = io_in[0];
	assign \mchip.clock  = io_in[12];
	assign \mchip.io_in  = io_in[11:0];
	assign \mchip.io_out  = {4'h0, \mchip.chr_out_valid , \mchip.chr_out , \mchip.the_beepbooper , \mchip.no_walk , \mchip.the_beepbooper , \mchip.green , \mchip.yellow , \mchip.red };
	assign \mchip.reset  = io_in[13];
	assign \mchip.walk  = \mchip.the_beepbooper ;
endmodule
module d04_example_aes128sca (
	io_in,
	io_out
);
	wire _0000_;
	wire _0001_;
	wire _0002_;
	wire _0003_;
	wire _0004_;
	wire _0005_;
	wire _0006_;
	wire _0007_;
	wire _0008_;
	wire _0009_;
	wire _0010_;
	wire _0011_;
	wire _0012_;
	wire _0013_;
	wire _0014_;
	wire _0015_;
	wire _0016_;
	wire _0017_;
	wire _0018_;
	wire _0019_;
	wire _0020_;
	wire _0021_;
	wire _0022_;
	wire _0023_;
	wire _0024_;
	wire _0025_;
	wire _0026_;
	wire _0027_;
	wire _0028_;
	wire _0029_;
	wire _0030_;
	wire _0031_;
	wire _0032_;
	wire _0033_;
	wire _0034_;
	wire _0035_;
	wire _0036_;
	wire _0037_;
	wire _0038_;
	wire _0039_;
	wire _0040_;
	wire _0041_;
	wire _0042_;
	wire _0043_;
	wire _0044_;
	wire _0045_;
	wire _0046_;
	wire _0047_;
	wire _0048_;
	wire _0049_;
	wire _0050_;
	wire _0051_;
	wire _0052_;
	wire _0053_;
	wire _0054_;
	wire _0055_;
	wire _0056_;
	wire _0057_;
	wire _0058_;
	wire _0059_;
	wire _0060_;
	wire _0061_;
	wire _0062_;
	wire _0063_;
	wire _0064_;
	wire _0065_;
	wire _0066_;
	wire _0067_;
	wire _0068_;
	wire _0069_;
	wire _0070_;
	wire _0071_;
	wire _0072_;
	wire _0073_;
	wire _0074_;
	wire _0075_;
	wire _0076_;
	wire _0077_;
	wire _0078_;
	wire _0079_;
	wire _0080_;
	wire _0081_;
	wire _0082_;
	wire _0083_;
	wire _0084_;
	wire _0085_;
	wire _0086_;
	wire _0087_;
	wire _0088_;
	wire _0089_;
	wire _0090_;
	wire _0091_;
	wire _0092_;
	wire _0093_;
	wire _0094_;
	wire _0095_;
	wire _0096_;
	wire _0097_;
	wire _0098_;
	wire _0099_;
	wire _0100_;
	wire _0101_;
	wire _0102_;
	wire _0103_;
	wire _0104_;
	wire _0105_;
	wire _0106_;
	wire _0107_;
	wire _0108_;
	wire _0109_;
	wire _0110_;
	wire _0111_;
	wire _0112_;
	wire _0113_;
	wire _0114_;
	wire _0115_;
	wire _0116_;
	wire _0117_;
	wire _0118_;
	wire _0119_;
	wire _0120_;
	wire _0121_;
	wire _0122_;
	wire _0123_;
	wire _0124_;
	wire _0125_;
	wire _0126_;
	wire _0127_;
	wire _0128_;
	wire _0129_;
	wire _0130_;
	wire _0131_;
	wire _0132_;
	wire _0133_;
	wire _0134_;
	wire _0135_;
	wire _0136_;
	wire _0137_;
	wire _0138_;
	wire _0139_;
	wire _0140_;
	wire _0141_;
	wire _0142_;
	wire _0143_;
	wire _0144_;
	wire _0145_;
	wire _0146_;
	wire _0147_;
	wire _0148_;
	wire _0149_;
	wire _0150_;
	wire _0151_;
	wire _0152_;
	wire _0153_;
	wire _0154_;
	wire _0155_;
	wire _0156_;
	wire _0157_;
	wire _0158_;
	wire _0159_;
	wire _0160_;
	wire _0161_;
	wire _0162_;
	wire _0163_;
	wire _0164_;
	wire _0165_;
	wire _0166_;
	wire _0167_;
	wire _0168_;
	wire _0169_;
	wire _0170_;
	wire _0171_;
	wire _0172_;
	wire _0173_;
	wire _0174_;
	wire _0175_;
	wire _0176_;
	wire _0177_;
	wire _0178_;
	wire _0179_;
	wire _0180_;
	wire _0181_;
	wire _0182_;
	wire _0183_;
	wire _0184_;
	wire _0185_;
	wire _0186_;
	wire _0187_;
	wire _0188_;
	wire _0189_;
	wire _0190_;
	wire _0191_;
	wire _0192_;
	wire _0193_;
	wire _0194_;
	wire _0195_;
	wire _0196_;
	wire _0197_;
	wire _0198_;
	wire _0199_;
	wire _0200_;
	wire _0201_;
	wire _0202_;
	wire _0203_;
	wire _0204_;
	wire _0205_;
	wire _0206_;
	wire _0207_;
	wire _0208_;
	wire _0209_;
	wire _0210_;
	wire _0211_;
	wire _0212_;
	wire _0213_;
	wire _0214_;
	wire _0215_;
	wire _0216_;
	wire _0217_;
	wire _0218_;
	wire _0219_;
	wire _0220_;
	wire _0221_;
	wire _0222_;
	wire _0223_;
	wire _0224_;
	wire _0225_;
	wire _0226_;
	wire _0227_;
	wire _0228_;
	wire _0229_;
	wire _0230_;
	wire _0231_;
	wire _0232_;
	wire _0233_;
	wire _0234_;
	wire _0235_;
	wire _0236_;
	wire _0237_;
	wire _0238_;
	wire _0239_;
	wire _0240_;
	wire _0241_;
	wire _0242_;
	wire _0243_;
	wire _0244_;
	wire _0245_;
	wire _0246_;
	wire _0247_;
	wire _0248_;
	wire _0249_;
	wire _0250_;
	wire _0251_;
	wire _0252_;
	wire _0253_;
	wire _0254_;
	wire _0255_;
	wire _0256_;
	wire _0257_;
	wire _0258_;
	wire _0259_;
	wire _0260_;
	wire _0261_;
	wire _0262_;
	wire _0263_;
	wire _0264_;
	wire _0265_;
	wire _0266_;
	wire _0267_;
	wire _0268_;
	wire _0269_;
	wire _0270_;
	wire _0271_;
	wire _0272_;
	wire _0273_;
	wire _0274_;
	wire _0275_;
	wire _0276_;
	wire _0277_;
	wire _0278_;
	wire _0279_;
	wire _0280_;
	wire _0281_;
	wire _0282_;
	wire _0283_;
	wire _0284_;
	wire _0285_;
	wire _0286_;
	wire _0287_;
	wire _0288_;
	wire _0289_;
	wire _0290_;
	wire _0291_;
	wire _0292_;
	wire _0293_;
	wire _0294_;
	wire _0295_;
	wire _0296_;
	wire _0297_;
	wire _0298_;
	wire _0299_;
	wire _0300_;
	wire _0301_;
	wire _0302_;
	wire _0303_;
	wire _0304_;
	wire _0305_;
	wire _0306_;
	wire _0307_;
	wire _0308_;
	wire _0309_;
	wire _0310_;
	wire _0311_;
	wire _0312_;
	wire _0313_;
	wire _0314_;
	wire _0315_;
	wire _0316_;
	wire _0317_;
	wire _0318_;
	wire _0319_;
	wire _0320_;
	wire _0321_;
	wire _0322_;
	wire _0323_;
	wire _0324_;
	wire _0325_;
	wire _0326_;
	wire _0327_;
	wire _0328_;
	wire _0329_;
	wire _0330_;
	wire _0331_;
	wire _0332_;
	wire _0333_;
	wire _0334_;
	wire _0335_;
	wire _0336_;
	wire _0337_;
	wire _0338_;
	wire _0339_;
	wire _0340_;
	wire _0341_;
	wire _0342_;
	wire _0343_;
	wire _0344_;
	wire _0345_;
	wire _0346_;
	wire _0347_;
	wire _0348_;
	wire _0349_;
	wire _0350_;
	wire _0351_;
	wire _0352_;
	wire _0353_;
	wire _0354_;
	wire _0355_;
	wire _0356_;
	wire _0357_;
	wire _0358_;
	wire _0359_;
	wire _0360_;
	wire _0361_;
	wire _0362_;
	wire _0363_;
	wire _0364_;
	wire _0365_;
	wire _0366_;
	wire _0367_;
	wire _0368_;
	wire _0369_;
	wire _0370_;
	wire _0371_;
	wire _0372_;
	wire _0373_;
	wire _0374_;
	wire _0375_;
	wire _0376_;
	wire _0377_;
	wire _0378_;
	wire _0379_;
	wire _0380_;
	wire _0381_;
	wire _0382_;
	wire _0383_;
	wire _0384_;
	wire _0385_;
	wire _0386_;
	wire _0387_;
	wire _0388_;
	wire _0389_;
	wire _0390_;
	wire _0391_;
	wire _0392_;
	wire _0393_;
	wire _0394_;
	wire _0395_;
	wire _0396_;
	wire _0397_;
	wire _0398_;
	wire _0399_;
	wire _0400_;
	wire _0401_;
	wire _0402_;
	wire _0403_;
	wire _0404_;
	wire _0405_;
	wire _0406_;
	wire _0407_;
	wire _0408_;
	wire _0409_;
	wire _0410_;
	wire _0411_;
	wire _0412_;
	wire _0413_;
	wire _0414_;
	wire _0415_;
	wire _0416_;
	wire _0417_;
	wire _0418_;
	wire _0419_;
	wire _0420_;
	wire _0421_;
	wire _0422_;
	wire _0423_;
	wire _0424_;
	wire _0425_;
	wire _0426_;
	wire _0427_;
	wire _0428_;
	wire _0429_;
	wire _0430_;
	wire _0431_;
	wire _0432_;
	wire _0433_;
	wire _0434_;
	wire _0435_;
	wire _0436_;
	wire _0437_;
	wire _0438_;
	wire _0439_;
	wire _0440_;
	wire _0441_;
	wire _0442_;
	wire _0443_;
	wire _0444_;
	wire _0445_;
	wire _0446_;
	wire _0447_;
	wire _0448_;
	wire _0449_;
	wire _0450_;
	wire _0451_;
	wire _0452_;
	wire _0453_;
	wire _0454_;
	wire _0455_;
	wire _0456_;
	wire _0457_;
	wire _0458_;
	wire _0459_;
	wire _0460_;
	wire _0461_;
	wire _0462_;
	wire _0463_;
	wire _0464_;
	wire _0465_;
	wire _0466_;
	wire _0467_;
	wire _0468_;
	wire _0469_;
	wire _0470_;
	wire _0471_;
	wire _0472_;
	wire _0473_;
	wire _0474_;
	wire _0475_;
	wire _0476_;
	wire _0477_;
	wire _0478_;
	wire _0479_;
	wire _0480_;
	wire _0481_;
	wire _0482_;
	wire _0483_;
	wire _0484_;
	wire _0485_;
	wire _0486_;
	wire _0487_;
	wire _0488_;
	wire _0489_;
	wire _0490_;
	wire _0491_;
	wire _0492_;
	wire _0493_;
	wire _0494_;
	wire _0495_;
	wire _0496_;
	wire _0497_;
	wire _0498_;
	wire _0499_;
	wire _0500_;
	wire _0501_;
	wire _0502_;
	wire _0503_;
	wire _0504_;
	wire _0505_;
	wire _0506_;
	wire _0507_;
	wire _0508_;
	wire _0509_;
	wire _0510_;
	wire _0511_;
	wire _0512_;
	wire _0513_;
	wire _0514_;
	wire _0515_;
	wire _0516_;
	wire _0517_;
	wire _0518_;
	wire _0519_;
	wire _0520_;
	wire _0521_;
	wire _0522_;
	wire _0523_;
	wire _0524_;
	wire _0525_;
	wire _0526_;
	wire _0527_;
	wire _0528_;
	wire _0529_;
	wire _0530_;
	wire _0531_;
	wire _0532_;
	wire _0533_;
	wire _0534_;
	wire _0535_;
	wire _0536_;
	wire _0537_;
	wire _0538_;
	wire _0539_;
	wire _0540_;
	wire _0541_;
	wire _0542_;
	wire _0543_;
	wire _0544_;
	wire _0545_;
	wire _0546_;
	wire _0547_;
	wire _0548_;
	wire _0549_;
	wire _0550_;
	wire _0551_;
	wire _0552_;
	wire _0553_;
	wire _0554_;
	wire _0555_;
	wire _0556_;
	wire _0557_;
	wire _0558_;
	wire _0559_;
	wire _0560_;
	wire _0561_;
	wire _0562_;
	wire _0563_;
	wire _0564_;
	wire _0565_;
	wire _0566_;
	wire _0567_;
	wire _0568_;
	wire _0569_;
	wire _0570_;
	wire _0571_;
	wire _0572_;
	wire _0573_;
	wire _0574_;
	wire _0575_;
	wire _0576_;
	wire _0577_;
	wire _0578_;
	wire _0579_;
	wire _0580_;
	wire _0581_;
	wire _0582_;
	wire _0583_;
	wire _0584_;
	wire _0585_;
	wire _0586_;
	wire _0587_;
	wire _0588_;
	wire _0589_;
	wire _0590_;
	wire _0591_;
	wire _0592_;
	wire _0593_;
	wire _0594_;
	wire _0595_;
	wire _0596_;
	wire _0597_;
	wire _0598_;
	wire _0599_;
	wire _0600_;
	wire _0601_;
	wire _0602_;
	wire _0603_;
	wire _0604_;
	wire _0605_;
	wire _0606_;
	wire _0607_;
	wire _0608_;
	wire _0609_;
	wire _0610_;
	wire _0611_;
	wire _0612_;
	wire _0613_;
	wire _0614_;
	wire _0615_;
	wire _0616_;
	wire _0617_;
	wire _0618_;
	wire _0619_;
	wire _0620_;
	wire _0621_;
	wire _0622_;
	wire _0623_;
	wire _0624_;
	wire _0625_;
	wire _0626_;
	wire _0627_;
	wire _0628_;
	wire _0629_;
	wire _0630_;
	wire _0631_;
	wire _0632_;
	wire _0633_;
	wire _0634_;
	wire _0635_;
	wire _0636_;
	wire _0637_;
	wire _0638_;
	wire _0639_;
	wire _0640_;
	wire _0641_;
	wire _0642_;
	wire _0643_;
	wire _0644_;
	wire _0645_;
	wire _0646_;
	wire _0647_;
	wire _0648_;
	wire _0649_;
	wire _0650_;
	wire _0651_;
	wire _0652_;
	wire _0653_;
	wire _0654_;
	wire _0655_;
	wire _0656_;
	wire _0657_;
	wire _0658_;
	wire _0659_;
	wire _0660_;
	wire _0661_;
	wire _0662_;
	wire _0663_;
	wire _0664_;
	wire _0665_;
	wire _0666_;
	wire _0667_;
	wire _0668_;
	wire _0669_;
	wire _0670_;
	wire _0671_;
	wire _0672_;
	wire _0673_;
	wire _0674_;
	wire _0675_;
	wire _0676_;
	wire _0677_;
	wire _0678_;
	wire _0679_;
	wire _0680_;
	wire _0681_;
	wire _0682_;
	wire _0683_;
	wire _0684_;
	wire _0685_;
	wire _0686_;
	wire _0687_;
	wire _0688_;
	wire _0689_;
	wire _0690_;
	wire _0691_;
	wire _0692_;
	wire _0693_;
	wire _0694_;
	wire _0695_;
	wire _0696_;
	wire _0697_;
	wire _0698_;
	wire _0699_;
	wire _0700_;
	wire _0701_;
	wire _0702_;
	wire _0703_;
	wire _0704_;
	wire _0705_;
	wire _0706_;
	wire _0707_;
	wire _0708_;
	wire _0709_;
	wire _0710_;
	wire _0711_;
	wire _0712_;
	wire _0713_;
	wire _0714_;
	wire _0715_;
	wire _0716_;
	wire _0717_;
	wire _0718_;
	wire _0719_;
	wire _0720_;
	wire _0721_;
	wire _0722_;
	wire _0723_;
	wire _0724_;
	wire _0725_;
	wire _0726_;
	wire _0727_;
	wire _0728_;
	wire _0729_;
	wire _0730_;
	wire _0731_;
	wire _0732_;
	wire _0733_;
	wire _0734_;
	wire _0735_;
	wire _0736_;
	wire _0737_;
	wire _0738_;
	wire _0739_;
	wire _0740_;
	wire _0741_;
	wire _0742_;
	wire _0743_;
	wire _0744_;
	wire _0745_;
	wire _0746_;
	wire _0747_;
	wire _0748_;
	wire _0749_;
	wire _0750_;
	wire _0751_;
	wire _0752_;
	wire _0753_;
	wire _0754_;
	wire _0755_;
	wire _0756_;
	wire _0757_;
	wire _0758_;
	wire _0759_;
	wire _0760_;
	wire _0761_;
	wire _0762_;
	wire _0763_;
	wire _0764_;
	wire _0765_;
	wire _0766_;
	wire _0767_;
	wire _0768_;
	wire _0769_;
	wire _0770_;
	wire _0771_;
	wire _0772_;
	wire _0773_;
	wire _0774_;
	wire _0775_;
	wire _0776_;
	wire _0777_;
	wire _0778_;
	wire _0779_;
	wire _0780_;
	wire _0781_;
	wire _0782_;
	wire _0783_;
	wire _0784_;
	wire _0785_;
	wire _0786_;
	wire _0787_;
	wire _0788_;
	wire _0789_;
	wire _0790_;
	wire _0791_;
	wire _0792_;
	wire _0793_;
	wire _0794_;
	wire _0795_;
	wire _0796_;
	wire _0797_;
	wire _0798_;
	wire _0799_;
	wire _0800_;
	wire _0801_;
	wire _0802_;
	wire _0803_;
	wire _0804_;
	wire _0805_;
	wire _0806_;
	wire _0807_;
	wire _0808_;
	wire _0809_;
	wire _0810_;
	wire _0811_;
	wire _0812_;
	wire _0813_;
	wire _0814_;
	wire _0815_;
	wire _0816_;
	wire _0817_;
	wire _0818_;
	wire _0819_;
	wire _0820_;
	wire _0821_;
	wire _0822_;
	wire _0823_;
	wire _0824_;
	wire _0825_;
	wire _0826_;
	wire _0827_;
	wire _0828_;
	wire _0829_;
	wire _0830_;
	wire _0831_;
	wire _0832_;
	wire _0833_;
	wire _0834_;
	wire _0835_;
	wire _0836_;
	wire _0837_;
	wire _0838_;
	wire _0839_;
	wire _0840_;
	wire _0841_;
	wire _0842_;
	wire _0843_;
	wire _0844_;
	wire _0845_;
	wire _0846_;
	wire _0847_;
	wire _0848_;
	wire _0849_;
	wire _0850_;
	wire _0851_;
	wire _0852_;
	wire _0853_;
	wire _0854_;
	wire _0855_;
	wire _0856_;
	wire _0857_;
	wire _0858_;
	wire _0859_;
	wire _0860_;
	wire _0861_;
	wire _0862_;
	wire _0863_;
	wire _0864_;
	wire _0865_;
	wire _0866_;
	wire _0867_;
	wire _0868_;
	wire _0869_;
	wire _0870_;
	wire _0871_;
	wire _0872_;
	wire _0873_;
	wire _0874_;
	wire _0875_;
	wire _0876_;
	wire _0877_;
	wire _0878_;
	wire _0879_;
	wire _0880_;
	wire _0881_;
	wire _0882_;
	wire _0883_;
	wire _0884_;
	wire _0885_;
	wire _0886_;
	wire _0887_;
	wire _0888_;
	wire _0889_;
	wire _0890_;
	wire _0891_;
	wire _0892_;
	wire _0893_;
	wire _0894_;
	wire _0895_;
	wire _0896_;
	wire _0897_;
	wire _0898_;
	wire _0899_;
	wire _0900_;
	wire _0901_;
	wire _0902_;
	wire _0903_;
	wire _0904_;
	wire _0905_;
	wire _0906_;
	wire _0907_;
	wire _0908_;
	wire _0909_;
	wire _0910_;
	wire _0911_;
	wire _0912_;
	wire _0913_;
	wire _0914_;
	wire _0915_;
	wire _0916_;
	wire _0917_;
	wire _0918_;
	wire _0919_;
	wire _0920_;
	wire _0921_;
	wire _0922_;
	wire _0923_;
	wire _0924_;
	wire _0925_;
	wire _0926_;
	wire _0927_;
	wire _0928_;
	wire _0929_;
	wire _0930_;
	wire _0931_;
	wire _0932_;
	wire _0933_;
	wire _0934_;
	wire _0935_;
	wire _0936_;
	wire _0937_;
	wire _0938_;
	wire _0939_;
	wire _0940_;
	wire _0941_;
	wire _0942_;
	wire _0943_;
	wire _0944_;
	wire _0945_;
	wire _0946_;
	wire _0947_;
	wire _0948_;
	wire _0949_;
	wire _0950_;
	wire _0951_;
	wire _0952_;
	wire _0953_;
	wire _0954_;
	wire _0955_;
	wire _0956_;
	wire _0957_;
	wire _0958_;
	wire _0959_;
	wire _0960_;
	wire _0961_;
	wire _0962_;
	wire _0963_;
	wire _0964_;
	wire _0965_;
	wire _0966_;
	wire _0967_;
	wire _0968_;
	wire _0969_;
	wire _0970_;
	wire _0971_;
	wire _0972_;
	wire _0973_;
	wire _0974_;
	wire _0975_;
	wire _0976_;
	wire _0977_;
	wire _0978_;
	wire _0979_;
	wire _0980_;
	wire _0981_;
	wire _0982_;
	wire _0983_;
	wire _0984_;
	wire _0985_;
	wire _0986_;
	wire _0987_;
	wire _0988_;
	wire _0989_;
	wire _0990_;
	wire _0991_;
	wire _0992_;
	wire _0993_;
	wire _0994_;
	wire _0995_;
	wire _0996_;
	wire _0997_;
	wire _0998_;
	wire _0999_;
	wire _1000_;
	wire _1001_;
	wire _1002_;
	wire _1003_;
	wire _1004_;
	wire _1005_;
	wire _1006_;
	wire _1007_;
	wire _1008_;
	wire _1009_;
	wire _1010_;
	wire _1011_;
	wire _1012_;
	wire _1013_;
	wire _1014_;
	wire _1015_;
	wire _1016_;
	wire _1017_;
	wire _1018_;
	wire _1019_;
	wire _1020_;
	wire _1021_;
	wire _1022_;
	wire _1023_;
	wire _1024_;
	wire _1025_;
	wire _1026_;
	wire _1027_;
	wire _1028_;
	wire _1029_;
	wire _1030_;
	wire _1031_;
	wire _1032_;
	wire _1033_;
	wire _1034_;
	wire _1035_;
	wire _1036_;
	wire _1037_;
	wire _1038_;
	wire _1039_;
	wire _1040_;
	wire _1041_;
	wire _1042_;
	wire _1043_;
	wire _1044_;
	wire _1045_;
	wire _1046_;
	wire _1047_;
	wire _1048_;
	wire _1049_;
	wire _1050_;
	wire _1051_;
	wire _1052_;
	wire _1053_;
	wire _1054_;
	wire _1055_;
	wire _1056_;
	wire _1057_;
	wire _1058_;
	wire _1059_;
	wire _1060_;
	wire _1061_;
	wire _1062_;
	wire _1063_;
	wire _1064_;
	wire _1065_;
	wire _1066_;
	wire _1067_;
	wire _1068_;
	wire _1069_;
	wire _1070_;
	wire _1071_;
	wire _1072_;
	wire _1073_;
	wire _1074_;
	wire _1075_;
	wire _1076_;
	wire _1077_;
	wire _1078_;
	wire _1079_;
	wire _1080_;
	wire _1081_;
	wire _1082_;
	wire _1083_;
	wire _1084_;
	wire _1085_;
	wire _1086_;
	wire _1087_;
	wire _1088_;
	wire _1089_;
	wire _1090_;
	wire _1091_;
	wire _1092_;
	wire _1093_;
	wire _1094_;
	wire _1095_;
	wire _1096_;
	wire _1097_;
	wire _1098_;
	wire _1099_;
	wire _1100_;
	wire _1101_;
	wire _1102_;
	wire _1103_;
	wire _1104_;
	wire _1105_;
	wire _1106_;
	wire _1107_;
	wire _1108_;
	wire _1109_;
	wire _1110_;
	wire _1111_;
	wire _1112_;
	wire _1113_;
	wire _1114_;
	wire _1115_;
	wire _1116_;
	wire _1117_;
	wire _1118_;
	wire _1119_;
	wire _1120_;
	wire _1121_;
	wire _1122_;
	wire _1123_;
	wire _1124_;
	wire _1125_;
	wire _1126_;
	wire _1127_;
	wire _1128_;
	wire _1129_;
	wire _1130_;
	wire _1131_;
	wire _1132_;
	wire _1133_;
	wire _1134_;
	wire _1135_;
	wire _1136_;
	wire _1137_;
	wire _1138_;
	wire _1139_;
	wire _1140_;
	wire _1141_;
	wire _1142_;
	wire _1143_;
	wire _1144_;
	wire _1145_;
	wire _1146_;
	wire _1147_;
	wire _1148_;
	wire _1149_;
	wire _1150_;
	wire _1151_;
	wire _1152_;
	wire _1153_;
	wire _1154_;
	wire _1155_;
	wire _1156_;
	wire _1157_;
	wire _1158_;
	wire _1159_;
	wire _1160_;
	wire _1161_;
	wire _1162_;
	wire _1163_;
	wire _1164_;
	wire _1165_;
	wire _1166_;
	wire _1167_;
	wire _1168_;
	wire _1169_;
	wire _1170_;
	wire _1171_;
	wire _1172_;
	wire _1173_;
	wire _1174_;
	wire _1175_;
	wire _1176_;
	wire _1177_;
	wire _1178_;
	wire _1179_;
	wire _1180_;
	wire _1181_;
	wire _1182_;
	wire _1183_;
	wire _1184_;
	wire _1185_;
	wire _1186_;
	wire _1187_;
	wire _1188_;
	wire _1189_;
	wire _1190_;
	wire _1191_;
	wire _1192_;
	wire _1193_;
	wire _1194_;
	wire _1195_;
	wire _1196_;
	wire _1197_;
	wire _1198_;
	wire _1199_;
	wire _1200_;
	wire _1201_;
	wire _1202_;
	wire _1203_;
	wire _1204_;
	wire _1205_;
	wire _1206_;
	wire _1207_;
	wire _1208_;
	wire _1209_;
	wire _1210_;
	wire _1211_;
	wire _1212_;
	wire _1213_;
	wire _1214_;
	wire _1215_;
	wire _1216_;
	wire _1217_;
	wire _1218_;
	wire _1219_;
	wire _1220_;
	wire _1221_;
	wire _1222_;
	wire _1223_;
	wire _1224_;
	wire _1225_;
	wire _1226_;
	wire _1227_;
	wire _1228_;
	wire _1229_;
	wire _1230_;
	wire _1231_;
	wire _1232_;
	wire _1233_;
	wire _1234_;
	wire _1235_;
	wire _1236_;
	wire _1237_;
	wire _1238_;
	wire _1239_;
	wire _1240_;
	wire _1241_;
	wire _1242_;
	wire _1243_;
	wire _1244_;
	wire _1245_;
	wire _1246_;
	wire _1247_;
	wire _1248_;
	wire _1249_;
	wire _1250_;
	wire _1251_;
	wire _1252_;
	wire _1253_;
	wire _1254_;
	wire _1255_;
	wire _1256_;
	wire _1257_;
	wire _1258_;
	wire _1259_;
	wire _1260_;
	wire _1261_;
	wire _1262_;
	wire _1263_;
	wire _1264_;
	wire _1265_;
	wire _1266_;
	wire _1267_;
	wire _1268_;
	wire _1269_;
	wire _1270_;
	wire _1271_;
	wire _1272_;
	wire _1273_;
	wire _1274_;
	wire _1275_;
	wire _1276_;
	wire _1277_;
	wire _1278_;
	wire _1279_;
	wire _1280_;
	wire _1281_;
	wire _1282_;
	wire _1283_;
	wire _1284_;
	wire _1285_;
	wire _1286_;
	wire _1287_;
	wire _1288_;
	wire _1289_;
	wire _1290_;
	wire _1291_;
	wire _1292_;
	wire _1293_;
	wire _1294_;
	wire _1295_;
	wire _1296_;
	wire _1297_;
	wire _1298_;
	wire _1299_;
	wire _1300_;
	wire _1301_;
	wire _1302_;
	wire _1303_;
	wire _1304_;
	wire _1305_;
	wire _1306_;
	wire _1307_;
	wire _1308_;
	wire _1309_;
	wire _1310_;
	wire _1311_;
	wire _1312_;
	wire _1313_;
	wire _1314_;
	wire _1315_;
	wire _1316_;
	wire _1317_;
	wire _1318_;
	wire _1319_;
	wire _1320_;
	wire _1321_;
	wire _1322_;
	wire _1323_;
	wire _1324_;
	wire _1325_;
	wire _1326_;
	wire _1327_;
	wire _1328_;
	wire _1329_;
	wire _1330_;
	wire _1331_;
	wire _1332_;
	wire _1333_;
	wire _1334_;
	wire _1335_;
	wire _1336_;
	wire _1337_;
	wire _1338_;
	wire _1339_;
	wire _1340_;
	wire _1341_;
	wire _1342_;
	wire _1343_;
	wire _1344_;
	wire _1345_;
	wire _1346_;
	wire _1347_;
	wire _1348_;
	wire _1349_;
	wire _1350_;
	wire _1351_;
	wire _1352_;
	wire _1353_;
	wire _1354_;
	wire _1355_;
	wire _1356_;
	wire _1357_;
	wire _1358_;
	wire _1359_;
	wire _1360_;
	wire _1361_;
	wire _1362_;
	wire _1363_;
	wire _1364_;
	wire _1365_;
	wire _1366_;
	wire _1367_;
	wire _1368_;
	wire _1369_;
	wire _1370_;
	wire _1371_;
	wire _1372_;
	wire _1373_;
	wire _1374_;
	wire _1375_;
	wire _1376_;
	wire _1377_;
	wire _1378_;
	wire _1379_;
	wire _1380_;
	wire _1381_;
	wire _1382_;
	wire _1383_;
	wire _1384_;
	wire _1385_;
	wire _1386_;
	wire _1387_;
	wire _1388_;
	wire _1389_;
	wire _1390_;
	wire _1391_;
	wire _1392_;
	wire _1393_;
	wire _1394_;
	wire _1395_;
	wire _1396_;
	wire _1397_;
	wire _1398_;
	wire _1399_;
	wire _1400_;
	wire _1401_;
	wire _1402_;
	wire _1403_;
	wire _1404_;
	wire _1405_;
	wire _1406_;
	wire _1407_;
	wire _1408_;
	wire _1409_;
	wire _1410_;
	wire _1411_;
	wire _1412_;
	wire _1413_;
	wire _1414_;
	wire _1415_;
	wire _1416_;
	wire _1417_;
	wire _1418_;
	wire _1419_;
	wire _1420_;
	wire _1421_;
	wire _1422_;
	wire _1423_;
	wire _1424_;
	wire _1425_;
	wire _1426_;
	wire _1427_;
	wire _1428_;
	wire _1429_;
	wire _1430_;
	wire _1431_;
	wire _1432_;
	wire _1433_;
	wire _1434_;
	wire _1435_;
	wire _1436_;
	wire _1437_;
	wire _1438_;
	wire _1439_;
	wire _1440_;
	wire _1441_;
	wire _1442_;
	wire _1443_;
	wire _1444_;
	wire _1445_;
	wire _1446_;
	wire _1447_;
	wire _1448_;
	wire _1449_;
	wire _1450_;
	wire _1451_;
	wire _1452_;
	wire _1453_;
	wire _1454_;
	wire _1455_;
	wire _1456_;
	wire _1457_;
	wire _1458_;
	wire _1459_;
	wire _1460_;
	wire _1461_;
	wire _1462_;
	wire _1463_;
	wire _1464_;
	wire _1465_;
	wire _1466_;
	wire _1467_;
	wire _1468_;
	wire _1469_;
	wire _1470_;
	wire _1471_;
	wire _1472_;
	wire _1473_;
	wire _1474_;
	wire _1475_;
	wire _1476_;
	wire _1477_;
	wire _1478_;
	wire _1479_;
	wire _1480_;
	wire _1481_;
	wire _1482_;
	wire _1483_;
	wire _1484_;
	wire _1485_;
	wire _1486_;
	wire _1487_;
	wire _1488_;
	wire _1489_;
	wire _1490_;
	wire _1491_;
	wire _1492_;
	wire _1493_;
	wire _1494_;
	wire _1495_;
	wire _1496_;
	wire _1497_;
	wire _1498_;
	wire _1499_;
	wire _1500_;
	wire _1501_;
	wire _1502_;
	wire _1503_;
	wire _1504_;
	wire _1505_;
	wire _1506_;
	wire _1507_;
	wire _1508_;
	wire _1509_;
	wire _1510_;
	wire _1511_;
	wire _1512_;
	wire _1513_;
	wire _1514_;
	wire _1515_;
	wire _1516_;
	wire _1517_;
	wire _1518_;
	wire _1519_;
	wire _1520_;
	wire _1521_;
	wire _1522_;
	wire _1523_;
	wire _1524_;
	wire _1525_;
	wire _1526_;
	wire _1527_;
	wire _1528_;
	wire _1529_;
	wire _1530_;
	wire _1531_;
	wire _1532_;
	wire _1533_;
	wire _1534_;
	wire _1535_;
	wire _1536_;
	wire _1537_;
	wire _1538_;
	wire _1539_;
	wire _1540_;
	wire _1541_;
	wire _1542_;
	wire _1543_;
	wire _1544_;
	wire _1545_;
	wire _1546_;
	wire _1547_;
	wire _1548_;
	wire _1549_;
	wire _1550_;
	wire _1551_;
	wire _1552_;
	wire _1553_;
	wire _1554_;
	wire _1555_;
	wire _1556_;
	wire _1557_;
	wire _1558_;
	wire _1559_;
	wire _1560_;
	wire _1561_;
	wire _1562_;
	wire _1563_;
	wire _1564_;
	wire _1565_;
	wire _1566_;
	wire _1567_;
	wire _1568_;
	wire _1569_;
	wire _1570_;
	wire _1571_;
	wire _1572_;
	wire _1573_;
	wire _1574_;
	wire _1575_;
	wire _1576_;
	wire _1577_;
	wire _1578_;
	wire _1579_;
	wire _1580_;
	wire _1581_;
	wire _1582_;
	wire _1583_;
	wire _1584_;
	wire _1585_;
	wire _1586_;
	wire _1587_;
	wire _1588_;
	wire _1589_;
	wire _1590_;
	wire _1591_;
	wire _1592_;
	wire _1593_;
	wire _1594_;
	wire _1595_;
	wire _1596_;
	wire _1597_;
	wire _1598_;
	wire _1599_;
	wire _1600_;
	wire _1601_;
	wire _1602_;
	wire _1603_;
	wire _1604_;
	wire _1605_;
	wire _1606_;
	wire _1607_;
	wire _1608_;
	wire _1609_;
	wire _1610_;
	wire _1611_;
	wire _1612_;
	wire _1613_;
	wire _1614_;
	wire _1615_;
	wire _1616_;
	wire _1617_;
	wire _1618_;
	wire _1619_;
	wire _1620_;
	wire _1621_;
	wire _1622_;
	wire _1623_;
	wire _1624_;
	wire _1625_;
	wire _1626_;
	wire _1627_;
	wire _1628_;
	wire _1629_;
	wire _1630_;
	wire _1631_;
	wire _1632_;
	wire _1633_;
	wire _1634_;
	wire _1635_;
	wire _1636_;
	wire _1637_;
	wire _1638_;
	wire _1639_;
	wire _1640_;
	wire _1641_;
	wire _1642_;
	wire _1643_;
	wire _1644_;
	wire _1645_;
	wire _1646_;
	wire _1647_;
	wire _1648_;
	wire _1649_;
	wire _1650_;
	wire _1651_;
	wire _1652_;
	wire _1653_;
	wire _1654_;
	wire _1655_;
	wire _1656_;
	wire _1657_;
	wire _1658_;
	wire _1659_;
	wire _1660_;
	wire _1661_;
	wire _1662_;
	wire _1663_;
	wire _1664_;
	wire _1665_;
	wire _1666_;
	wire _1667_;
	wire _1668_;
	wire _1669_;
	wire _1670_;
	wire _1671_;
	wire _1672_;
	wire _1673_;
	wire _1674_;
	wire _1675_;
	wire _1676_;
	wire _1677_;
	wire _1678_;
	wire _1679_;
	wire _1680_;
	wire _1681_;
	wire _1682_;
	wire _1683_;
	wire _1684_;
	wire _1685_;
	wire _1686_;
	wire _1687_;
	wire _1688_;
	wire _1689_;
	wire _1690_;
	wire _1691_;
	wire _1692_;
	wire _1693_;
	wire _1694_;
	wire _1695_;
	wire _1696_;
	wire _1697_;
	wire _1698_;
	wire _1699_;
	wire _1700_;
	wire _1701_;
	wire _1702_;
	wire _1703_;
	wire _1704_;
	wire _1705_;
	wire _1706_;
	wire _1707_;
	wire _1708_;
	wire _1709_;
	wire _1710_;
	wire _1711_;
	wire _1712_;
	wire _1713_;
	wire _1714_;
	wire _1715_;
	wire _1716_;
	wire _1717_;
	wire _1718_;
	wire _1719_;
	wire _1720_;
	wire _1721_;
	wire _1722_;
	wire _1723_;
	wire _1724_;
	wire _1725_;
	wire _1726_;
	wire _1727_;
	wire _1728_;
	wire _1729_;
	wire _1730_;
	wire _1731_;
	wire _1732_;
	wire _1733_;
	wire _1734_;
	wire _1735_;
	wire _1736_;
	wire _1737_;
	wire _1738_;
	wire _1739_;
	wire _1740_;
	input wire [13:0] io_in;
	output wire [13:0] io_out;
	wire [7:0] \mchip.byte_in ;
	wire [7:0] \mchip.byte_out ;
	wire \mchip.clock ;
	reg [127:0] \mchip.internal ;
	wire [11:0] \mchip.io_in ;
	wire [11:0] \mchip.io_out ;
	wire \mchip.is_active ;
	reg [127:0] \mchip.key ;
	wire \mchip.key_in ;
	reg \mchip.key_in_last ;
	reg [127:0] \mchip.plaintext ;
	wire \mchip.plaintext_in ;
	reg \mchip.plaintext_in_last ;
	wire \mchip.reset ;
	wire [7:0] \mchip.sbox.s ;
	wire [7:0] \mchip.sbox.sbox_in ;
	wire [7:0] \mchip.sbox.sbox_out ;
	wire [67:0] \mchip.sbox.t ;
	wire [7:0] \mchip.sbox.u ;
	wire [21:0] \mchip.sbox.y ;
	wire [17:0] \mchip.sbox.z ;
	wire [7:0] \mchip.sbox_out ;
	wire \mchip.start ;
	reg [6:0] \mchip.state ;
	assign _1304_ = ~(\mchip.state [5] | \mchip.state [4]);
	assign _1305_ = _1304_ & ~\mchip.state [6];
	assign _1306_ = ~(\mchip.state [2] | \mchip.state [3]);
	assign _1307_ = ~(\mchip.state [0] | \mchip.state [1]);
	assign _1308_ = ~(_1307_ & _1306_);
	assign \mchip.is_active  = _1308_ | ~_1305_;
	assign _0136_ = io_in[10] & ~\mchip.is_active ;
	assign _1309_ = ~\mchip.state [0];
	assign _1310_ = \mchip.state [6] | \mchip.state [5];
	assign _1311_ = _1310_ | _1309_;
	assign _1312_ = \mchip.state [4] | \mchip.state [3];
	assign _1313_ = \mchip.state [2] | \mchip.state [1];
	assign _1314_ = _1313_ | _1312_;
	assign _1315_ = _1314_ | _1311_;
	assign _1316_ = _1315_ | io_in[10];
	assign _0002_ = _0136_ | ~_1316_;
	assign _1317_ = ~(_1314_ | _1310_);
	assign _1318_ = ~_1317_;
	assign _1319_ = io_in[13] | ~_1316_;
	assign _0001_ = _1319_ | _1318_;
	assign _0000_ = io_in[13] | ~_1317_;
	assign _1320_ = ~_1304_;
	assign _1321_ = ~_1306_;
	assign _1322_ = \mchip.state [2] & ~\mchip.state [3];
	assign _1323_ = _1322_ & _1307_;
	assign _1324_ = _1321_ & ~_1323_;
	assign _1325_ = _1324_ | _1320_;
	assign _1326_ = _1325_ | \mchip.state [6];
	assign _1327_ = _1323_ & _1305_;
	assign _1328_ = _1327_ | _1326_;
	assign _1329_ = ~\mchip.state [6];
	assign _1330_ = \mchip.state [4] & ~\mchip.state [5];
	assign _1331_ = ~(_1330_ & _1329_);
	assign _1332_ = _1323_ & ~_1331_;
	assign _1333_ = _1330_ & ~_1324_;
	assign _1334_ = _1320_ & ~_1333_;
	assign _1335_ = _1334_ | \mchip.state [6];
	assign _1336_ = _1335_ | _1332_;
	assign _0137_ = _1328_ & ~_1336_;
	assign _0135_ = io_in[9] & ~\mchip.plaintext_in_last ;
	assign _0134_ = io_in[8] & ~\mchip.key_in_last ;
	assign _1337_ = \mchip.key [14] ^ \mchip.plaintext [14];
	assign _1338_ = \mchip.state [5] & ~\mchip.state [4];
	assign _1339_ = _1338_ & ~\mchip.state [6];
	assign _1340_ = \mchip.state [3] & ~\mchip.state [2];
	assign _1341_ = _1340_ & _1307_;
	assign _1342_ = ~(_1341_ & _1339_);
	assign _1343_ = (_1342_ ? \mchip.internal [14] : _1337_);
	assign _1344_ = \mchip.state [2] & \mchip.state [1];
	assign _1345_ = _1313_ & ~_1344_;
	assign _1346_ = ~\mchip.state [3];
	assign _1347_ = _1344_ ^ _1346_;
	assign _1348_ = ~(_1347_ | _1345_);
	assign _1349_ = \mchip.state [1] & ~\mchip.state [0];
	assign _1350_ = ~_1349_;
	assign _1351_ = _1348_ & ~_1350_;
	assign _1352_ = ~\mchip.state [4];
	assign _1353_ = _1346_ & ~_1344_;
	assign _1354_ = _1353_ ^ _1352_;
	assign _1355_ = ~\mchip.state [5];
	assign _1356_ = \mchip.state [4] & \mchip.state [3];
	assign _1357_ = \mchip.state [3] | ~\mchip.state [4];
	assign _1358_ = _1344_ & ~_1357_;
	assign _1359_ = _1358_ | _1356_;
	assign _1360_ = _1359_ ^ _1355_;
	assign _1361_ = _1360_ | _1354_;
	assign _1362_ = _1351_ & ~_1361_;
	assign _1363_ = _1355_ & ~_1359_;
	assign _1364_ = _1363_ ^ \mchip.state [6];
	assign _1365_ = _1362_ & ~_1364_;
	assign _1366_ = ~(_1359_ | _1310_);
	assign _1367_ = ~(_1366_ ^ _1365_);
	assign _1368_ = (\mchip.state [0] ? \mchip.internal [127] : \mchip.internal [126]);
	assign _1369_ = (\mchip.state [0] ? \mchip.internal [125] : \mchip.internal [124]);
	assign _1370_ = (\mchip.state [1] ? _1369_ : _1368_);
	assign _1371_ = (\mchip.state [0] ? \mchip.internal [123] : \mchip.internal [122]);
	assign _1372_ = (\mchip.state [0] ? \mchip.internal [121] : \mchip.internal [120]);
	assign _1373_ = (\mchip.state [1] ? _1372_ : _1371_);
	assign _1374_ = (_1345_ ? _1370_ : _1373_);
	assign _1375_ = (\mchip.state [0] ? \mchip.internal [119] : \mchip.internal [118]);
	assign _1376_ = (\mchip.state [0] ? \mchip.internal [117] : \mchip.internal [116]);
	assign _1377_ = (\mchip.state [1] ? _1376_ : _1375_);
	assign _1378_ = (\mchip.state [0] ? \mchip.internal [115] : \mchip.internal [114]);
	assign _1379_ = (\mchip.state [0] ? \mchip.internal [113] : \mchip.internal [112]);
	assign _1380_ = (\mchip.state [1] ? _1379_ : _1378_);
	assign _1381_ = (_1345_ ? _1377_ : _1380_);
	assign _1382_ = (_1347_ ? _1374_ : _1381_);
	assign _1383_ = (\mchip.state [0] ? \mchip.internal [111] : \mchip.internal [110]);
	assign _1384_ = (\mchip.state [0] ? \mchip.internal [109] : \mchip.internal [108]);
	assign _1385_ = (\mchip.state [1] ? _1384_ : _1383_);
	assign _1386_ = (\mchip.state [0] ? \mchip.internal [107] : \mchip.internal [106]);
	assign _1387_ = (\mchip.state [0] ? \mchip.internal [105] : \mchip.internal [104]);
	assign _1388_ = (\mchip.state [1] ? _1387_ : _1386_);
	assign _1389_ = (_1345_ ? _1385_ : _1388_);
	assign _1390_ = (\mchip.state [0] ? \mchip.internal [103] : \mchip.internal [102]);
	assign _1391_ = (\mchip.state [0] ? \mchip.internal [101] : \mchip.internal [100]);
	assign _1392_ = (\mchip.state [1] ? _1391_ : _1390_);
	assign _1393_ = (\mchip.state [0] ? \mchip.internal [99] : \mchip.internal [98]);
	assign _1394_ = (\mchip.state [0] ? \mchip.internal [97] : \mchip.internal [96]);
	assign _1395_ = (\mchip.state [1] ? _1394_ : _1393_);
	assign _1396_ = (_1345_ ? _1392_ : _1395_);
	assign _1397_ = (_1347_ ? _1389_ : _1396_);
	assign _1398_ = (_1354_ ? _1382_ : _1397_);
	assign _1399_ = (\mchip.state [0] ? \mchip.internal [95] : \mchip.internal [94]);
	assign _1400_ = (\mchip.state [0] ? \mchip.internal [93] : \mchip.internal [92]);
	assign _1401_ = (\mchip.state [1] ? _1400_ : _1399_);
	assign _1402_ = (\mchip.state [0] ? \mchip.internal [91] : \mchip.internal [90]);
	assign _1403_ = (\mchip.state [0] ? \mchip.internal [89] : \mchip.internal [88]);
	assign _1404_ = (\mchip.state [1] ? _1403_ : _1402_);
	assign _1405_ = (_1345_ ? _1401_ : _1404_);
	assign _1406_ = (\mchip.state [0] ? \mchip.internal [87] : \mchip.internal [86]);
	assign _1407_ = (\mchip.state [0] ? \mchip.internal [85] : \mchip.internal [84]);
	assign _1408_ = (\mchip.state [1] ? _1407_ : _1406_);
	assign _1409_ = (\mchip.state [0] ? \mchip.internal [83] : \mchip.internal [82]);
	assign _1410_ = (\mchip.state [0] ? \mchip.internal [81] : \mchip.internal [80]);
	assign _1411_ = (\mchip.state [1] ? _1410_ : _1409_);
	assign _1412_ = (_1345_ ? _1408_ : _1411_);
	assign _1413_ = (_1347_ ? _1405_ : _1412_);
	assign _1414_ = (\mchip.state [0] ? \mchip.internal [79] : \mchip.internal [78]);
	assign _1415_ = (\mchip.state [0] ? \mchip.internal [77] : \mchip.internal [76]);
	assign _1416_ = (\mchip.state [1] ? _1415_ : _1414_);
	assign _1417_ = (\mchip.state [0] ? \mchip.internal [75] : \mchip.internal [74]);
	assign _1418_ = (\mchip.state [0] ? \mchip.internal [73] : \mchip.internal [72]);
	assign _1419_ = (\mchip.state [1] ? _1418_ : _1417_);
	assign _1420_ = (_1345_ ? _1416_ : _1419_);
	assign _1421_ = (\mchip.state [0] ? \mchip.internal [71] : \mchip.internal [70]);
	assign _1422_ = (\mchip.state [0] ? \mchip.internal [69] : \mchip.internal [68]);
	assign _1423_ = (\mchip.state [1] ? _1422_ : _1421_);
	assign _1424_ = (\mchip.state [0] ? \mchip.internal [67] : \mchip.internal [66]);
	assign _1425_ = (\mchip.state [0] ? \mchip.internal [65] : \mchip.internal [64]);
	assign _1426_ = (\mchip.state [1] ? _1425_ : _1424_);
	assign _1427_ = (_1345_ ? _1423_ : _1426_);
	assign _1428_ = (_1347_ ? _1420_ : _1427_);
	assign _1429_ = (_1354_ ? _1413_ : _1428_);
	assign _1430_ = (_1360_ ? _1398_ : _1429_);
	assign _1431_ = (\mchip.state [0] ? \mchip.internal [63] : \mchip.internal [62]);
	assign _1432_ = (\mchip.state [0] ? \mchip.internal [61] : \mchip.internal [60]);
	assign _1433_ = (\mchip.state [1] ? _1432_ : _1431_);
	assign _1434_ = (\mchip.state [0] ? \mchip.internal [59] : \mchip.internal [58]);
	assign _1435_ = (\mchip.state [0] ? \mchip.internal [57] : \mchip.internal [56]);
	assign _1436_ = (\mchip.state [1] ? _1435_ : _1434_);
	assign _1437_ = (_1345_ ? _1433_ : _1436_);
	assign _1438_ = (\mchip.state [0] ? \mchip.internal [55] : \mchip.internal [54]);
	assign _1439_ = (\mchip.state [0] ? \mchip.internal [53] : \mchip.internal [52]);
	assign _1440_ = (\mchip.state [1] ? _1439_ : _1438_);
	assign _1441_ = (\mchip.state [0] ? \mchip.internal [51] : \mchip.internal [50]);
	assign _1442_ = (\mchip.state [0] ? \mchip.internal [49] : \mchip.internal [48]);
	assign _1443_ = (\mchip.state [1] ? _1442_ : _1441_);
	assign _1444_ = (_1345_ ? _1440_ : _1443_);
	assign _1445_ = (_1347_ ? _1437_ : _1444_);
	assign _1446_ = (\mchip.state [0] ? \mchip.internal [47] : \mchip.internal [46]);
	assign _1447_ = (\mchip.state [0] ? \mchip.internal [45] : \mchip.internal [44]);
	assign _1448_ = (\mchip.state [1] ? _1447_ : _1446_);
	assign _1449_ = (\mchip.state [0] ? \mchip.internal [43] : \mchip.internal [42]);
	assign _1450_ = (\mchip.state [0] ? \mchip.internal [41] : \mchip.internal [40]);
	assign _1451_ = (\mchip.state [1] ? _1450_ : _1449_);
	assign _1452_ = (_1345_ ? _1448_ : _1451_);
	assign _1453_ = (\mchip.state [0] ? \mchip.internal [39] : \mchip.internal [38]);
	assign _1454_ = (\mchip.state [0] ? \mchip.internal [37] : \mchip.internal [36]);
	assign _1455_ = (\mchip.state [1] ? _1454_ : _1453_);
	assign _1456_ = (\mchip.state [0] ? \mchip.internal [35] : \mchip.internal [34]);
	assign _1457_ = (\mchip.state [0] ? \mchip.internal [33] : \mchip.internal [32]);
	assign _1458_ = (\mchip.state [1] ? _1457_ : _1456_);
	assign _1459_ = (_1345_ ? _1455_ : _1458_);
	assign _1460_ = (_1347_ ? _1452_ : _1459_);
	assign _1461_ = (_1354_ ? _1445_ : _1460_);
	assign _1462_ = (\mchip.state [0] ? \mchip.internal [31] : \mchip.internal [30]);
	assign _1463_ = (\mchip.state [0] ? \mchip.internal [29] : \mchip.internal [28]);
	assign _1464_ = (\mchip.state [1] ? _1463_ : _1462_);
	assign _1465_ = (\mchip.state [0] ? \mchip.internal [27] : \mchip.internal [26]);
	assign _1466_ = (\mchip.state [0] ? \mchip.internal [25] : \mchip.internal [24]);
	assign _1467_ = (\mchip.state [1] ? _1466_ : _1465_);
	assign _1468_ = (_1345_ ? _1464_ : _1467_);
	assign _1469_ = (\mchip.state [0] ? \mchip.internal [23] : \mchip.internal [22]);
	assign _1470_ = (\mchip.state [0] ? \mchip.internal [21] : \mchip.internal [20]);
	assign _1471_ = (\mchip.state [1] ? _1470_ : _1469_);
	assign _1472_ = (\mchip.state [0] ? \mchip.internal [19] : \mchip.internal [18]);
	assign _1473_ = (\mchip.state [0] ? \mchip.internal [17] : \mchip.internal [16]);
	assign _1474_ = (\mchip.state [1] ? _1473_ : _1472_);
	assign _1475_ = (_1345_ ? _1471_ : _1474_);
	assign _1476_ = (_1347_ ? _1468_ : _1475_);
	assign _1477_ = (\mchip.state [0] ? \mchip.internal [15] : \mchip.internal [14]);
	assign _1478_ = (\mchip.state [0] ? \mchip.internal [13] : \mchip.internal [12]);
	assign _1479_ = (\mchip.state [1] ? _1478_ : _1477_);
	assign _1480_ = (\mchip.state [0] ? \mchip.internal [11] : \mchip.internal [10]);
	assign _1481_ = (\mchip.state [0] ? \mchip.internal [9] : \mchip.internal [8]);
	assign _1482_ = (\mchip.state [1] ? _1481_ : _1480_);
	assign _1483_ = (_1345_ ? _1479_ : _1482_);
	assign _1484_ = (\mchip.state [0] ? \mchip.internal [7] : \mchip.internal [6]);
	assign _1485_ = (\mchip.state [0] ? \mchip.internal [5] : \mchip.internal [4]);
	assign _1486_ = (\mchip.state [1] ? _1485_ : _1484_);
	assign _1487_ = (\mchip.state [0] ? \mchip.internal [3] : \mchip.internal [2]);
	assign _1488_ = (\mchip.state [0] ? \mchip.internal [1] : \mchip.internal [0]);
	assign _1489_ = (\mchip.state [1] ? _1488_ : _1487_);
	assign _1490_ = (_1345_ ? _1486_ : _1489_);
	assign _1491_ = (_1347_ ? _1483_ : _1490_);
	assign _1492_ = (_1354_ ? _1476_ : _1491_);
	assign _1493_ = (_1360_ ? _1461_ : _1492_);
	assign _1494_ = (_1364_ ? _1430_ : _1493_);
	assign _1495_ = _1366_ | ~_1494_;
	assign _1496_ = _1366_ | _1364_;
	assign _1497_ = _1496_ | _1361_;
	assign _1498_ = _1351_ & ~_1497_;
	assign _1499_ = ~(_1498_ ^ _1366_);
	assign _1500_ = _1495_ | ~_1499_;
	assign _1501_ = _1500_ | \mchip.state [0];
	assign _1502_ = ~(\mchip.state [0] ^ \mchip.state [1]);
	assign _1503_ = ~_1502_;
	assign _1504_ = _1503_ | _1501_;
	assign _1505_ = _1349_ ^ _1345_;
	assign _1506_ = ~_1505_;
	assign _1507_ = _1506_ | _1504_;
	assign _1508_ = _1349_ & ~_1345_;
	assign _1509_ = ~(_1508_ ^ _1347_);
	assign _1510_ = _1509_ | _1507_;
	assign _1511_ = ~(_1354_ ^ _1351_);
	assign _1512_ = ~_1511_;
	assign _1513_ = _1512_ | _1510_;
	assign _1514_ = _1351_ & ~_1354_;
	assign _1515_ = ~(_1514_ ^ _1360_);
	assign _1516_ = ~_1515_;
	assign _1517_ = _1516_ | _1513_;
	assign _1518_ = ~(_1364_ ^ _1362_);
	assign _1519_ = ~_1518_;
	assign _1520_ = _1519_ | _1517_;
	assign _1521_ = _1367_ & ~_1520_;
	assign _1522_ = _1498_ | _1366_;
	assign _1523_ = _1522_ | \mchip.state [0];
	assign _1524_ = _1523_ | ~_1502_;
	assign _1525_ = _1524_ | _1506_;
	assign _1526_ = _1525_ | _1509_;
	assign _1527_ = _1526_ | _1512_;
	assign _1528_ = _1527_ | _1516_;
	assign _1529_ = _1528_ | _1519_;
	assign _1530_ = _1367_ & ~_1529_;
	assign _1531_ = _1343_ & ~_1530_;
	assign _1532_ = _1531_ | _1521_;
	assign _1533_ = ~(_1349_ & _1322_);
	assign _1534_ = _1339_ & ~_1533_;
	assign _1535_ = \mchip.state [0] & \mchip.state [1];
	assign _1536_ = _1322_ & ~_1535_;
	assign _1537_ = _1321_ & ~_1536_;
	assign _1538_ = _1338_ & ~_1537_;
	assign _1539_ = \mchip.state [5] & ~_1538_;
	assign _1540_ = _1539_ | \mchip.state [6];
	assign _1541_ = _1540_ | _1534_;
	assign _1542_ = _1533_ | _1331_;
	assign _1543_ = _1330_ & ~_1537_;
	assign _1544_ = _1320_ & ~_1543_;
	assign _1545_ = _1544_ | \mchip.state [6];
	assign _1546_ = _1542_ & ~_1545_;
	assign _1547_ = _1546_ | _1541_;
	assign _0039_ = (_1547_ ? _1343_ : _1532_);
	assign _1548_ = \mchip.key [15] ^ \mchip.plaintext [15];
	assign _1549_ = (_1342_ ? \mchip.internal [15] : _1548_);
	assign _1550_ = _1500_ | _1309_;
	assign _1551_ = _1550_ | _1502_;
	assign _1552_ = _1551_ | _1506_;
	assign _1553_ = _1552_ | _1509_;
	assign _1554_ = _1553_ | _1512_;
	assign _1555_ = _1554_ | _1516_;
	assign _1556_ = _1555_ | _1519_;
	assign _1557_ = _1367_ & ~_1556_;
	assign _1558_ = _1522_ | _1309_;
	assign _1559_ = _1558_ | _1502_;
	assign _1560_ = _1559_ | _1506_;
	assign _1561_ = _1560_ | _1509_;
	assign _1562_ = _1561_ | _1512_;
	assign _1563_ = _1562_ | _1516_;
	assign _1564_ = _1563_ | _1519_;
	assign _1565_ = _1367_ & ~_1564_;
	assign _1566_ = _1549_ & ~_1565_;
	assign _1567_ = _1566_ | _1557_;
	assign _0040_ = (_1547_ ? _1549_ : _1567_);
	assign _1568_ = \mchip.key [16] ^ \mchip.plaintext [16];
	assign _1569_ = (_1342_ ? \mchip.internal [16] : _1568_);
	assign _1570_ = _1502_ | _1501_;
	assign _1571_ = _1570_ | _1506_;
	assign _1572_ = _1571_ | _1509_;
	assign _1573_ = _1572_ | _1512_;
	assign _1574_ = _1573_ | _1516_;
	assign _1575_ = _1574_ | _1519_;
	assign _1576_ = _1367_ & ~_1575_;
	assign _1577_ = _1523_ | _1502_;
	assign _1578_ = _1577_ | _1506_;
	assign _1579_ = _1578_ | _1509_;
	assign _1580_ = _1579_ | _1512_;
	assign _1581_ = _1580_ | _1516_;
	assign _1582_ = _1581_ | _1519_;
	assign _1583_ = _1367_ & ~_1582_;
	assign _1584_ = _1569_ & ~_1583_;
	assign _1585_ = _1584_ | _1576_;
	assign _0041_ = (_1547_ ? _1569_ : _1585_);
	assign _1586_ = \mchip.key [17] ^ \mchip.plaintext [17];
	assign _1587_ = (_1342_ ? \mchip.internal [17] : _1586_);
	assign _1588_ = ~_1509_;
	assign _1589_ = _1550_ | _1503_;
	assign _1590_ = _1589_ | _1505_;
	assign _1591_ = _1590_ | _1588_;
	assign _1592_ = _1591_ | _1511_;
	assign _1593_ = _1592_ | _1516_;
	assign _1594_ = _1593_ | _1519_;
	assign _1595_ = _1367_ & ~_1594_;
	assign _1596_ = _1558_ | ~_1502_;
	assign _1597_ = _1596_ | ~_1506_;
	assign _1598_ = _1597_ | _1588_;
	assign _1599_ = _1598_ | _1511_;
	assign _1600_ = _1599_ | _1516_;
	assign _1601_ = _1600_ | _1519_;
	assign _1602_ = _1367_ & ~_1601_;
	assign _1603_ = _1587_ & ~_1602_;
	assign _1604_ = _1603_ | _1595_;
	assign _0042_ = (_1547_ ? _1587_ : _1604_);
	assign _1605_ = \mchip.key [18] ^ \mchip.plaintext [18];
	assign _1606_ = (_1342_ ? \mchip.internal [18] : _1605_);
	assign _1607_ = _1505_ | _1504_;
	assign _1608_ = _1607_ | _1588_;
	assign _1609_ = _1608_ | _1511_;
	assign _1610_ = _1609_ | _1516_;
	assign _1611_ = _1610_ | _1519_;
	assign _1612_ = _1367_ & ~_1611_;
	assign _1613_ = _1524_ | ~_1506_;
	assign _1614_ = _1613_ | _1588_;
	assign _1615_ = _1614_ | _1511_;
	assign _1616_ = _1615_ | _1516_;
	assign _1617_ = _1616_ | _1519_;
	assign _1618_ = _1367_ & ~_1617_;
	assign _1619_ = _1606_ & ~_1618_;
	assign _1620_ = _1619_ | _1612_;
	assign _0043_ = (_1547_ ? _1606_ : _1620_);
	assign _1621_ = \mchip.key [19] ^ \mchip.plaintext [19];
	assign _1622_ = (_1342_ ? \mchip.internal [19] : _1621_);
	assign _1623_ = _1551_ | _1505_;
	assign _1624_ = _1623_ | _1588_;
	assign _1625_ = _1624_ | _1511_;
	assign _1626_ = _1625_ | _1516_;
	assign _1627_ = _1626_ | _1519_;
	assign _1628_ = _1367_ & ~_1627_;
	assign _1629_ = _1559_ | ~_1506_;
	assign _1630_ = _1629_ | _1588_;
	assign _1631_ = _1630_ | _1511_;
	assign _1632_ = _1631_ | _1516_;
	assign _1633_ = _1632_ | _1519_;
	assign _1634_ = _1367_ & ~_1633_;
	assign _1635_ = _1622_ & ~_1634_;
	assign _1636_ = _1635_ | _1628_;
	assign _0044_ = (_1547_ ? _1622_ : _1636_);
	assign _1637_ = \mchip.key [20] ^ \mchip.plaintext [20];
	assign _1638_ = (_1342_ ? \mchip.internal [20] : _1637_);
	assign _1639_ = _1570_ | _1505_;
	assign _1640_ = _1639_ | _1588_;
	assign _1641_ = _1640_ | _1511_;
	assign _1642_ = _1641_ | _1516_;
	assign _1643_ = _1642_ | _1519_;
	assign _1644_ = _1367_ & ~_1643_;
	assign _1645_ = _1577_ | ~_1506_;
	assign _1646_ = _1645_ | _1588_;
	assign _1647_ = _1646_ | _1511_;
	assign _1648_ = _1647_ | _1516_;
	assign _1649_ = _1648_ | _1519_;
	assign _1650_ = _1367_ & ~_1649_;
	assign _1651_ = _1638_ & ~_1650_;
	assign _1652_ = _1651_ | _1644_;
	assign _0046_ = (_1547_ ? _1638_ : _1652_);
	assign _1653_ = \mchip.key [21] ^ \mchip.plaintext [21];
	assign _1654_ = (_1342_ ? \mchip.internal [21] : _1653_);
	assign _1655_ = _1589_ | _1506_;
	assign _1656_ = _1655_ | _1588_;
	assign _1657_ = _1656_ | _1511_;
	assign _1658_ = _1657_ | _1516_;
	assign _1659_ = _1658_ | _1519_;
	assign _1660_ = _1367_ & ~_1659_;
	assign _1661_ = _1596_ | _1506_;
	assign _1662_ = _1661_ | _1588_;
	assign _1663_ = _1662_ | _1511_;
	assign _1664_ = _1663_ | _1516_;
	assign _1665_ = _1664_ | _1519_;
	assign _1666_ = _1367_ & ~_1665_;
	assign _1667_ = _1654_ & ~_1666_;
	assign _1668_ = _1667_ | _1660_;
	assign _0047_ = (_1547_ ? _1654_ : _1668_);
	assign _1669_ = \mchip.key [22] ^ \mchip.plaintext [22];
	assign _1670_ = (_1342_ ? \mchip.internal [22] : _1669_);
	assign _1671_ = _1588_ | _1507_;
	assign _1672_ = _1671_ | _1511_;
	assign _1673_ = _1672_ | _1516_;
	assign _1674_ = _1673_ | _1519_;
	assign _1675_ = _1367_ & ~_1674_;
	assign _1676_ = _1525_ | _1588_;
	assign _1677_ = _1676_ | _1511_;
	assign _1678_ = _1677_ | _1516_;
	assign _1679_ = _1678_ | _1519_;
	assign _1680_ = _1367_ & ~_1679_;
	assign _1681_ = _1670_ & ~_1680_;
	assign _1682_ = _1681_ | _1675_;
	assign _0048_ = (_1547_ ? _1670_ : _1682_);
	assign _1683_ = \mchip.key [23] ^ \mchip.plaintext [23];
	assign _1684_ = (_1342_ ? \mchip.internal [23] : _1683_);
	assign _1685_ = _1552_ | _1588_;
	assign _1686_ = _1685_ | _1511_;
	assign _1687_ = _1686_ | _1516_;
	assign _1688_ = _1687_ | _1519_;
	assign _1689_ = _1367_ & ~_1688_;
	assign _1690_ = _1560_ | _1588_;
	assign _1691_ = _1690_ | _1511_;
	assign _1692_ = _1691_ | _1516_;
	assign _1693_ = _1692_ | _1519_;
	assign _1694_ = _1367_ & ~_1693_;
	assign _1695_ = _1684_ & ~_1694_;
	assign _1696_ = _1695_ | _1689_;
	assign _0049_ = (_1547_ ? _1684_ : _1696_);
	assign _1697_ = \mchip.key [24] ^ \mchip.plaintext [24];
	assign _1698_ = (_1342_ ? \mchip.internal [24] : _1697_);
	assign _1699_ = _1571_ | _1588_;
	assign _1700_ = _1699_ | _1511_;
	assign _1701_ = _1700_ | _1516_;
	assign _1702_ = _1701_ | _1519_;
	assign _1703_ = _1367_ & ~_1702_;
	assign _1704_ = _1578_ | _1588_;
	assign _1705_ = _1704_ | _1511_;
	assign _1706_ = _1705_ | _1516_;
	assign _1707_ = _1706_ | _1519_;
	assign _1708_ = _1367_ & ~_1707_;
	assign _1709_ = _1698_ & ~_1708_;
	assign _1710_ = _1709_ | _1703_;
	assign _0050_ = (_1547_ ? _1698_ : _1710_);
	assign _1711_ = \mchip.key [25] ^ \mchip.plaintext [25];
	assign _1712_ = (_1342_ ? \mchip.internal [25] : _1711_);
	assign _1713_ = _1590_ | _1509_;
	assign _1714_ = _1713_ | _1511_;
	assign _1715_ = _1714_ | _1516_;
	assign _1716_ = _1715_ | _1519_;
	assign _1717_ = _1367_ & ~_1716_;
	assign _1718_ = _1597_ | _1509_;
	assign _1719_ = _1718_ | _1511_;
	assign _1720_ = _1719_ | _1516_;
	assign _1721_ = _1720_ | _1519_;
	assign _1722_ = _1367_ & ~_1721_;
	assign _1723_ = _1712_ & ~_1722_;
	assign _1724_ = _1723_ | _1717_;
	assign _0051_ = (_1547_ ? _1712_ : _1724_);
	assign _1725_ = \mchip.key [26] ^ \mchip.plaintext [26];
	assign _1726_ = (_1342_ ? \mchip.internal [26] : _1725_);
	assign _1727_ = _1607_ | _1509_;
	assign _1728_ = _1727_ | _1511_;
	assign _1729_ = _1728_ | _1516_;
	assign _1730_ = _1729_ | _1519_;
	assign _1731_ = _1367_ & ~_1730_;
	assign _1732_ = _1613_ | _1509_;
	assign _1733_ = _1732_ | _1511_;
	assign _1734_ = _1733_ | _1516_;
	assign _1735_ = _1734_ | _1519_;
	assign _1736_ = _1367_ & ~_1735_;
	assign _1737_ = _1726_ & ~_1736_;
	assign _1738_ = _1737_ | _1731_;
	assign _0052_ = (_1547_ ? _1726_ : _1738_);
	assign _1739_ = \mchip.key [27] ^ \mchip.plaintext [27];
	assign _0142_ = (_1342_ ? \mchip.internal [27] : _1739_);
	assign _0143_ = _1623_ | _1509_;
	assign _0144_ = _0143_ | _1511_;
	assign _0145_ = _0144_ | _1516_;
	assign _0146_ = _0145_ | _1519_;
	assign _0147_ = _1367_ & ~_0146_;
	assign _0148_ = _1629_ | _1509_;
	assign _0149_ = _0148_ | _1511_;
	assign _0150_ = _0149_ | _1516_;
	assign _0151_ = _0150_ | _1519_;
	assign _0152_ = _1367_ & ~_0151_;
	assign _0153_ = _0142_ & ~_0152_;
	assign _0154_ = _0153_ | _0147_;
	assign _0053_ = (_1547_ ? _0142_ : _0154_);
	assign _0155_ = \mchip.key [28] ^ \mchip.plaintext [28];
	assign _0156_ = (_1342_ ? \mchip.internal [28] : _0155_);
	assign _0157_ = _1639_ | _1509_;
	assign _0158_ = _0157_ | _1511_;
	assign _0159_ = _0158_ | _1516_;
	assign _0160_ = _0159_ | _1519_;
	assign _0161_ = _1367_ & ~_0160_;
	assign _0162_ = _1645_ | _1509_;
	assign _0163_ = _0162_ | _1511_;
	assign _0164_ = _0163_ | _1516_;
	assign _0165_ = _0164_ | _1519_;
	assign _0166_ = _1367_ & ~_0165_;
	assign _0167_ = _0156_ & ~_0166_;
	assign _0168_ = _0167_ | _0161_;
	assign _0054_ = (_1547_ ? _0156_ : _0168_);
	assign _0169_ = \mchip.key [29] ^ \mchip.plaintext [29];
	assign _0170_ = (_1342_ ? \mchip.internal [29] : _0169_);
	assign _0171_ = _1655_ | _1509_;
	assign _0172_ = _0171_ | _1511_;
	assign _0173_ = _0172_ | _1516_;
	assign _0174_ = _0173_ | _1519_;
	assign _0175_ = _1367_ & ~_0174_;
	assign _0176_ = _1661_ | _1509_;
	assign _0177_ = _0176_ | _1511_;
	assign _0178_ = _0177_ | _1516_;
	assign _0179_ = _0178_ | _1519_;
	assign _0180_ = _1367_ & ~_0179_;
	assign _0181_ = _0170_ & ~_0180_;
	assign _0182_ = _0181_ | _0175_;
	assign _0055_ = (_1547_ ? _0170_ : _0182_);
	assign _0183_ = \mchip.key [30] ^ \mchip.plaintext [30];
	assign _0184_ = (_1342_ ? \mchip.internal [30] : _0183_);
	assign _0185_ = _1511_ | _1510_;
	assign _0186_ = _0185_ | _1516_;
	assign _0187_ = _0186_ | _1519_;
	assign _0188_ = _1367_ & ~_0187_;
	assign _0189_ = _1526_ | _1511_;
	assign _0190_ = _0189_ | _1516_;
	assign _0191_ = _0190_ | _1519_;
	assign _0192_ = _1367_ & ~_0191_;
	assign _0193_ = _0184_ & ~_0192_;
	assign _0194_ = _0193_ | _0188_;
	assign _0057_ = (_1547_ ? _0184_ : _0194_);
	assign _0195_ = \mchip.key [31] ^ \mchip.plaintext [31];
	assign _0196_ = (_1342_ ? \mchip.internal [31] : _0195_);
	assign _0197_ = _1553_ | _1511_;
	assign _0198_ = _0197_ | _1516_;
	assign _0199_ = _0198_ | _1519_;
	assign _0200_ = _1367_ & ~_0199_;
	assign _0201_ = _1561_ | _1511_;
	assign _0202_ = _0201_ | _1516_;
	assign _0203_ = _0202_ | _1519_;
	assign _0204_ = _1367_ & ~_0203_;
	assign _0205_ = _0196_ & ~_0204_;
	assign _0206_ = _0205_ | _0200_;
	assign _0058_ = (_1547_ ? _0196_ : _0206_);
	assign _0207_ = \mchip.key [32] ^ \mchip.plaintext [32];
	assign _0208_ = (_1342_ ? \mchip.internal [32] : _0207_);
	assign _0209_ = _1572_ | _1511_;
	assign _0210_ = _0209_ | _1516_;
	assign _0211_ = _0210_ | _1519_;
	assign _0212_ = _1367_ & ~_0211_;
	assign _0213_ = _1579_ | _1511_;
	assign _0214_ = _0213_ | _1516_;
	assign _0215_ = _0214_ | _1519_;
	assign _0216_ = _1367_ & ~_0215_;
	assign _0217_ = _0208_ & ~_0216_;
	assign _0218_ = _0217_ | _0212_;
	assign _0059_ = (_1547_ ? _0208_ : _0218_);
	assign _0219_ = \mchip.key [33] ^ \mchip.plaintext [33];
	assign _0220_ = (_1342_ ? \mchip.internal [33] : _0219_);
	assign _0221_ = _1591_ | _1512_;
	assign _0222_ = _0221_ | _1515_;
	assign _0223_ = _0222_ | _1519_;
	assign _0224_ = _1367_ & ~_0223_;
	assign _0225_ = _1598_ | _1512_;
	assign _0226_ = _0225_ | _1515_;
	assign _0227_ = _0226_ | _1519_;
	assign _0228_ = _1367_ & ~_0227_;
	assign _0229_ = _0220_ & ~_0228_;
	assign _0230_ = _0229_ | _0224_;
	assign _0060_ = (_1547_ ? _0220_ : _0230_);
	assign _0231_ = \mchip.key [34] ^ \mchip.plaintext [34];
	assign _0232_ = (_1342_ ? \mchip.internal [34] : _0231_);
	assign _0233_ = _1608_ | _1512_;
	assign _0234_ = _0233_ | _1515_;
	assign _0235_ = _0234_ | _1519_;
	assign _0236_ = _1367_ & ~_0235_;
	assign _0237_ = _1614_ | _1512_;
	assign _0238_ = _0237_ | _1515_;
	assign _0239_ = _0238_ | _1519_;
	assign _0240_ = _1367_ & ~_0239_;
	assign _0241_ = _0232_ & ~_0240_;
	assign _0242_ = _0241_ | _0236_;
	assign _0061_ = (_1547_ ? _0232_ : _0242_);
	assign _0243_ = \mchip.key [35] ^ \mchip.plaintext [35];
	assign _0244_ = (_1342_ ? \mchip.internal [35] : _0243_);
	assign _0245_ = _1624_ | _1512_;
	assign _0246_ = _0245_ | _1515_;
	assign _0247_ = _0246_ | _1519_;
	assign _0248_ = _1367_ & ~_0247_;
	assign _0249_ = _1630_ | _1512_;
	assign _0250_ = _0249_ | _1515_;
	assign _0251_ = _0250_ | _1519_;
	assign _0252_ = _1367_ & ~_0251_;
	assign _0253_ = _0244_ & ~_0252_;
	assign _0254_ = _0253_ | _0248_;
	assign _0062_ = (_1547_ ? _0244_ : _0254_);
	assign _0255_ = \mchip.key [36] ^ \mchip.plaintext [36];
	assign _0256_ = (_1342_ ? \mchip.internal [36] : _0255_);
	assign _0257_ = _1640_ | _1512_;
	assign _0258_ = _0257_ | _1515_;
	assign _0259_ = _0258_ | _1519_;
	assign _0260_ = _1367_ & ~_0259_;
	assign _0261_ = _1646_ | _1512_;
	assign _0262_ = _0261_ | _1515_;
	assign _0263_ = _0262_ | _1519_;
	assign _0264_ = _1367_ & ~_0263_;
	assign _0265_ = _0256_ & ~_0264_;
	assign _0266_ = _0265_ | _0260_;
	assign _0063_ = (_1547_ ? _0256_ : _0266_);
	assign _0267_ = \mchip.key [37] ^ \mchip.plaintext [37];
	assign _0268_ = (_1342_ ? \mchip.internal [37] : _0267_);
	assign _0269_ = _1656_ | _1512_;
	assign _0270_ = _0269_ | _1515_;
	assign _0271_ = _0270_ | _1519_;
	assign _0272_ = _1367_ & ~_0271_;
	assign _0273_ = _1662_ | _1512_;
	assign _0274_ = _0273_ | _1515_;
	assign _0275_ = _0274_ | _1519_;
	assign _0276_ = _1367_ & ~_0275_;
	assign _0277_ = _0268_ & ~_0276_;
	assign _0278_ = _0277_ | _0272_;
	assign _0064_ = (_1547_ ? _0268_ : _0278_);
	assign _0279_ = \mchip.key [38] ^ \mchip.plaintext [38];
	assign _0280_ = (_1342_ ? \mchip.internal [38] : _0279_);
	assign _0281_ = _1671_ | _1512_;
	assign _0282_ = _0281_ | _1515_;
	assign _0283_ = _0282_ | _1519_;
	assign _0284_ = _1367_ & ~_0283_;
	assign _0285_ = _1676_ | _1512_;
	assign _0286_ = _0285_ | _1515_;
	assign _0287_ = _0286_ | _1519_;
	assign _0288_ = _1367_ & ~_0287_;
	assign _0289_ = _0280_ & ~_0288_;
	assign _0290_ = _0289_ | _0284_;
	assign _0065_ = (_1547_ ? _0280_ : _0290_);
	assign _0291_ = \mchip.key [39] ^ \mchip.plaintext [39];
	assign _0292_ = (_1342_ ? \mchip.internal [39] : _0291_);
	assign _0293_ = _1685_ | _1512_;
	assign _0294_ = _0293_ | _1515_;
	assign _0295_ = _0294_ | _1519_;
	assign _0296_ = _1367_ & ~_0295_;
	assign _0297_ = _1690_ | _1512_;
	assign _0298_ = _0297_ | _1515_;
	assign _0299_ = _0298_ | _1519_;
	assign _0300_ = _1367_ & ~_0299_;
	assign _0301_ = _0292_ & ~_0300_;
	assign _0302_ = _0301_ | _0296_;
	assign _0066_ = (_1547_ ? _0292_ : _0302_);
	assign _0303_ = \mchip.key [40] ^ \mchip.plaintext [40];
	assign _0304_ = (_1342_ ? \mchip.internal [40] : _0303_);
	assign _0305_ = _1699_ | _1512_;
	assign _0306_ = _0305_ | _1515_;
	assign _0307_ = _0306_ | _1519_;
	assign _0308_ = _1367_ & ~_0307_;
	assign _0309_ = _1704_ | _1512_;
	assign _0310_ = _0309_ | _1515_;
	assign _0311_ = _0310_ | _1519_;
	assign _0312_ = _1367_ & ~_0311_;
	assign _0313_ = _0304_ & ~_0312_;
	assign _0314_ = _0313_ | _0308_;
	assign _0068_ = (_1547_ ? _0304_ : _0314_);
	assign _0315_ = \mchip.key [41] ^ \mchip.plaintext [41];
	assign _0316_ = (_1342_ ? \mchip.internal [41] : _0315_);
	assign _0317_ = _1713_ | _1512_;
	assign _0318_ = _0317_ | _1515_;
	assign _0319_ = _0318_ | _1519_;
	assign _0320_ = _1367_ & ~_0319_;
	assign _0321_ = _1718_ | _1512_;
	assign _0322_ = _0321_ | _1515_;
	assign _0323_ = _0322_ | _1519_;
	assign _0324_ = _1367_ & ~_0323_;
	assign _0325_ = _0316_ & ~_0324_;
	assign _0326_ = _0325_ | _0320_;
	assign _0069_ = (_1547_ ? _0316_ : _0326_);
	assign _0327_ = \mchip.key [42] ^ \mchip.plaintext [42];
	assign _0328_ = (_1342_ ? \mchip.internal [42] : _0327_);
	assign _0329_ = _1727_ | _1512_;
	assign _0330_ = _0329_ | _1515_;
	assign _0331_ = _0330_ | _1519_;
	assign _0332_ = _1367_ & ~_0331_;
	assign _0333_ = _1732_ | _1512_;
	assign _0334_ = _0333_ | _1515_;
	assign _0335_ = _0334_ | _1519_;
	assign _0336_ = _1367_ & ~_0335_;
	assign _0337_ = _0328_ & ~_0336_;
	assign _0338_ = _0337_ | _0332_;
	assign _0070_ = (_1547_ ? _0328_ : _0338_);
	assign _0339_ = \mchip.key [43] ^ \mchip.plaintext [43];
	assign _0340_ = (_1342_ ? \mchip.internal [43] : _0339_);
	assign _0341_ = _0143_ | _1512_;
	assign _0342_ = _0341_ | _1515_;
	assign _0343_ = _0342_ | _1519_;
	assign _0344_ = _1367_ & ~_0343_;
	assign _0345_ = _0148_ | _1512_;
	assign _0346_ = _0345_ | _1515_;
	assign _0347_ = _0346_ | _1519_;
	assign _0348_ = _1367_ & ~_0347_;
	assign _0349_ = _0340_ & ~_0348_;
	assign _0350_ = _0349_ | _0344_;
	assign _0071_ = (_1547_ ? _0340_ : _0350_);
	assign _0351_ = \mchip.key [44] ^ \mchip.plaintext [44];
	assign _0352_ = (_1342_ ? \mchip.internal [44] : _0351_);
	assign _0353_ = _0157_ | _1512_;
	assign _0354_ = _0353_ | _1515_;
	assign _0355_ = _0354_ | _1519_;
	assign _0356_ = _1367_ & ~_0355_;
	assign _0357_ = _0162_ | _1512_;
	assign _0358_ = _0357_ | _1515_;
	assign _0359_ = _0358_ | _1519_;
	assign _0360_ = _1367_ & ~_0359_;
	assign _0361_ = _0352_ & ~_0360_;
	assign _0362_ = _0361_ | _0356_;
	assign _0072_ = (_1547_ ? _0352_ : _0362_);
	assign _0363_ = \mchip.key [45] ^ \mchip.plaintext [45];
	assign _0364_ = (_1342_ ? \mchip.internal [45] : _0363_);
	assign _0365_ = _0171_ | _1512_;
	assign _0366_ = _0365_ | _1515_;
	assign _0367_ = _0366_ | _1519_;
	assign _0368_ = _1367_ & ~_0367_;
	assign _0369_ = _0176_ | _1512_;
	assign _0370_ = _0369_ | _1515_;
	assign _0371_ = _0370_ | _1519_;
	assign _0372_ = _1367_ & ~_0371_;
	assign _0373_ = _0364_ & ~_0372_;
	assign _0374_ = _0373_ | _0368_;
	assign _0073_ = (_1547_ ? _0364_ : _0374_);
	assign _0375_ = \mchip.key [46] ^ \mchip.plaintext [46];
	assign _0376_ = (_1342_ ? \mchip.internal [46] : _0375_);
	assign _0377_ = _1515_ | _1513_;
	assign _0378_ = _0377_ | _1519_;
	assign _0379_ = _1367_ & ~_0378_;
	assign _0380_ = _1527_ | _1515_;
	assign _0381_ = _0380_ | _1519_;
	assign _0382_ = _1367_ & ~_0381_;
	assign _0383_ = _0376_ & ~_0382_;
	assign _0384_ = _0383_ | _0379_;
	assign _0074_ = (_1547_ ? _0376_ : _0384_);
	assign _0385_ = \mchip.key [47] ^ \mchip.plaintext [47];
	assign _0386_ = (_1342_ ? \mchip.internal [47] : _0385_);
	assign _0387_ = _1554_ | _1515_;
	assign _0388_ = _0387_ | _1519_;
	assign _0389_ = _1367_ & ~_0388_;
	assign _0390_ = _1562_ | _1515_;
	assign _0391_ = _0390_ | _1519_;
	assign _0392_ = _1367_ & ~_0391_;
	assign _0393_ = _0386_ & ~_0392_;
	assign _0394_ = _0393_ | _0389_;
	assign _0075_ = (_1547_ ? _0386_ : _0394_);
	assign _0395_ = \mchip.key [48] ^ \mchip.plaintext [48];
	assign _0396_ = (_1342_ ? \mchip.internal [48] : _0395_);
	assign _0397_ = _1573_ | _1515_;
	assign _0398_ = _0397_ | _1519_;
	assign _0399_ = _1367_ & ~_0398_;
	assign _0400_ = _1580_ | _1515_;
	assign _0401_ = _0400_ | _1519_;
	assign _0402_ = _1367_ & ~_0401_;
	assign _0403_ = _0396_ & ~_0402_;
	assign _0404_ = _0403_ | _0399_;
	assign _0076_ = (_1547_ ? _0396_ : _0404_);
	assign _0405_ = \mchip.key [49] ^ \mchip.plaintext [49];
	assign _0406_ = (_1342_ ? \mchip.internal [49] : _0405_);
	assign _0407_ = _1592_ | _1515_;
	assign _0408_ = _0407_ | _1519_;
	assign _0409_ = _1367_ & ~_0408_;
	assign _0410_ = _1599_ | _1515_;
	assign _0411_ = _0410_ | _1519_;
	assign _0412_ = _1367_ & ~_0411_;
	assign _0413_ = _0406_ & ~_0412_;
	assign _0414_ = _0413_ | _0409_;
	assign _0077_ = (_1547_ ? _0406_ : _0414_);
	assign _0415_ = \mchip.key [50] ^ \mchip.plaintext [50];
	assign _0416_ = (_1342_ ? \mchip.internal [50] : _0415_);
	assign _0417_ = _1609_ | _1515_;
	assign _0418_ = _0417_ | _1519_;
	assign _0419_ = _1367_ & ~_0418_;
	assign _0420_ = _1615_ | _1515_;
	assign _0421_ = _0420_ | _1519_;
	assign _0422_ = _1367_ & ~_0421_;
	assign _0423_ = _0416_ & ~_0422_;
	assign _0424_ = _0423_ | _0419_;
	assign _0079_ = (_1547_ ? _0416_ : _0424_);
	assign _0425_ = \mchip.key [51] ^ \mchip.plaintext [51];
	assign _0426_ = (_1342_ ? \mchip.internal [51] : _0425_);
	assign _0427_ = _1625_ | _1515_;
	assign _0428_ = _0427_ | _1519_;
	assign _0429_ = _1367_ & ~_0428_;
	assign _0430_ = _1631_ | _1515_;
	assign _0431_ = _0430_ | _1519_;
	assign _0432_ = _1367_ & ~_0431_;
	assign _0433_ = _0426_ & ~_0432_;
	assign _0434_ = _0433_ | _0429_;
	assign _0080_ = (_1547_ ? _0426_ : _0434_);
	assign _0435_ = \mchip.key [52] ^ \mchip.plaintext [52];
	assign _0436_ = (_1342_ ? \mchip.internal [52] : _0435_);
	assign _0437_ = _1641_ | _1515_;
	assign _0438_ = _0437_ | _1519_;
	assign _0439_ = _1367_ & ~_0438_;
	assign _0440_ = _1647_ | _1515_;
	assign _0441_ = _0440_ | _1519_;
	assign _0442_ = _1367_ & ~_0441_;
	assign _0443_ = _0436_ & ~_0442_;
	assign _0444_ = _0443_ | _0439_;
	assign _0081_ = (_1547_ ? _0436_ : _0444_);
	assign _0445_ = \mchip.key [53] ^ \mchip.plaintext [53];
	assign _0446_ = (_1342_ ? \mchip.internal [53] : _0445_);
	assign _0447_ = _1657_ | _1515_;
	assign _0448_ = _0447_ | _1519_;
	assign _0449_ = _1367_ & ~_0448_;
	assign _0450_ = _1663_ | _1515_;
	assign _0451_ = _0450_ | _1519_;
	assign _0452_ = _1367_ & ~_0451_;
	assign _0453_ = _0446_ & ~_0452_;
	assign _0454_ = _0453_ | _0449_;
	assign _0082_ = (_1547_ ? _0446_ : _0454_);
	assign _0455_ = \mchip.key [54] ^ \mchip.plaintext [54];
	assign _0456_ = (_1342_ ? \mchip.internal [54] : _0455_);
	assign _0457_ = _1672_ | _1515_;
	assign _0458_ = _0457_ | _1519_;
	assign _0459_ = _1367_ & ~_0458_;
	assign _0460_ = _1677_ | _1515_;
	assign _0461_ = _0460_ | _1519_;
	assign _0462_ = _1367_ & ~_0461_;
	assign _0463_ = _0456_ & ~_0462_;
	assign _0464_ = _0463_ | _0459_;
	assign _0083_ = (_1547_ ? _0456_ : _0464_);
	assign _0465_ = \mchip.key [55] ^ \mchip.plaintext [55];
	assign _0466_ = (_1342_ ? \mchip.internal [55] : _0465_);
	assign _0467_ = _1686_ | _1515_;
	assign _0468_ = _0467_ | _1519_;
	assign _0469_ = _1367_ & ~_0468_;
	assign _0470_ = _1691_ | _1515_;
	assign _0471_ = _0470_ | _1519_;
	assign _0472_ = _1367_ & ~_0471_;
	assign _0473_ = _0466_ & ~_0472_;
	assign _0474_ = _0473_ | _0469_;
	assign _0084_ = (_1547_ ? _0466_ : _0474_);
	assign _0475_ = \mchip.key [56] ^ \mchip.plaintext [56];
	assign _0476_ = (_1342_ ? \mchip.internal [56] : _0475_);
	assign _0477_ = _1700_ | _1515_;
	assign _0478_ = _0477_ | _1519_;
	assign _0479_ = _1367_ & ~_0478_;
	assign _0480_ = _1705_ | _1515_;
	assign _0481_ = _0480_ | _1519_;
	assign _0482_ = _1367_ & ~_0481_;
	assign _0483_ = _0476_ & ~_0482_;
	assign _0484_ = _0483_ | _0479_;
	assign _0085_ = (_1547_ ? _0476_ : _0484_);
	assign _0485_ = \mchip.key [57] ^ \mchip.plaintext [57];
	assign _0486_ = (_1342_ ? \mchip.internal [57] : _0485_);
	assign _0487_ = _1714_ | _1515_;
	assign _0488_ = _0487_ | _1519_;
	assign _0489_ = _1367_ & ~_0488_;
	assign _0490_ = _1719_ | _1515_;
	assign _0491_ = _0490_ | _1519_;
	assign _0492_ = _1367_ & ~_0491_;
	assign _0493_ = _0486_ & ~_0492_;
	assign _0494_ = _0493_ | _0489_;
	assign _0086_ = (_1547_ ? _0486_ : _0494_);
	assign _0495_ = \mchip.key [58] ^ \mchip.plaintext [58];
	assign _0496_ = (_1342_ ? \mchip.internal [58] : _0495_);
	assign _0497_ = _1728_ | _1515_;
	assign _0498_ = _0497_ | _1519_;
	assign _0499_ = _1367_ & ~_0498_;
	assign _0500_ = _1733_ | _1515_;
	assign _0501_ = _0500_ | _1519_;
	assign _0502_ = _1367_ & ~_0501_;
	assign _0503_ = _0496_ & ~_0502_;
	assign _0504_ = _0503_ | _0499_;
	assign _0087_ = (_1547_ ? _0496_ : _0504_);
	assign _0505_ = \mchip.key [59] ^ \mchip.plaintext [59];
	assign _0506_ = (_1342_ ? \mchip.internal [59] : _0505_);
	assign _0507_ = _0144_ | _1515_;
	assign _0508_ = _0507_ | _1519_;
	assign _0509_ = _1367_ & ~_0508_;
	assign _0510_ = _0149_ | _1515_;
	assign _0511_ = _0510_ | _1519_;
	assign _0512_ = _1367_ & ~_0511_;
	assign _0513_ = _0506_ & ~_0512_;
	assign _0514_ = _0513_ | _0509_;
	assign _0088_ = (_1547_ ? _0506_ : _0514_);
	assign _0515_ = \mchip.key [60] ^ \mchip.plaintext [60];
	assign _0516_ = (_1342_ ? \mchip.internal [60] : _0515_);
	assign _0517_ = _0158_ | _1515_;
	assign _0518_ = _0517_ | _1519_;
	assign _0519_ = _1367_ & ~_0518_;
	assign _0520_ = _0163_ | _1515_;
	assign _0521_ = _0520_ | _1519_;
	assign _0522_ = _1367_ & ~_0521_;
	assign _0523_ = _0516_ & ~_0522_;
	assign _0524_ = _0523_ | _0519_;
	assign _0090_ = (_1547_ ? _0516_ : _0524_);
	assign _0525_ = \mchip.key [61] ^ \mchip.plaintext [61];
	assign _0526_ = (_1342_ ? \mchip.internal [61] : _0525_);
	assign _0527_ = _0172_ | _1515_;
	assign _0528_ = _0527_ | _1519_;
	assign _0529_ = _1367_ & ~_0528_;
	assign _0530_ = _0177_ | _1515_;
	assign _0531_ = _0530_ | _1519_;
	assign _0532_ = _1367_ & ~_0531_;
	assign _0533_ = _0526_ & ~_0532_;
	assign _0534_ = _0533_ | _0529_;
	assign _0091_ = (_1547_ ? _0526_ : _0534_);
	assign _0535_ = \mchip.key [62] ^ \mchip.plaintext [62];
	assign _0536_ = (_1342_ ? \mchip.internal [62] : _0535_);
	assign _0537_ = _0185_ | _1515_;
	assign _0538_ = _0537_ | _1519_;
	assign _0539_ = _1367_ & ~_0538_;
	assign _0540_ = _0189_ | _1515_;
	assign _0541_ = _0540_ | _1519_;
	assign _0542_ = _1367_ & ~_0541_;
	assign _0543_ = _0536_ & ~_0542_;
	assign _0544_ = _0543_ | _0539_;
	assign _0092_ = (_1547_ ? _0536_ : _0544_);
	assign _0545_ = \mchip.key [63] ^ \mchip.plaintext [63];
	assign _0546_ = (_1342_ ? \mchip.internal [63] : _0545_);
	assign _0547_ = _0197_ | _1515_;
	assign _0548_ = _0547_ | _1519_;
	assign _0549_ = _1367_ & ~_0548_;
	assign _0550_ = _0201_ | _1515_;
	assign _0551_ = _0550_ | _1519_;
	assign _0552_ = _1367_ & ~_0551_;
	assign _0553_ = _0546_ & ~_0552_;
	assign _0554_ = _0553_ | _0549_;
	assign _0093_ = (_1547_ ? _0546_ : _0554_);
	assign _0555_ = \mchip.key [64] ^ \mchip.plaintext [64];
	assign _0556_ = (_1342_ ? \mchip.internal [64] : _0555_);
	assign _0557_ = _0209_ | _1515_;
	assign _0558_ = _0557_ | _1519_;
	assign _0559_ = _1367_ & ~_0558_;
	assign _0560_ = _0213_ | _1515_;
	assign _0561_ = _0560_ | _1519_;
	assign _0562_ = _1367_ & ~_0561_;
	assign _0563_ = _0556_ & ~_0562_;
	assign _0564_ = _0563_ | _0559_;
	assign _0094_ = (_1547_ ? _0556_ : _0564_);
	assign _0565_ = \mchip.key [65] ^ \mchip.plaintext [65];
	assign _0566_ = (_1342_ ? \mchip.internal [65] : _0565_);
	assign _0567_ = _0221_ | _1516_;
	assign _0568_ = _0567_ | _1518_;
	assign _0569_ = _1367_ & ~_0568_;
	assign _0570_ = _0225_ | _1516_;
	assign _0571_ = _0570_ | _1518_;
	assign _0572_ = _1367_ & ~_0571_;
	assign _0573_ = _0566_ & ~_0572_;
	assign _0574_ = _0573_ | _0569_;
	assign _0095_ = (_1547_ ? _0566_ : _0574_);
	assign _0575_ = \mchip.key [66] ^ \mchip.plaintext [66];
	assign _0576_ = (_1342_ ? \mchip.internal [66] : _0575_);
	assign _0577_ = _0233_ | _1516_;
	assign _0578_ = _0577_ | _1518_;
	assign _0579_ = _1367_ & ~_0578_;
	assign _0580_ = _0237_ | _1516_;
	assign _0581_ = _0580_ | _1518_;
	assign _0582_ = _1367_ & ~_0581_;
	assign _0583_ = _0576_ & ~_0582_;
	assign _0584_ = _0583_ | _0579_;
	assign _0096_ = (_1547_ ? _0576_ : _0584_);
	assign _0585_ = \mchip.key [67] ^ \mchip.plaintext [67];
	assign _0586_ = (_1342_ ? \mchip.internal [67] : _0585_);
	assign _0587_ = _0245_ | _1516_;
	assign _0588_ = _0587_ | _1518_;
	assign _0589_ = _1367_ & ~_0588_;
	assign _0590_ = _0249_ | _1516_;
	assign _0591_ = _0590_ | _1518_;
	assign _0592_ = _1367_ & ~_0591_;
	assign _0593_ = _0586_ & ~_0592_;
	assign _0594_ = _0593_ | _0589_;
	assign _0097_ = (_1547_ ? _0586_ : _0594_);
	assign _0595_ = \mchip.key [68] ^ \mchip.plaintext [68];
	assign _0596_ = (_1342_ ? \mchip.internal [68] : _0595_);
	assign _0597_ = _0257_ | _1516_;
	assign _0598_ = _0597_ | _1518_;
	assign _0599_ = _1367_ & ~_0598_;
	assign _0600_ = _0261_ | _1516_;
	assign _0601_ = _0600_ | _1518_;
	assign _0602_ = _1367_ & ~_0601_;
	assign _0603_ = _0596_ & ~_0602_;
	assign _0604_ = _0603_ | _0599_;
	assign _0098_ = (_1547_ ? _0596_ : _0604_);
	assign _0605_ = \mchip.key [69] ^ \mchip.plaintext [69];
	assign _0606_ = (_1342_ ? \mchip.internal [69] : _0605_);
	assign _0607_ = _0269_ | _1516_;
	assign _0608_ = _0607_ | _1518_;
	assign _0609_ = _1367_ & ~_0608_;
	assign _0610_ = _0273_ | _1516_;
	assign _0611_ = _0610_ | _1518_;
	assign _0612_ = _1367_ & ~_0611_;
	assign _0613_ = _0606_ & ~_0612_;
	assign _0614_ = _0613_ | _0609_;
	assign _0099_ = (_1547_ ? _0606_ : _0614_);
	assign _0615_ = \mchip.key [70] ^ \mchip.plaintext [70];
	assign _0616_ = (_1342_ ? \mchip.internal [70] : _0615_);
	assign _0617_ = _0281_ | _1516_;
	assign _0618_ = _0617_ | _1518_;
	assign _0619_ = _1367_ & ~_0618_;
	assign _0620_ = _0285_ | _1516_;
	assign _0621_ = _0620_ | _1518_;
	assign _0622_ = _1367_ & ~_0621_;
	assign _0623_ = _0616_ & ~_0622_;
	assign _0624_ = _0623_ | _0619_;
	assign _0101_ = (_1547_ ? _0616_ : _0624_);
	assign _0625_ = \mchip.key [71] ^ \mchip.plaintext [71];
	assign _0626_ = (_1342_ ? \mchip.internal [71] : _0625_);
	assign _0627_ = _0293_ | _1516_;
	assign _0628_ = _0627_ | _1518_;
	assign _0629_ = _1367_ & ~_0628_;
	assign _0630_ = _0297_ | _1516_;
	assign _0631_ = _0630_ | _1518_;
	assign _0632_ = _1367_ & ~_0631_;
	assign _0633_ = _0626_ & ~_0632_;
	assign _0634_ = _0633_ | _0629_;
	assign _0102_ = (_1547_ ? _0626_ : _0634_);
	assign _0635_ = \mchip.key [72] ^ \mchip.plaintext [72];
	assign _0636_ = (_1342_ ? \mchip.internal [72] : _0635_);
	assign _0637_ = _0305_ | _1516_;
	assign _0638_ = _0637_ | _1518_;
	assign _0639_ = _1367_ & ~_0638_;
	assign _0640_ = _0309_ | _1516_;
	assign _0641_ = _0640_ | _1518_;
	assign _0642_ = _1367_ & ~_0641_;
	assign _0643_ = _0636_ & ~_0642_;
	assign _0644_ = _0643_ | _0639_;
	assign _0103_ = (_1547_ ? _0636_ : _0644_);
	assign _0645_ = \mchip.key [73] ^ \mchip.plaintext [73];
	assign _0646_ = (_1342_ ? \mchip.internal [73] : _0645_);
	assign _0647_ = _0317_ | _1516_;
	assign _0648_ = _0647_ | _1518_;
	assign _0649_ = _1367_ & ~_0648_;
	assign _0650_ = _0321_ | _1516_;
	assign _0651_ = _0650_ | _1518_;
	assign _0652_ = _1367_ & ~_0651_;
	assign _0653_ = _0646_ & ~_0652_;
	assign _0654_ = _0653_ | _0649_;
	assign _0104_ = (_1547_ ? _0646_ : _0654_);
	assign _0655_ = \mchip.key [74] ^ \mchip.plaintext [74];
	assign _0656_ = (_1342_ ? \mchip.internal [74] : _0655_);
	assign _0657_ = _0329_ | _1516_;
	assign _0658_ = _0657_ | _1518_;
	assign _0659_ = _1367_ & ~_0658_;
	assign _0660_ = _0333_ | _1516_;
	assign _0661_ = _0660_ | _1518_;
	assign _0662_ = _1367_ & ~_0661_;
	assign _0663_ = _0656_ & ~_0662_;
	assign _0664_ = _0663_ | _0659_;
	assign _0105_ = (_1547_ ? _0656_ : _0664_);
	assign _0665_ = \mchip.key [75] ^ \mchip.plaintext [75];
	assign _0666_ = (_1342_ ? \mchip.internal [75] : _0665_);
	assign _0667_ = _0341_ | _1516_;
	assign _0668_ = _0667_ | _1518_;
	assign _0669_ = _1367_ & ~_0668_;
	assign _0670_ = _0345_ | _1516_;
	assign _0671_ = _0670_ | _1518_;
	assign _0672_ = _1367_ & ~_0671_;
	assign _0673_ = _0666_ & ~_0672_;
	assign _0674_ = _0673_ | _0669_;
	assign _0106_ = (_1547_ ? _0666_ : _0674_);
	assign _0675_ = \mchip.key [76] ^ \mchip.plaintext [76];
	assign _0676_ = (_1342_ ? \mchip.internal [76] : _0675_);
	assign _0677_ = _0353_ | _1516_;
	assign _0678_ = _0677_ | _1518_;
	assign _0679_ = _1367_ & ~_0678_;
	assign _0680_ = _0357_ | _1516_;
	assign _0681_ = _0680_ | _1518_;
	assign _0682_ = _1367_ & ~_0681_;
	assign _0683_ = _0676_ & ~_0682_;
	assign _0684_ = _0683_ | _0679_;
	assign _0107_ = (_1547_ ? _0676_ : _0684_);
	assign _0685_ = \mchip.key [77] ^ \mchip.plaintext [77];
	assign _0686_ = (_1342_ ? \mchip.internal [77] : _0685_);
	assign _0687_ = _0365_ | _1516_;
	assign _0688_ = _0687_ | _1518_;
	assign _0689_ = _1367_ & ~_0688_;
	assign _0690_ = _0369_ | _1516_;
	assign _0691_ = _0690_ | _1518_;
	assign _0692_ = _1367_ & ~_0691_;
	assign _0693_ = _0686_ & ~_0692_;
	assign _0694_ = _0693_ | _0689_;
	assign _0108_ = (_1547_ ? _0686_ : _0694_);
	assign _0695_ = \mchip.key [78] ^ \mchip.plaintext [78];
	assign _0696_ = (_1342_ ? \mchip.internal [78] : _0695_);
	assign _0697_ = _1518_ | _1517_;
	assign _0698_ = _1367_ & ~_0697_;
	assign _0699_ = _1528_ | _1518_;
	assign _0700_ = _1367_ & ~_0699_;
	assign _0701_ = _0696_ & ~_0700_;
	assign _0702_ = _0701_ | _0698_;
	assign _0109_ = (_1547_ ? _0696_ : _0702_);
	assign _0703_ = \mchip.key [79] ^ \mchip.plaintext [79];
	assign _0704_ = (_1342_ ? \mchip.internal [79] : _0703_);
	assign _0705_ = _1555_ | _1518_;
	assign _0706_ = _1367_ & ~_0705_;
	assign _0707_ = _1563_ | _1518_;
	assign _0708_ = _1367_ & ~_0707_;
	assign _0709_ = _0704_ & ~_0708_;
	assign _0710_ = _0709_ | _0706_;
	assign _0110_ = (_1547_ ? _0704_ : _0710_);
	assign _0711_ = \mchip.key [80] ^ \mchip.plaintext [80];
	assign _0712_ = (_1342_ ? \mchip.internal [80] : _0711_);
	assign _0713_ = _1574_ | _1518_;
	assign _0714_ = _1367_ & ~_0713_;
	assign _0715_ = _1581_ | _1518_;
	assign _0716_ = _1367_ & ~_0715_;
	assign _0717_ = _0712_ & ~_0716_;
	assign _0718_ = _0717_ | _0714_;
	assign _0112_ = (_1547_ ? _0712_ : _0718_);
	assign _0719_ = \mchip.key [81] ^ \mchip.plaintext [81];
	assign _0720_ = (_1342_ ? \mchip.internal [81] : _0719_);
	assign _0721_ = _1593_ | _1518_;
	assign _0722_ = _1367_ & ~_0721_;
	assign _0723_ = _1600_ | _1518_;
	assign _0724_ = _1367_ & ~_0723_;
	assign _0725_ = _0720_ & ~_0724_;
	assign _0726_ = _0725_ | _0722_;
	assign _0113_ = (_1547_ ? _0720_ : _0726_);
	assign _0727_ = \mchip.key [82] ^ \mchip.plaintext [82];
	assign _0728_ = (_1342_ ? \mchip.internal [82] : _0727_);
	assign _0729_ = _1610_ | _1518_;
	assign _0730_ = _1367_ & ~_0729_;
	assign _0731_ = _1616_ | _1518_;
	assign _0732_ = _1367_ & ~_0731_;
	assign _0733_ = _0728_ & ~_0732_;
	assign _0734_ = _0733_ | _0730_;
	assign _0114_ = (_1547_ ? _0728_ : _0734_);
	assign _0735_ = \mchip.key [83] ^ \mchip.plaintext [83];
	assign _0736_ = (_1342_ ? \mchip.internal [83] : _0735_);
	assign _0737_ = _1626_ | _1518_;
	assign _0738_ = _1367_ & ~_0737_;
	assign _0739_ = _1632_ | _1518_;
	assign _0740_ = _1367_ & ~_0739_;
	assign _0741_ = _0736_ & ~_0740_;
	assign _0742_ = _0741_ | _0738_;
	assign _0115_ = (_1547_ ? _0736_ : _0742_);
	assign _0743_ = \mchip.key [84] ^ \mchip.plaintext [84];
	assign _0744_ = (_1342_ ? \mchip.internal [84] : _0743_);
	assign _0745_ = _1642_ | _1518_;
	assign _0746_ = _1367_ & ~_0745_;
	assign _0747_ = _1648_ | _1518_;
	assign _0748_ = _1367_ & ~_0747_;
	assign _0749_ = _0744_ & ~_0748_;
	assign _0750_ = _0749_ | _0746_;
	assign _0116_ = (_1547_ ? _0744_ : _0750_);
	assign _0751_ = \mchip.key [85] ^ \mchip.plaintext [85];
	assign _0752_ = (_1342_ ? \mchip.internal [85] : _0751_);
	assign _0753_ = _1658_ | _1518_;
	assign _0754_ = _1367_ & ~_0753_;
	assign _0755_ = _1664_ | _1518_;
	assign _0756_ = _1367_ & ~_0755_;
	assign _0757_ = _0752_ & ~_0756_;
	assign _0758_ = _0757_ | _0754_;
	assign _0117_ = (_1547_ ? _0752_ : _0758_);
	assign _0759_ = \mchip.key [86] ^ \mchip.plaintext [86];
	assign _0760_ = (_1342_ ? \mchip.internal [86] : _0759_);
	assign _0761_ = _1673_ | _1518_;
	assign _0762_ = _1367_ & ~_0761_;
	assign _0763_ = _1678_ | _1518_;
	assign _0764_ = _1367_ & ~_0763_;
	assign _0765_ = _0760_ & ~_0764_;
	assign _0766_ = _0765_ | _0762_;
	assign _0118_ = (_1547_ ? _0760_ : _0766_);
	assign _0767_ = \mchip.key [87] ^ \mchip.plaintext [87];
	assign _0768_ = (_1342_ ? \mchip.internal [87] : _0767_);
	assign _0769_ = _1687_ | _1518_;
	assign _0770_ = _1367_ & ~_0769_;
	assign _0771_ = _1692_ | _1518_;
	assign _0772_ = _1367_ & ~_0771_;
	assign _0773_ = _0768_ & ~_0772_;
	assign _0774_ = _0773_ | _0770_;
	assign _0119_ = (_1547_ ? _0768_ : _0774_);
	assign _0775_ = \mchip.key [88] ^ \mchip.plaintext [88];
	assign _0776_ = (_1342_ ? \mchip.internal [88] : _0775_);
	assign _0777_ = _1701_ | _1518_;
	assign _0778_ = _1367_ & ~_0777_;
	assign _0779_ = _1706_ | _1518_;
	assign _0780_ = _1367_ & ~_0779_;
	assign _0781_ = _0776_ & ~_0780_;
	assign _0782_ = _0781_ | _0778_;
	assign _0120_ = (_1547_ ? _0776_ : _0782_);
	assign _0783_ = \mchip.key [89] ^ \mchip.plaintext [89];
	assign _0784_ = (_1342_ ? \mchip.internal [89] : _0783_);
	assign _0785_ = _1715_ | _1518_;
	assign _0786_ = _1367_ & ~_0785_;
	assign _0787_ = _1720_ | _1518_;
	assign _0788_ = _1367_ & ~_0787_;
	assign _0789_ = _0784_ & ~_0788_;
	assign _0790_ = _0789_ | _0786_;
	assign _0121_ = (_1547_ ? _0784_ : _0790_);
	assign _0791_ = \mchip.key [90] ^ \mchip.plaintext [90];
	assign _0792_ = (_1342_ ? \mchip.internal [90] : _0791_);
	assign _0793_ = _1729_ | _1518_;
	assign _0794_ = _1367_ & ~_0793_;
	assign _0795_ = _1734_ | _1518_;
	assign _0796_ = _1367_ & ~_0795_;
	assign _0797_ = _0792_ & ~_0796_;
	assign _0798_ = _0797_ | _0794_;
	assign _0123_ = (_1547_ ? _0792_ : _0798_);
	assign _0799_ = \mchip.key [91] ^ \mchip.plaintext [91];
	assign _0800_ = (_1342_ ? \mchip.internal [91] : _0799_);
	assign _0801_ = _0145_ | _1518_;
	assign _0802_ = _1367_ & ~_0801_;
	assign _0803_ = _0150_ | _1518_;
	assign _0804_ = _1367_ & ~_0803_;
	assign _0805_ = _0800_ & ~_0804_;
	assign _0806_ = _0805_ | _0802_;
	assign _0124_ = (_1547_ ? _0800_ : _0806_);
	assign _0807_ = \mchip.key [92] ^ \mchip.plaintext [92];
	assign _0808_ = (_1342_ ? \mchip.internal [92] : _0807_);
	assign _0809_ = _0159_ | _1518_;
	assign _0810_ = _1367_ & ~_0809_;
	assign _0811_ = _0164_ | _1518_;
	assign _0812_ = _1367_ & ~_0811_;
	assign _0813_ = _0808_ & ~_0812_;
	assign _0814_ = _0813_ | _0810_;
	assign _0125_ = (_1547_ ? _0808_ : _0814_);
	assign _0815_ = \mchip.key [93] ^ \mchip.plaintext [93];
	assign _0816_ = (_1342_ ? \mchip.internal [93] : _0815_);
	assign _0817_ = _0173_ | _1518_;
	assign _0818_ = _1367_ & ~_0817_;
	assign _0819_ = _0178_ | _1518_;
	assign _0820_ = _1367_ & ~_0819_;
	assign _0821_ = _0816_ & ~_0820_;
	assign _0822_ = _0821_ | _0818_;
	assign _0126_ = (_1547_ ? _0816_ : _0822_);
	assign _0823_ = \mchip.key [94] ^ \mchip.plaintext [94];
	assign _0824_ = (_1342_ ? \mchip.internal [94] : _0823_);
	assign _0825_ = _0186_ | _1518_;
	assign _0826_ = _1367_ & ~_0825_;
	assign _0827_ = _0190_ | _1518_;
	assign _0828_ = _1367_ & ~_0827_;
	assign _0829_ = _0824_ & ~_0828_;
	assign _0830_ = _0829_ | _0826_;
	assign _0127_ = (_1547_ ? _0824_ : _0830_);
	assign _0831_ = \mchip.key [95] ^ \mchip.plaintext [95];
	assign _0832_ = (_1342_ ? \mchip.internal [95] : _0831_);
	assign _0833_ = _0198_ | _1518_;
	assign _0834_ = _1367_ & ~_0833_;
	assign _0835_ = _0202_ | _1518_;
	assign _0836_ = _1367_ & ~_0835_;
	assign _0837_ = _0832_ & ~_0836_;
	assign _0838_ = _0837_ | _0834_;
	assign _0128_ = (_1547_ ? _0832_ : _0838_);
	assign _0839_ = \mchip.key [96] ^ \mchip.plaintext [96];
	assign _0840_ = (_1342_ ? \mchip.internal [96] : _0839_);
	assign _0841_ = _0210_ | _1518_;
	assign _0842_ = _1367_ & ~_0841_;
	assign _0843_ = _0214_ | _1518_;
	assign _0844_ = _1367_ & ~_0843_;
	assign _0845_ = _0840_ & ~_0844_;
	assign _0846_ = _0845_ | _0842_;
	assign _0129_ = (_1547_ ? _0840_ : _0846_);
	assign _0847_ = \mchip.key [97] ^ \mchip.plaintext [97];
	assign _0848_ = (_1342_ ? \mchip.internal [97] : _0847_);
	assign _0849_ = _0222_ | _1518_;
	assign _0850_ = _1367_ & ~_0849_;
	assign _0851_ = _0226_ | _1518_;
	assign _0852_ = _1367_ & ~_0851_;
	assign _0853_ = _0848_ & ~_0852_;
	assign _0854_ = _0853_ | _0850_;
	assign _0130_ = (_1547_ ? _0848_ : _0854_);
	assign _0855_ = \mchip.key [98] ^ \mchip.plaintext [98];
	assign _0856_ = (_1342_ ? \mchip.internal [98] : _0855_);
	assign _0857_ = _0234_ | _1518_;
	assign _0858_ = _1367_ & ~_0857_;
	assign _0859_ = _0238_ | _1518_;
	assign _0860_ = _1367_ & ~_0859_;
	assign _0861_ = _0856_ & ~_0860_;
	assign _0862_ = _0861_ | _0858_;
	assign _0131_ = (_1547_ ? _0856_ : _0862_);
	assign _0863_ = \mchip.key [99] ^ \mchip.plaintext [99];
	assign _0864_ = (_1342_ ? \mchip.internal [99] : _0863_);
	assign _0865_ = _0246_ | _1518_;
	assign _0866_ = _1367_ & ~_0865_;
	assign _0867_ = _0250_ | _1518_;
	assign _0868_ = _1367_ & ~_0867_;
	assign _0869_ = _0864_ & ~_0868_;
	assign _0870_ = _0869_ | _0866_;
	assign _0132_ = (_1547_ ? _0864_ : _0870_);
	assign _0871_ = \mchip.key [100] ^ \mchip.plaintext [100];
	assign _0872_ = (_1342_ ? \mchip.internal [100] : _0871_);
	assign _0873_ = _0258_ | _1518_;
	assign _0874_ = _1367_ & ~_0873_;
	assign _0875_ = _0262_ | _1518_;
	assign _0876_ = _1367_ & ~_0875_;
	assign _0877_ = _0872_ & ~_0876_;
	assign _0878_ = _0877_ | _0874_;
	assign _0007_ = (_1547_ ? _0872_ : _0878_);
	assign _0879_ = \mchip.key [101] ^ \mchip.plaintext [101];
	assign _0880_ = (_1342_ ? \mchip.internal [101] : _0879_);
	assign _0881_ = _0270_ | _1518_;
	assign _0882_ = _1367_ & ~_0881_;
	assign _0883_ = _0274_ | _1518_;
	assign _0884_ = _1367_ & ~_0883_;
	assign _0885_ = _0880_ & ~_0884_;
	assign _0886_ = _0885_ | _0882_;
	assign _0008_ = (_1547_ ? _0880_ : _0886_);
	assign _0887_ = \mchip.key [102] ^ \mchip.plaintext [102];
	assign _0888_ = (_1342_ ? \mchip.internal [102] : _0887_);
	assign _0889_ = _0282_ | _1518_;
	assign _0890_ = _1367_ & ~_0889_;
	assign _0891_ = _0286_ | _1518_;
	assign _0892_ = _1367_ & ~_0891_;
	assign _0893_ = _0888_ & ~_0892_;
	assign _0894_ = _0893_ | _0890_;
	assign _0009_ = (_1547_ ? _0888_ : _0894_);
	assign _0895_ = \mchip.key [103] ^ \mchip.plaintext [103];
	assign _0896_ = (_1342_ ? \mchip.internal [103] : _0895_);
	assign _0897_ = _0294_ | _1518_;
	assign _0898_ = _1367_ & ~_0897_;
	assign _0899_ = _0298_ | _1518_;
	assign _0900_ = _1367_ & ~_0899_;
	assign _0901_ = _0896_ & ~_0900_;
	assign _0902_ = _0901_ | _0898_;
	assign _0010_ = (_1547_ ? _0896_ : _0902_);
	assign _0903_ = \mchip.key [104] ^ \mchip.plaintext [104];
	assign _0904_ = (_1342_ ? \mchip.internal [104] : _0903_);
	assign _0905_ = _0306_ | _1518_;
	assign _0906_ = _1367_ & ~_0905_;
	assign _0907_ = _0310_ | _1518_;
	assign _0908_ = _1367_ & ~_0907_;
	assign _0909_ = _0904_ & ~_0908_;
	assign _0910_ = _0909_ | _0906_;
	assign _0011_ = (_1547_ ? _0904_ : _0910_);
	assign _0911_ = \mchip.key [105] ^ \mchip.plaintext [105];
	assign _0912_ = (_1342_ ? \mchip.internal [105] : _0911_);
	assign _0913_ = _0318_ | _1518_;
	assign _0914_ = _1367_ & ~_0913_;
	assign _0915_ = _0322_ | _1518_;
	assign _0916_ = _1367_ & ~_0915_;
	assign _0917_ = _0912_ & ~_0916_;
	assign _0918_ = _0917_ | _0914_;
	assign _0012_ = (_1547_ ? _0912_ : _0918_);
	assign _0919_ = \mchip.key [106] ^ \mchip.plaintext [106];
	assign _0920_ = (_1342_ ? \mchip.internal [106] : _0919_);
	assign _0921_ = _0330_ | _1518_;
	assign _0922_ = _1367_ & ~_0921_;
	assign _0923_ = _0334_ | _1518_;
	assign _0924_ = _1367_ & ~_0923_;
	assign _0925_ = _0920_ & ~_0924_;
	assign _0926_ = _0925_ | _0922_;
	assign _0013_ = (_1547_ ? _0920_ : _0926_);
	assign _0927_ = \mchip.key [107] ^ \mchip.plaintext [107];
	assign _0928_ = (_1342_ ? \mchip.internal [107] : _0927_);
	assign _0929_ = _0342_ | _1518_;
	assign _0930_ = _1367_ & ~_0929_;
	assign _0931_ = _0346_ | _1518_;
	assign _0932_ = _1367_ & ~_0931_;
	assign _0933_ = _0928_ & ~_0932_;
	assign _0934_ = _0933_ | _0930_;
	assign _0014_ = (_1547_ ? _0928_ : _0934_);
	assign _0935_ = \mchip.key [108] ^ \mchip.plaintext [108];
	assign _0936_ = (_1342_ ? \mchip.internal [108] : _0935_);
	assign _0937_ = _0354_ | _1518_;
	assign _0938_ = _1367_ & ~_0937_;
	assign _0939_ = _0358_ | _1518_;
	assign _0940_ = _1367_ & ~_0939_;
	assign _0941_ = _0936_ & ~_0940_;
	assign _0942_ = _0941_ | _0938_;
	assign _0015_ = (_1547_ ? _0936_ : _0942_);
	assign _0943_ = \mchip.key [109] ^ \mchip.plaintext [109];
	assign _0944_ = (_1342_ ? \mchip.internal [109] : _0943_);
	assign _0945_ = _0366_ | _1518_;
	assign _0946_ = _1367_ & ~_0945_;
	assign _0947_ = _0370_ | _1518_;
	assign _0948_ = _1367_ & ~_0947_;
	assign _0949_ = _0944_ & ~_0948_;
	assign _0950_ = _0949_ | _0946_;
	assign _0016_ = (_1547_ ? _0944_ : _0950_);
	assign _0951_ = \mchip.key [110] ^ \mchip.plaintext [110];
	assign _0952_ = (_1342_ ? \mchip.internal [110] : _0951_);
	assign _0953_ = _0377_ | _1518_;
	assign _0954_ = _1367_ & ~_0953_;
	assign _0955_ = _0380_ | _1518_;
	assign _0956_ = _1367_ & ~_0955_;
	assign _0957_ = _0952_ & ~_0956_;
	assign _0958_ = _0957_ | _0954_;
	assign _0018_ = (_1547_ ? _0952_ : _0958_);
	assign _0959_ = \mchip.key [111] ^ \mchip.plaintext [111];
	assign _0960_ = (_1342_ ? \mchip.internal [111] : _0959_);
	assign _0961_ = _0387_ | _1518_;
	assign _0962_ = _1367_ & ~_0961_;
	assign _0963_ = _0390_ | _1518_;
	assign _0964_ = _1367_ & ~_0963_;
	assign _0965_ = _0960_ & ~_0964_;
	assign _0966_ = _0965_ | _0962_;
	assign _0019_ = (_1547_ ? _0960_ : _0966_);
	assign _0967_ = \mchip.key [112] ^ \mchip.plaintext [112];
	assign _0968_ = (_1342_ ? \mchip.internal [112] : _0967_);
	assign _0969_ = _0397_ | _1518_;
	assign _0970_ = _1367_ & ~_0969_;
	assign _0971_ = _0400_ | _1518_;
	assign _0972_ = _1367_ & ~_0971_;
	assign _0973_ = _0968_ & ~_0972_;
	assign _0974_ = _0973_ | _0970_;
	assign _0020_ = (_1547_ ? _0968_ : _0974_);
	assign _0975_ = \mchip.key [113] ^ \mchip.plaintext [113];
	assign _0976_ = (_1342_ ? \mchip.internal [113] : _0975_);
	assign _0977_ = _0407_ | _1518_;
	assign _0978_ = _1367_ & ~_0977_;
	assign _0979_ = _0410_ | _1518_;
	assign _0980_ = _1367_ & ~_0979_;
	assign _0981_ = _0976_ & ~_0980_;
	assign _0982_ = _0981_ | _0978_;
	assign _0021_ = (_1547_ ? _0976_ : _0982_);
	assign _0983_ = \mchip.key [114] ^ \mchip.plaintext [114];
	assign _0984_ = (_1342_ ? \mchip.internal [114] : _0983_);
	assign _0985_ = _0417_ | _1518_;
	assign _0986_ = _1367_ & ~_0985_;
	assign _0987_ = _0420_ | _1518_;
	assign _0988_ = _1367_ & ~_0987_;
	assign _0989_ = _0984_ & ~_0988_;
	assign _0990_ = _0989_ | _0986_;
	assign _0022_ = (_1547_ ? _0984_ : _0990_);
	assign _0991_ = \mchip.key [115] ^ \mchip.plaintext [115];
	assign _0992_ = (_1342_ ? \mchip.internal [115] : _0991_);
	assign _0993_ = _0427_ | _1518_;
	assign _0994_ = _1367_ & ~_0993_;
	assign _0995_ = _0430_ | _1518_;
	assign _0996_ = _1367_ & ~_0995_;
	assign _0997_ = _0992_ & ~_0996_;
	assign _0998_ = _0997_ | _0994_;
	assign _0023_ = (_1547_ ? _0992_ : _0998_);
	assign _0999_ = \mchip.key [116] ^ \mchip.plaintext [116];
	assign _1000_ = (_1342_ ? \mchip.internal [116] : _0999_);
	assign _1001_ = _0437_ | _1518_;
	assign _1002_ = _1367_ & ~_1001_;
	assign _1003_ = _0440_ | _1518_;
	assign _1004_ = _1367_ & ~_1003_;
	assign _1005_ = _1000_ & ~_1004_;
	assign _1006_ = _1005_ | _1002_;
	assign _0024_ = (_1547_ ? _1000_ : _1006_);
	assign _1007_ = \mchip.key [117] ^ \mchip.plaintext [117];
	assign _1008_ = (_1342_ ? \mchip.internal [117] : _1007_);
	assign _1009_ = _0447_ | _1518_;
	assign _1010_ = _1367_ & ~_1009_;
	assign _1011_ = _0450_ | _1518_;
	assign _1012_ = _1367_ & ~_1011_;
	assign _1013_ = _1008_ & ~_1012_;
	assign _1014_ = _1013_ | _1010_;
	assign _0025_ = (_1547_ ? _1008_ : _1014_);
	assign _1015_ = \mchip.key [118] ^ \mchip.plaintext [118];
	assign _1016_ = (_1342_ ? \mchip.internal [118] : _1015_);
	assign _1017_ = _0457_ | _1518_;
	assign _1018_ = _1367_ & ~_1017_;
	assign _1019_ = _0460_ | _1518_;
	assign _1020_ = _1367_ & ~_1019_;
	assign _1021_ = _1016_ & ~_1020_;
	assign _1022_ = _1021_ | _1018_;
	assign _0026_ = (_1547_ ? _1016_ : _1022_);
	assign _1023_ = \mchip.key [119] ^ \mchip.plaintext [119];
	assign _1024_ = (_1342_ ? \mchip.internal [119] : _1023_);
	assign _1025_ = _0467_ | _1518_;
	assign _1026_ = _1367_ & ~_1025_;
	assign _1027_ = _0470_ | _1518_;
	assign _1028_ = _1367_ & ~_1027_;
	assign _1029_ = _1024_ & ~_1028_;
	assign _1030_ = _1029_ | _1026_;
	assign _0027_ = (_1547_ ? _1024_ : _1030_);
	assign _1031_ = \mchip.key [120] ^ \mchip.plaintext [120];
	assign _1032_ = (_1342_ ? \mchip.internal [120] : _1031_);
	assign _1033_ = _0477_ | _1518_;
	assign _1034_ = _1367_ & ~_1033_;
	assign _1035_ = _0480_ | _1518_;
	assign _1036_ = _1367_ & ~_1035_;
	assign _1037_ = _1032_ & ~_1036_;
	assign _1038_ = _1037_ | _1034_;
	assign _0029_ = (_1547_ ? _1032_ : _1038_);
	assign _1039_ = \mchip.key [121] ^ \mchip.plaintext [121];
	assign _1040_ = (_1342_ ? \mchip.internal [121] : _1039_);
	assign _1041_ = _0487_ | _1518_;
	assign _1042_ = _1367_ & ~_1041_;
	assign _1043_ = _0490_ | _1518_;
	assign _1044_ = _1367_ & ~_1043_;
	assign _1045_ = _1040_ & ~_1044_;
	assign _1046_ = _1045_ | _1042_;
	assign _0030_ = (_1547_ ? _1040_ : _1046_);
	assign _1047_ = \mchip.key [122] ^ \mchip.plaintext [122];
	assign _1048_ = (_1342_ ? \mchip.internal [122] : _1047_);
	assign _1049_ = _0497_ | _1518_;
	assign _1050_ = _1367_ & ~_1049_;
	assign _1051_ = _0500_ | _1518_;
	assign _1052_ = _1367_ & ~_1051_;
	assign _1053_ = _1048_ & ~_1052_;
	assign _1054_ = _1053_ | _1050_;
	assign _0031_ = (_1547_ ? _1048_ : _1054_);
	assign _1055_ = \mchip.key [123] ^ \mchip.plaintext [123];
	assign _1056_ = (_1342_ ? \mchip.internal [123] : _1055_);
	assign _1057_ = _0507_ | _1518_;
	assign _1058_ = _1367_ & ~_1057_;
	assign _1059_ = _0510_ | _1518_;
	assign _1060_ = _1367_ & ~_1059_;
	assign _1061_ = _1056_ & ~_1060_;
	assign _1062_ = _1061_ | _1058_;
	assign _0032_ = (_1547_ ? _1056_ : _1062_);
	assign _1063_ = \mchip.key [124] ^ \mchip.plaintext [124];
	assign _1064_ = (_1342_ ? \mchip.internal [124] : _1063_);
	assign _1065_ = _0517_ | _1518_;
	assign _1066_ = _1367_ & ~_1065_;
	assign _1067_ = _0520_ | _1518_;
	assign _1068_ = _1367_ & ~_1067_;
	assign _1069_ = _1064_ & ~_1068_;
	assign _1070_ = _1069_ | _1066_;
	assign _0033_ = (_1547_ ? _1064_ : _1070_);
	assign _1071_ = \mchip.key [125] ^ \mchip.plaintext [125];
	assign _1072_ = (_1342_ ? \mchip.internal [125] : _1071_);
	assign _1073_ = _0527_ | _1518_;
	assign _1074_ = _1367_ & ~_1073_;
	assign _1075_ = _0530_ | _1518_;
	assign _1076_ = _1367_ & ~_1075_;
	assign _1077_ = _1072_ & ~_1076_;
	assign _1078_ = _1077_ | _1074_;
	assign _0034_ = (_1547_ ? _1072_ : _1078_);
	assign _1079_ = \mchip.key [126] ^ \mchip.plaintext [126];
	assign _1080_ = (_1342_ ? \mchip.internal [126] : _1079_);
	assign _1081_ = _0537_ | _1518_;
	assign _1082_ = _1367_ & ~_1081_;
	assign _1083_ = _0540_ | _1518_;
	assign _1084_ = _1367_ & ~_1083_;
	assign _1085_ = _1080_ & ~_1084_;
	assign _1086_ = _1085_ | _1082_;
	assign _0035_ = (_1547_ ? _1080_ : _1086_);
	assign _1087_ = \mchip.key [127] ^ \mchip.plaintext [127];
	assign _1088_ = (_1342_ ? \mchip.internal [127] : _1087_);
	assign _1089_ = _0547_ | _1518_;
	assign _1090_ = _1367_ & ~_1089_;
	assign _1091_ = _0550_ | _1518_;
	assign _1092_ = _1367_ & ~_1091_;
	assign _1093_ = _1088_ & ~_1092_;
	assign _1094_ = _1093_ | _1090_;
	assign _0036_ = (_1547_ ? _1088_ : _1094_);
	assign _1095_ = _1306_ & _1304_;
	assign _1096_ = _1095_ & ~\mchip.state [6];
	assign _1097_ = (\mchip.state [1] ? _1368_ : _1369_);
	assign _1098_ = (\mchip.state [1] ? _1371_ : _1372_);
	assign _1099_ = (\mchip.state [2] ? _1098_ : _1097_);
	assign _1100_ = ~(_1340_ | _1322_);
	assign _1101_ = (\mchip.state [1] ? _1375_ : _1376_);
	assign _1102_ = (\mchip.state [1] ? _1378_ : _1379_);
	assign _1103_ = (\mchip.state [2] ? _1102_ : _1101_);
	assign _1104_ = (_1100_ ? _1099_ : _1103_);
	assign _1105_ = _1306_ ^ \mchip.state [4];
	assign _1106_ = (\mchip.state [1] ? _1383_ : _1384_);
	assign _1107_ = (\mchip.state [1] ? _1386_ : _1387_);
	assign _1108_ = (\mchip.state [2] ? _1107_ : _1106_);
	assign _1109_ = (\mchip.state [1] ? _1390_ : _1391_);
	assign _1110_ = (\mchip.state [1] ? _1393_ : _1394_);
	assign _1111_ = (\mchip.state [2] ? _1110_ : _1109_);
	assign _1112_ = (_1100_ ? _1108_ : _1111_);
	assign _1113_ = (_1105_ ? _1104_ : _1112_);
	assign _1114_ = _1306_ & ~\mchip.state [4];
	assign _1115_ = _1114_ ^ \mchip.state [5];
	assign _1116_ = (\mchip.state [1] ? _1399_ : _1400_);
	assign _1117_ = (\mchip.state [1] ? _1402_ : _1403_);
	assign _1118_ = (\mchip.state [2] ? _1117_ : _1116_);
	assign _1119_ = (\mchip.state [1] ? _1406_ : _1407_);
	assign _1120_ = (\mchip.state [1] ? _1409_ : _1410_);
	assign _1121_ = (\mchip.state [2] ? _1120_ : _1119_);
	assign _1122_ = (_1100_ ? _1118_ : _1121_);
	assign _1123_ = (\mchip.state [1] ? _1414_ : _1415_);
	assign _1124_ = (\mchip.state [1] ? _1417_ : _1418_);
	assign _1125_ = (\mchip.state [2] ? _1124_ : _1123_);
	assign _1126_ = (\mchip.state [1] ? _1421_ : _1422_);
	assign _1127_ = (\mchip.state [1] ? _1424_ : _1425_);
	assign _1128_ = (\mchip.state [2] ? _1127_ : _1126_);
	assign _1129_ = (_1100_ ? _1125_ : _1128_);
	assign _1130_ = (_1105_ ? _1122_ : _1129_);
	assign _1131_ = (_1115_ ? _1113_ : _1130_);
	assign _1132_ = _1095_ ^ \mchip.state [6];
	assign _1133_ = (\mchip.state [1] ? _1431_ : _1432_);
	assign _1134_ = (\mchip.state [1] ? _1434_ : _1435_);
	assign _1135_ = (\mchip.state [2] ? _1134_ : _1133_);
	assign _1136_ = (\mchip.state [1] ? _1438_ : _1439_);
	assign _1137_ = (\mchip.state [1] ? _1441_ : _1442_);
	assign _1138_ = (\mchip.state [2] ? _1137_ : _1136_);
	assign _1139_ = (_1100_ ? _1135_ : _1138_);
	assign _1140_ = (\mchip.state [1] ? _1446_ : _1447_);
	assign _1141_ = (\mchip.state [1] ? _1449_ : _1450_);
	assign _1142_ = (\mchip.state [2] ? _1141_ : _1140_);
	assign _1143_ = (\mchip.state [1] ? _1453_ : _1454_);
	assign _1144_ = (\mchip.state [1] ? _1456_ : _1457_);
	assign _1145_ = (\mchip.state [2] ? _1144_ : _1143_);
	assign _1146_ = (_1100_ ? _1142_ : _1145_);
	assign _1147_ = (_1105_ ? _1139_ : _1146_);
	assign _1148_ = (\mchip.state [1] ? _1462_ : _1463_);
	assign _1149_ = (\mchip.state [1] ? _1465_ : _1466_);
	assign _1150_ = (\mchip.state [2] ? _1149_ : _1148_);
	assign _1151_ = (\mchip.state [1] ? _1469_ : _1470_);
	assign _1152_ = (\mchip.state [1] ? _1472_ : _1473_);
	assign _1153_ = (\mchip.state [2] ? _1152_ : _1151_);
	assign _1154_ = (_1100_ ? _1150_ : _1153_);
	assign _1155_ = (\mchip.state [1] ? _1477_ : _1478_);
	assign _1156_ = (\mchip.state [1] ? _1480_ : _1481_);
	assign _1157_ = (\mchip.state [2] ? _1156_ : _1155_);
	assign _1158_ = (\mchip.state [1] ? _1484_ : _1485_);
	assign _1159_ = (\mchip.state [1] ? _1487_ : _1488_);
	assign _1160_ = (\mchip.state [2] ? _1159_ : _1158_);
	assign _1161_ = (_1100_ ? _1157_ : _1160_);
	assign _1162_ = (_1105_ ? _1154_ : _1161_);
	assign _1163_ = (_1115_ ? _1147_ : _1162_);
	assign _1164_ = (_1132_ ? _1131_ : _1163_);
	assign _1740_ = _1164_ & ~_1096_;
	assign _1165_ = _1503_ | _1317_;
	assign _0003_ = _1316_ & ~_1165_;
	assign _1166_ = _1307_ & _1306_;
	assign _1167_ = _1166_ ^ _1352_;
	assign _1168_ = _1167_ | _1317_;
	assign _0004_ = _1316_ & ~_1168_;
	assign _1169_ = _1166_ & ~\mchip.state [4];
	assign _1170_ = _1169_ ^ _1355_;
	assign _1171_ = _1170_ | _1317_;
	assign _0005_ = _1316_ & ~_1171_;
	assign _0138_ = _1309_ & ~_1317_;
	assign _1172_ = _1307_ ^ \mchip.state [2];
	assign _0139_ = _1172_ & ~_1317_;
	assign _1173_ = _1307_ & ~\mchip.state [2];
	assign _1174_ = _1173_ ^ \mchip.state [3];
	assign _0140_ = _1174_ & ~_1317_;
	assign _1175_ = _1166_ & ~_1320_;
	assign _1176_ = _1175_ ^ _1329_;
	assign _0141_ = _1318_ & ~_1176_;
	assign _1177_ = \mchip.key [0] ^ \mchip.plaintext [0];
	assign _1178_ = (_1342_ ? \mchip.internal [0] : _1177_);
	assign _1179_ = ~_1367_;
	assign _1180_ = _1499_ | _1495_;
	assign _1181_ = _1180_ | \mchip.state [0];
	assign _1182_ = _1181_ | _1502_;
	assign _1183_ = _1182_ | _1506_;
	assign _1184_ = _1183_ | _1509_;
	assign _1185_ = _1184_ | _1511_;
	assign _1186_ = _1185_ | _1515_;
	assign _1187_ = _1186_ | _1518_;
	assign _1188_ = _1179_ & ~_1187_;
	assign _1189_ = _1366_ | ~_1498_;
	assign _1190_ = _1189_ | \mchip.state [0];
	assign _1191_ = _1190_ | _1502_;
	assign _1192_ = _1191_ | _1506_;
	assign _1193_ = _1192_ | _1509_;
	assign _1194_ = _1193_ | _1511_;
	assign _1195_ = _1194_ | _1515_;
	assign _1196_ = _1195_ | _1518_;
	assign _1197_ = _1179_ & ~_1196_;
	assign _1198_ = _1178_ & ~_1197_;
	assign _1199_ = _1198_ | _1188_;
	assign _0006_ = (_1547_ ? _1178_ : _1199_);
	assign _1200_ = \mchip.key [1] ^ \mchip.plaintext [1];
	assign _1201_ = (_1342_ ? \mchip.internal [1] : _1200_);
	assign _1202_ = _0567_ | _1519_;
	assign _1203_ = _1367_ & ~_1202_;
	assign _1204_ = _0570_ | _1519_;
	assign _1205_ = _1367_ & ~_1204_;
	assign _1206_ = _1201_ & ~_1205_;
	assign _1207_ = _1206_ | _1203_;
	assign _0045_ = (_1547_ ? _1201_ : _1207_);
	assign _1208_ = \mchip.key [2] ^ \mchip.plaintext [2];
	assign _1209_ = (_1342_ ? \mchip.internal [2] : _1208_);
	assign _1210_ = _0577_ | _1519_;
	assign _1211_ = _1367_ & ~_1210_;
	assign _1212_ = _0580_ | _1519_;
	assign _1213_ = _1367_ & ~_1212_;
	assign _1214_ = _1209_ & ~_1213_;
	assign _1215_ = _1214_ | _1211_;
	assign _0056_ = (_1547_ ? _1209_ : _1215_);
	assign _1216_ = \mchip.key [3] ^ \mchip.plaintext [3];
	assign _1217_ = (_1342_ ? \mchip.internal [3] : _1216_);
	assign _1218_ = _0587_ | _1519_;
	assign _1219_ = _1367_ & ~_1218_;
	assign _1220_ = _0590_ | _1519_;
	assign _1221_ = _1367_ & ~_1220_;
	assign _1222_ = _1217_ & ~_1221_;
	assign _1223_ = _1222_ | _1219_;
	assign _0067_ = (_1547_ ? _1217_ : _1223_);
	assign _1224_ = \mchip.key [4] ^ \mchip.plaintext [4];
	assign _1225_ = (_1342_ ? \mchip.internal [4] : _1224_);
	assign _1226_ = _0597_ | _1519_;
	assign _1227_ = _1367_ & ~_1226_;
	assign _1228_ = _0600_ | _1519_;
	assign _1229_ = _1367_ & ~_1228_;
	assign _1230_ = _1225_ & ~_1229_;
	assign _1231_ = _1230_ | _1227_;
	assign _0078_ = (_1547_ ? _1225_ : _1231_);
	assign _1232_ = \mchip.key [5] ^ \mchip.plaintext [5];
	assign _1233_ = (_1342_ ? \mchip.internal [5] : _1232_);
	assign _1234_ = _0607_ | _1519_;
	assign _1235_ = _1367_ & ~_1234_;
	assign _1236_ = _0610_ | _1519_;
	assign _1237_ = _1367_ & ~_1236_;
	assign _1238_ = _1233_ & ~_1237_;
	assign _1239_ = _1238_ | _1235_;
	assign _0089_ = (_1547_ ? _1233_ : _1239_);
	assign _1240_ = \mchip.key [6] ^ \mchip.plaintext [6];
	assign _1241_ = (_1342_ ? \mchip.internal [6] : _1240_);
	assign _1242_ = _0617_ | _1519_;
	assign _1243_ = _1367_ & ~_1242_;
	assign _1244_ = _0620_ | _1519_;
	assign _1245_ = _1367_ & ~_1244_;
	assign _1246_ = _1241_ & ~_1245_;
	assign _1247_ = _1246_ | _1243_;
	assign _0100_ = (_1547_ ? _1241_ : _1247_);
	assign _1248_ = \mchip.key [7] ^ \mchip.plaintext [7];
	assign _1249_ = (_1342_ ? \mchip.internal [7] : _1248_);
	assign _1250_ = _0627_ | _1519_;
	assign _1251_ = _1367_ & ~_1250_;
	assign _1252_ = _0630_ | _1519_;
	assign _1253_ = _1367_ & ~_1252_;
	assign _1254_ = _1249_ & ~_1253_;
	assign _1255_ = _1254_ | _1251_;
	assign _0111_ = (_1547_ ? _1249_ : _1255_);
	assign _1256_ = \mchip.key [8] ^ \mchip.plaintext [8];
	assign _1257_ = (_1342_ ? \mchip.internal [8] : _1256_);
	assign _1258_ = _0637_ | _1519_;
	assign _1259_ = _1367_ & ~_1258_;
	assign _1260_ = _0640_ | _1519_;
	assign _1261_ = _1367_ & ~_1260_;
	assign _1262_ = _1257_ & ~_1261_;
	assign _1263_ = _1262_ | _1259_;
	assign _0122_ = (_1547_ ? _1257_ : _1263_);
	assign _1264_ = \mchip.key [9] ^ \mchip.plaintext [9];
	assign _1265_ = (_1342_ ? \mchip.internal [9] : _1264_);
	assign _1266_ = _0647_ | _1519_;
	assign _1267_ = _1367_ & ~_1266_;
	assign _1268_ = _0650_ | _1519_;
	assign _1269_ = _1367_ & ~_1268_;
	assign _1270_ = _1265_ & ~_1269_;
	assign _1271_ = _1270_ | _1267_;
	assign _0133_ = (_1547_ ? _1265_ : _1271_);
	assign _1272_ = \mchip.key [10] ^ \mchip.plaintext [10];
	assign _1273_ = (_1342_ ? \mchip.internal [10] : _1272_);
	assign _1274_ = _0657_ | _1519_;
	assign _1275_ = _1367_ & ~_1274_;
	assign _1276_ = _0660_ | _1519_;
	assign _1277_ = _1367_ & ~_1276_;
	assign _1278_ = _1273_ & ~_1277_;
	assign _1279_ = _1278_ | _1275_;
	assign _0017_ = (_1547_ ? _1273_ : _1279_);
	assign _1280_ = \mchip.key [11] ^ \mchip.plaintext [11];
	assign _1281_ = (_1342_ ? \mchip.internal [11] : _1280_);
	assign _1282_ = _0667_ | _1519_;
	assign _1283_ = _1367_ & ~_1282_;
	assign _1284_ = _0670_ | _1519_;
	assign _1285_ = _1367_ & ~_1284_;
	assign _1286_ = _1281_ & ~_1285_;
	assign _1287_ = _1286_ | _1283_;
	assign _0028_ = (_1547_ ? _1281_ : _1287_);
	assign _1288_ = \mchip.key [12] ^ \mchip.plaintext [12];
	assign _1289_ = (_1342_ ? \mchip.internal [12] : _1288_);
	assign _1290_ = _0677_ | _1519_;
	assign _1291_ = _1367_ & ~_1290_;
	assign _1292_ = _0680_ | _1519_;
	assign _1293_ = _1367_ & ~_1292_;
	assign _1294_ = _1289_ & ~_1293_;
	assign _1295_ = _1294_ | _1291_;
	assign _0037_ = (_1547_ ? _1289_ : _1295_);
	assign _1296_ = \mchip.key [13] ^ \mchip.plaintext [13];
	assign _1297_ = (_1342_ ? \mchip.internal [13] : _1296_);
	assign _1298_ = _0687_ | _1519_;
	assign _1299_ = _1367_ & ~_1298_;
	assign _1300_ = _0690_ | _1519_;
	assign _1301_ = _1367_ & ~_1300_;
	assign _1302_ = _1297_ & ~_1301_;
	assign _1303_ = _1302_ | _1299_;
	assign _0038_ = (_1547_ ? _1297_ : _1303_);
	always @(posedge io_in[12]) \mchip.plaintext_in_last  <= io_in[9];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [0] <= io_in[0];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [1] <= io_in[1];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [2] <= io_in[2];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [3] <= io_in[3];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [4] <= io_in[4];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [5] <= io_in[5];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [6] <= io_in[6];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [7] <= io_in[7];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [8] <= \mchip.plaintext [0];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [9] <= \mchip.plaintext [1];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [10] <= \mchip.plaintext [2];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [11] <= \mchip.plaintext [3];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [12] <= \mchip.plaintext [4];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [13] <= \mchip.plaintext [5];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [14] <= \mchip.plaintext [6];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [15] <= \mchip.plaintext [7];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [16] <= \mchip.plaintext [8];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [17] <= \mchip.plaintext [9];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [18] <= \mchip.plaintext [10];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [19] <= \mchip.plaintext [11];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [20] <= \mchip.plaintext [12];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [21] <= \mchip.plaintext [13];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [22] <= \mchip.plaintext [14];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [23] <= \mchip.plaintext [15];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [24] <= \mchip.plaintext [16];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [25] <= \mchip.plaintext [17];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [26] <= \mchip.plaintext [18];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [27] <= \mchip.plaintext [19];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [28] <= \mchip.plaintext [20];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [29] <= \mchip.plaintext [21];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [30] <= \mchip.plaintext [22];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [31] <= \mchip.plaintext [23];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [32] <= \mchip.plaintext [24];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [33] <= \mchip.plaintext [25];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [34] <= \mchip.plaintext [26];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [35] <= \mchip.plaintext [27];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [36] <= \mchip.plaintext [28];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [37] <= \mchip.plaintext [29];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [38] <= \mchip.plaintext [30];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [39] <= \mchip.plaintext [31];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [40] <= \mchip.plaintext [32];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [41] <= \mchip.plaintext [33];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [42] <= \mchip.plaintext [34];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [43] <= \mchip.plaintext [35];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [44] <= \mchip.plaintext [36];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [45] <= \mchip.plaintext [37];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [46] <= \mchip.plaintext [38];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [47] <= \mchip.plaintext [39];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [48] <= \mchip.plaintext [40];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [49] <= \mchip.plaintext [41];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [50] <= \mchip.plaintext [42];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [51] <= \mchip.plaintext [43];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [52] <= \mchip.plaintext [44];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [53] <= \mchip.plaintext [45];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [54] <= \mchip.plaintext [46];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [55] <= \mchip.plaintext [47];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [56] <= \mchip.plaintext [48];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [57] <= \mchip.plaintext [49];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [58] <= \mchip.plaintext [50];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [59] <= \mchip.plaintext [51];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [60] <= \mchip.plaintext [52];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [61] <= \mchip.plaintext [53];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [62] <= \mchip.plaintext [54];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [63] <= \mchip.plaintext [55];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [64] <= \mchip.plaintext [56];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [65] <= \mchip.plaintext [57];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [66] <= \mchip.plaintext [58];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [67] <= \mchip.plaintext [59];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [68] <= \mchip.plaintext [60];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [69] <= \mchip.plaintext [61];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [70] <= \mchip.plaintext [62];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [71] <= \mchip.plaintext [63];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [72] <= \mchip.plaintext [64];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [73] <= \mchip.plaintext [65];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [74] <= \mchip.plaintext [66];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [75] <= \mchip.plaintext [67];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [76] <= \mchip.plaintext [68];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [77] <= \mchip.plaintext [69];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [78] <= \mchip.plaintext [70];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [79] <= \mchip.plaintext [71];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [80] <= \mchip.plaintext [72];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [81] <= \mchip.plaintext [73];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [82] <= \mchip.plaintext [74];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [83] <= \mchip.plaintext [75];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [84] <= \mchip.plaintext [76];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [85] <= \mchip.plaintext [77];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [86] <= \mchip.plaintext [78];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [87] <= \mchip.plaintext [79];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [88] <= \mchip.plaintext [80];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [89] <= \mchip.plaintext [81];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [90] <= \mchip.plaintext [82];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [91] <= \mchip.plaintext [83];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [92] <= \mchip.plaintext [84];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [93] <= \mchip.plaintext [85];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [94] <= \mchip.plaintext [86];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [95] <= \mchip.plaintext [87];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [96] <= \mchip.plaintext [88];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [97] <= \mchip.plaintext [89];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [98] <= \mchip.plaintext [90];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [99] <= \mchip.plaintext [91];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [100] <= \mchip.plaintext [92];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [101] <= \mchip.plaintext [93];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [102] <= \mchip.plaintext [94];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [103] <= \mchip.plaintext [95];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [104] <= \mchip.plaintext [96];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [105] <= \mchip.plaintext [97];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [106] <= \mchip.plaintext [98];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [107] <= \mchip.plaintext [99];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [108] <= \mchip.plaintext [100];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [109] <= \mchip.plaintext [101];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [110] <= \mchip.plaintext [102];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [111] <= \mchip.plaintext [103];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [112] <= \mchip.plaintext [104];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [113] <= \mchip.plaintext [105];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [114] <= \mchip.plaintext [106];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [115] <= \mchip.plaintext [107];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [116] <= \mchip.plaintext [108];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [117] <= \mchip.plaintext [109];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [118] <= \mchip.plaintext [110];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [119] <= \mchip.plaintext [111];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [120] <= \mchip.plaintext [112];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [121] <= \mchip.plaintext [113];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [122] <= \mchip.plaintext [114];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [123] <= \mchip.plaintext [115];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [124] <= \mchip.plaintext [116];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [125] <= \mchip.plaintext [117];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [126] <= \mchip.plaintext [118];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.plaintext [127] <= \mchip.plaintext [119];
	always @(posedge io_in[12])
		if (_0136_)
			\mchip.state [1] <= 1'h1;
		else if (_0001_)
			\mchip.state [1] <= _0003_;
	always @(posedge io_in[12])
		if (_0136_)
			\mchip.state [4] <= 1'h1;
		else if (_0001_)
			\mchip.state [4] <= _0004_;
	always @(posedge io_in[12])
		if (_0136_)
			\mchip.state [5] <= 1'h1;
		else if (_0001_)
			\mchip.state [5] <= _0005_;
	always @(posedge io_in[12]) \mchip.key_in_last  <= io_in[8];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [0] <= io_in[0];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [1] <= io_in[1];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [2] <= io_in[2];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [3] <= io_in[3];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [4] <= io_in[4];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [5] <= io_in[5];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [6] <= io_in[6];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [7] <= io_in[7];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [8] <= \mchip.key [0];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [9] <= \mchip.key [1];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [10] <= \mchip.key [2];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [11] <= \mchip.key [3];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [12] <= \mchip.key [4];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [13] <= \mchip.key [5];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [14] <= \mchip.key [6];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [15] <= \mchip.key [7];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [16] <= \mchip.key [8];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [17] <= \mchip.key [9];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [18] <= \mchip.key [10];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [19] <= \mchip.key [11];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [20] <= \mchip.key [12];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [21] <= \mchip.key [13];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [22] <= \mchip.key [14];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [23] <= \mchip.key [15];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [24] <= \mchip.key [16];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [25] <= \mchip.key [17];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [26] <= \mchip.key [18];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [27] <= \mchip.key [19];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [28] <= \mchip.key [20];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [29] <= \mchip.key [21];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [30] <= \mchip.key [22];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [31] <= \mchip.key [23];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [32] <= \mchip.key [24];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [33] <= \mchip.key [25];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [34] <= \mchip.key [26];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [35] <= \mchip.key [27];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [36] <= \mchip.key [28];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [37] <= \mchip.key [29];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [38] <= \mchip.key [30];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [39] <= \mchip.key [31];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [40] <= \mchip.key [32];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [41] <= \mchip.key [33];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [42] <= \mchip.key [34];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [43] <= \mchip.key [35];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [44] <= \mchip.key [36];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [45] <= \mchip.key [37];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [46] <= \mchip.key [38];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [47] <= \mchip.key [39];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [48] <= \mchip.key [40];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [49] <= \mchip.key [41];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [50] <= \mchip.key [42];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [51] <= \mchip.key [43];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [52] <= \mchip.key [44];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [53] <= \mchip.key [45];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [54] <= \mchip.key [46];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [55] <= \mchip.key [47];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [56] <= \mchip.key [48];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [57] <= \mchip.key [49];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [58] <= \mchip.key [50];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [59] <= \mchip.key [51];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [60] <= \mchip.key [52];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [61] <= \mchip.key [53];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [62] <= \mchip.key [54];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [63] <= \mchip.key [55];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [64] <= \mchip.key [56];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [65] <= \mchip.key [57];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [66] <= \mchip.key [58];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [67] <= \mchip.key [59];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [68] <= \mchip.key [60];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [69] <= \mchip.key [61];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [70] <= \mchip.key [62];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [71] <= \mchip.key [63];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [72] <= \mchip.key [64];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [73] <= \mchip.key [65];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [74] <= \mchip.key [66];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [75] <= \mchip.key [67];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [76] <= \mchip.key [68];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [77] <= \mchip.key [69];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [78] <= \mchip.key [70];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [79] <= \mchip.key [71];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [80] <= \mchip.key [72];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [81] <= \mchip.key [73];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [82] <= \mchip.key [74];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [83] <= \mchip.key [75];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [84] <= \mchip.key [76];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [85] <= \mchip.key [77];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [86] <= \mchip.key [78];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [87] <= \mchip.key [79];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [88] <= \mchip.key [80];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [89] <= \mchip.key [81];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [90] <= \mchip.key [82];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [91] <= \mchip.key [83];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [92] <= \mchip.key [84];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [93] <= \mchip.key [85];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [94] <= \mchip.key [86];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [95] <= \mchip.key [87];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [96] <= \mchip.key [88];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [97] <= \mchip.key [89];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [98] <= \mchip.key [90];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [99] <= \mchip.key [91];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [100] <= \mchip.key [92];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [101] <= \mchip.key [93];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [102] <= \mchip.key [94];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [103] <= \mchip.key [95];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [104] <= \mchip.key [96];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [105] <= \mchip.key [97];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [106] <= \mchip.key [98];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [107] <= \mchip.key [99];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [108] <= \mchip.key [100];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [109] <= \mchip.key [101];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [110] <= \mchip.key [102];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [111] <= \mchip.key [103];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [112] <= \mchip.key [104];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [113] <= \mchip.key [105];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [114] <= \mchip.key [106];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [115] <= \mchip.key [107];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [116] <= \mchip.key [108];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [117] <= \mchip.key [109];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [118] <= \mchip.key [110];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [119] <= \mchip.key [111];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [120] <= \mchip.key [112];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [121] <= \mchip.key [113];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [122] <= \mchip.key [114];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [123] <= \mchip.key [115];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [124] <= \mchip.key [116];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [125] <= \mchip.key [117];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [126] <= \mchip.key [118];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.key [127] <= \mchip.key [119];
	always @(posedge io_in[12]) \mchip.internal [0] <= _0006_;
	always @(posedge io_in[12]) \mchip.internal [1] <= _0045_;
	always @(posedge io_in[12]) \mchip.internal [2] <= _0056_;
	always @(posedge io_in[12]) \mchip.internal [3] <= _0067_;
	always @(posedge io_in[12]) \mchip.internal [4] <= _0078_;
	always @(posedge io_in[12]) \mchip.internal [5] <= _0089_;
	always @(posedge io_in[12]) \mchip.internal [6] <= _0100_;
	always @(posedge io_in[12]) \mchip.internal [7] <= _0111_;
	always @(posedge io_in[12]) \mchip.internal [8] <= _0122_;
	always @(posedge io_in[12]) \mchip.internal [9] <= _0133_;
	always @(posedge io_in[12]) \mchip.internal [10] <= _0017_;
	always @(posedge io_in[12]) \mchip.internal [11] <= _0028_;
	always @(posedge io_in[12]) \mchip.internal [12] <= _0037_;
	always @(posedge io_in[12]) \mchip.internal [13] <= _0038_;
	always @(posedge io_in[12]) \mchip.internal [14] <= _0039_;
	always @(posedge io_in[12]) \mchip.internal [15] <= _0040_;
	always @(posedge io_in[12]) \mchip.internal [16] <= _0041_;
	always @(posedge io_in[12]) \mchip.internal [17] <= _0042_;
	always @(posedge io_in[12]) \mchip.internal [18] <= _0043_;
	always @(posedge io_in[12]) \mchip.internal [19] <= _0044_;
	always @(posedge io_in[12]) \mchip.internal [20] <= _0046_;
	always @(posedge io_in[12]) \mchip.internal [21] <= _0047_;
	always @(posedge io_in[12]) \mchip.internal [22] <= _0048_;
	always @(posedge io_in[12]) \mchip.internal [23] <= _0049_;
	always @(posedge io_in[12]) \mchip.internal [24] <= _0050_;
	always @(posedge io_in[12]) \mchip.internal [25] <= _0051_;
	always @(posedge io_in[12]) \mchip.internal [26] <= _0052_;
	always @(posedge io_in[12]) \mchip.internal [27] <= _0053_;
	always @(posedge io_in[12]) \mchip.internal [28] <= _0054_;
	always @(posedge io_in[12]) \mchip.internal [29] <= _0055_;
	always @(posedge io_in[12]) \mchip.internal [30] <= _0057_;
	always @(posedge io_in[12]) \mchip.internal [31] <= _0058_;
	always @(posedge io_in[12]) \mchip.internal [32] <= _0059_;
	always @(posedge io_in[12]) \mchip.internal [33] <= _0060_;
	always @(posedge io_in[12]) \mchip.internal [34] <= _0061_;
	always @(posedge io_in[12]) \mchip.internal [35] <= _0062_;
	always @(posedge io_in[12]) \mchip.internal [36] <= _0063_;
	always @(posedge io_in[12]) \mchip.internal [37] <= _0064_;
	always @(posedge io_in[12]) \mchip.internal [38] <= _0065_;
	always @(posedge io_in[12]) \mchip.internal [39] <= _0066_;
	always @(posedge io_in[12]) \mchip.internal [40] <= _0068_;
	always @(posedge io_in[12]) \mchip.internal [41] <= _0069_;
	always @(posedge io_in[12]) \mchip.internal [42] <= _0070_;
	always @(posedge io_in[12]) \mchip.internal [43] <= _0071_;
	always @(posedge io_in[12]) \mchip.internal [44] <= _0072_;
	always @(posedge io_in[12]) \mchip.internal [45] <= _0073_;
	always @(posedge io_in[12]) \mchip.internal [46] <= _0074_;
	always @(posedge io_in[12]) \mchip.internal [47] <= _0075_;
	always @(posedge io_in[12]) \mchip.internal [48] <= _0076_;
	always @(posedge io_in[12]) \mchip.internal [49] <= _0077_;
	always @(posedge io_in[12]) \mchip.internal [50] <= _0079_;
	always @(posedge io_in[12]) \mchip.internal [51] <= _0080_;
	always @(posedge io_in[12]) \mchip.internal [52] <= _0081_;
	always @(posedge io_in[12]) \mchip.internal [53] <= _0082_;
	always @(posedge io_in[12]) \mchip.internal [54] <= _0083_;
	always @(posedge io_in[12]) \mchip.internal [55] <= _0084_;
	always @(posedge io_in[12]) \mchip.internal [56] <= _0085_;
	always @(posedge io_in[12]) \mchip.internal [57] <= _0086_;
	always @(posedge io_in[12]) \mchip.internal [58] <= _0087_;
	always @(posedge io_in[12]) \mchip.internal [59] <= _0088_;
	always @(posedge io_in[12]) \mchip.internal [60] <= _0090_;
	always @(posedge io_in[12]) \mchip.internal [61] <= _0091_;
	always @(posedge io_in[12]) \mchip.internal [62] <= _0092_;
	always @(posedge io_in[12]) \mchip.internal [63] <= _0093_;
	always @(posedge io_in[12]) \mchip.internal [64] <= _0094_;
	always @(posedge io_in[12]) \mchip.internal [65] <= _0095_;
	always @(posedge io_in[12]) \mchip.internal [66] <= _0096_;
	always @(posedge io_in[12]) \mchip.internal [67] <= _0097_;
	always @(posedge io_in[12]) \mchip.internal [68] <= _0098_;
	always @(posedge io_in[12]) \mchip.internal [69] <= _0099_;
	always @(posedge io_in[12]) \mchip.internal [70] <= _0101_;
	always @(posedge io_in[12]) \mchip.internal [71] <= _0102_;
	always @(posedge io_in[12]) \mchip.internal [72] <= _0103_;
	always @(posedge io_in[12]) \mchip.internal [73] <= _0104_;
	always @(posedge io_in[12]) \mchip.internal [74] <= _0105_;
	always @(posedge io_in[12]) \mchip.internal [75] <= _0106_;
	always @(posedge io_in[12]) \mchip.internal [76] <= _0107_;
	always @(posedge io_in[12]) \mchip.internal [77] <= _0108_;
	always @(posedge io_in[12]) \mchip.internal [78] <= _0109_;
	always @(posedge io_in[12]) \mchip.internal [79] <= _0110_;
	always @(posedge io_in[12]) \mchip.internal [80] <= _0112_;
	always @(posedge io_in[12]) \mchip.internal [81] <= _0113_;
	always @(posedge io_in[12]) \mchip.internal [82] <= _0114_;
	always @(posedge io_in[12]) \mchip.internal [83] <= _0115_;
	always @(posedge io_in[12]) \mchip.internal [84] <= _0116_;
	always @(posedge io_in[12]) \mchip.internal [85] <= _0117_;
	always @(posedge io_in[12]) \mchip.internal [86] <= _0118_;
	always @(posedge io_in[12]) \mchip.internal [87] <= _0119_;
	always @(posedge io_in[12]) \mchip.internal [88] <= _0120_;
	always @(posedge io_in[12]) \mchip.internal [89] <= _0121_;
	always @(posedge io_in[12]) \mchip.internal [90] <= _0123_;
	always @(posedge io_in[12]) \mchip.internal [91] <= _0124_;
	always @(posedge io_in[12]) \mchip.internal [92] <= _0125_;
	always @(posedge io_in[12]) \mchip.internal [93] <= _0126_;
	always @(posedge io_in[12]) \mchip.internal [94] <= _0127_;
	always @(posedge io_in[12]) \mchip.internal [95] <= _0128_;
	always @(posedge io_in[12]) \mchip.internal [96] <= _0129_;
	always @(posedge io_in[12]) \mchip.internal [97] <= _0130_;
	always @(posedge io_in[12]) \mchip.internal [98] <= _0131_;
	always @(posedge io_in[12]) \mchip.internal [99] <= _0132_;
	always @(posedge io_in[12]) \mchip.internal [100] <= _0007_;
	always @(posedge io_in[12]) \mchip.internal [101] <= _0008_;
	always @(posedge io_in[12]) \mchip.internal [102] <= _0009_;
	always @(posedge io_in[12]) \mchip.internal [103] <= _0010_;
	always @(posedge io_in[12]) \mchip.internal [104] <= _0011_;
	always @(posedge io_in[12]) \mchip.internal [105] <= _0012_;
	always @(posedge io_in[12]) \mchip.internal [106] <= _0013_;
	always @(posedge io_in[12]) \mchip.internal [107] <= _0014_;
	always @(posedge io_in[12]) \mchip.internal [108] <= _0015_;
	always @(posedge io_in[12]) \mchip.internal [109] <= _0016_;
	always @(posedge io_in[12]) \mchip.internal [110] <= _0018_;
	always @(posedge io_in[12]) \mchip.internal [111] <= _0019_;
	always @(posedge io_in[12]) \mchip.internal [112] <= _0020_;
	always @(posedge io_in[12]) \mchip.internal [113] <= _0021_;
	always @(posedge io_in[12]) \mchip.internal [114] <= _0022_;
	always @(posedge io_in[12]) \mchip.internal [115] <= _0023_;
	always @(posedge io_in[12]) \mchip.internal [116] <= _0024_;
	always @(posedge io_in[12]) \mchip.internal [117] <= _0025_;
	always @(posedge io_in[12]) \mchip.internal [118] <= _0026_;
	always @(posedge io_in[12]) \mchip.internal [119] <= _0027_;
	always @(posedge io_in[12]) \mchip.internal [120] <= _0029_;
	always @(posedge io_in[12]) \mchip.internal [121] <= _0030_;
	always @(posedge io_in[12]) \mchip.internal [122] <= _0031_;
	always @(posedge io_in[12]) \mchip.internal [123] <= _0032_;
	always @(posedge io_in[12]) \mchip.internal [124] <= _0033_;
	always @(posedge io_in[12]) \mchip.internal [125] <= _0034_;
	always @(posedge io_in[12]) \mchip.internal [126] <= _0035_;
	always @(posedge io_in[12]) \mchip.internal [127] <= _0036_;
	always @(posedge io_in[12])
		if (_0002_)
			\mchip.state [0] <= 1'h0;
		else if (_0000_)
			\mchip.state [0] <= _0138_;
	always @(posedge io_in[12])
		if (_0002_)
			\mchip.state [2] <= 1'h0;
		else if (_0000_)
			\mchip.state [2] <= _0139_;
	always @(posedge io_in[12])
		if (_0002_)
			\mchip.state [3] <= 1'h0;
		else if (_0000_)
			\mchip.state [3] <= _0140_;
	always @(posedge io_in[12])
		if (_0002_)
			\mchip.state [6] <= 1'h0;
		else if (_0000_)
			\mchip.state [6] <= _0141_;
	reg \mchip.byte_out_reg[0] ;
	always @(posedge io_in[12])
		if (_0137_)
			\mchip.byte_out_reg[0]  <= _1740_;
	assign \mchip.byte_out [0] = \mchip.byte_out_reg[0] ;
	assign io_out = {5'h00, \mchip.is_active , 7'h00, \mchip.byte_out [0]};
	assign \mchip.byte_in  = io_in[7:0];
	assign \mchip.byte_out [7:1] = 7'h00;
	assign \mchip.clock  = io_in[12];
	assign \mchip.io_in  = io_in[11:0];
	assign \mchip.io_out  = {3'h0, \mchip.is_active , 7'h00, \mchip.byte_out [0]};
	assign \mchip.key_in  = io_in[8];
	assign \mchip.plaintext_in  = io_in[9];
	assign \mchip.reset  = io_in[13];
	assign \mchip.sbox.s  = 8'h82;
	assign \mchip.sbox.sbox_in  = 8'h00;
	assign \mchip.sbox.sbox_out  = 8'h82;
	assign \mchip.sbox.t  = 68'h00000000000000000;
	assign \mchip.sbox.u  = 8'h00;
	assign \mchip.sbox.y  = 22'h000000;
	assign \mchip.sbox.z  = 18'h00000;
	assign \mchip.sbox_out  = 8'h82;
	assign \mchip.start  = io_in[10];
endmodule
module d05_meta_info (
	io_in,
	io_out
);
	wire _00000_;
	wire _00001_;
	wire _00002_;
	wire _00003_;
	wire _00004_;
	wire _00005_;
	wire _00006_;
	wire _00007_;
	wire _00008_;
	wire _00009_;
	wire _00010_;
	wire _00011_;
	wire _00012_;
	wire _00013_;
	wire _00014_;
	wire _00015_;
	wire _00016_;
	wire _00017_;
	wire _00018_;
	wire _00019_;
	wire _00020_;
	wire _00021_;
	wire _00022_;
	wire _00023_;
	wire _00024_;
	wire _00025_;
	wire _00026_;
	wire _00027_;
	wire _00028_;
	wire _00029_;
	wire _00030_;
	wire _00031_;
	wire _00032_;
	wire _00033_;
	wire _00034_;
	wire _00035_;
	wire _00036_;
	wire _00037_;
	wire _00038_;
	wire _00039_;
	wire _00040_;
	wire _00041_;
	wire _00042_;
	wire _00043_;
	wire _00044_;
	wire _00045_;
	wire _00046_;
	wire _00047_;
	wire _00048_;
	wire _00049_;
	wire _00050_;
	wire _00051_;
	wire _00052_;
	wire _00053_;
	wire _00054_;
	wire _00055_;
	wire _00056_;
	wire _00057_;
	wire _00058_;
	wire _00059_;
	wire _00060_;
	wire _00061_;
	wire _00062_;
	wire _00063_;
	wire _00064_;
	wire _00065_;
	wire _00066_;
	wire _00067_;
	wire _00068_;
	wire _00069_;
	wire _00070_;
	wire _00071_;
	wire _00072_;
	wire _00073_;
	wire _00074_;
	wire _00075_;
	wire _00076_;
	wire _00077_;
	wire _00078_;
	wire _00079_;
	wire _00080_;
	wire _00081_;
	wire _00082_;
	wire _00083_;
	wire _00084_;
	wire _00085_;
	wire _00086_;
	wire _00087_;
	wire _00088_;
	wire _00089_;
	wire _00090_;
	wire _00091_;
	wire _00092_;
	wire _00093_;
	wire _00094_;
	wire _00095_;
	wire _00096_;
	wire _00097_;
	wire _00098_;
	wire _00099_;
	wire _00100_;
	wire _00101_;
	wire _00102_;
	wire _00103_;
	wire _00104_;
	wire _00105_;
	wire _00106_;
	wire _00107_;
	wire _00108_;
	wire _00109_;
	wire _00110_;
	wire _00111_;
	wire _00112_;
	wire _00113_;
	wire _00114_;
	wire _00115_;
	wire _00116_;
	wire _00117_;
	wire _00118_;
	wire _00119_;
	wire _00120_;
	wire _00121_;
	wire _00122_;
	wire _00123_;
	wire _00124_;
	wire _00125_;
	wire _00126_;
	wire _00127_;
	wire _00128_;
	wire _00129_;
	wire _00130_;
	wire _00131_;
	wire _00132_;
	wire _00133_;
	wire _00134_;
	wire _00135_;
	wire _00136_;
	wire _00137_;
	wire _00138_;
	wire _00139_;
	wire _00140_;
	wire _00141_;
	wire _00142_;
	wire _00143_;
	wire _00144_;
	wire _00145_;
	wire _00146_;
	wire _00147_;
	wire _00148_;
	wire _00149_;
	wire _00150_;
	wire _00151_;
	wire _00152_;
	wire _00153_;
	wire _00154_;
	wire _00155_;
	wire _00156_;
	wire _00157_;
	wire _00158_;
	wire _00159_;
	wire _00160_;
	wire _00161_;
	wire _00162_;
	wire _00163_;
	wire _00164_;
	wire _00165_;
	wire _00166_;
	wire _00167_;
	wire _00168_;
	wire _00169_;
	wire _00170_;
	wire _00171_;
	wire _00172_;
	wire _00173_;
	wire _00174_;
	wire _00175_;
	wire _00176_;
	wire _00177_;
	wire _00178_;
	wire _00179_;
	wire _00180_;
	wire _00181_;
	wire _00182_;
	wire _00183_;
	wire _00184_;
	wire _00185_;
	wire _00186_;
	wire _00187_;
	wire _00188_;
	wire _00189_;
	wire _00190_;
	wire _00191_;
	wire _00192_;
	wire _00193_;
	wire _00194_;
	wire _00195_;
	wire _00196_;
	wire _00197_;
	wire _00198_;
	wire _00199_;
	wire _00200_;
	wire _00201_;
	wire _00202_;
	wire _00203_;
	wire _00204_;
	wire _00205_;
	wire _00206_;
	wire _00207_;
	wire _00208_;
	wire _00209_;
	wire _00210_;
	wire _00211_;
	wire _00212_;
	wire _00213_;
	wire _00214_;
	wire _00215_;
	wire _00216_;
	wire _00217_;
	wire _00218_;
	wire _00219_;
	wire _00220_;
	wire _00221_;
	wire _00222_;
	wire _00223_;
	wire _00224_;
	wire _00225_;
	wire _00226_;
	wire _00227_;
	wire _00228_;
	wire _00229_;
	wire _00230_;
	wire _00231_;
	wire _00232_;
	wire _00233_;
	wire _00234_;
	wire _00235_;
	wire _00236_;
	wire _00237_;
	wire _00238_;
	wire _00239_;
	wire _00240_;
	wire _00241_;
	wire _00242_;
	wire _00243_;
	wire _00244_;
	wire _00245_;
	wire _00246_;
	wire _00247_;
	wire _00248_;
	wire _00249_;
	wire _00250_;
	wire _00251_;
	wire _00252_;
	wire _00253_;
	wire _00254_;
	wire _00255_;
	wire _00256_;
	wire _00257_;
	wire _00258_;
	wire _00259_;
	wire _00260_;
	wire _00261_;
	wire _00262_;
	wire _00263_;
	wire _00264_;
	wire _00265_;
	wire _00266_;
	wire _00267_;
	wire _00268_;
	wire _00269_;
	wire _00270_;
	wire _00271_;
	wire _00272_;
	wire _00273_;
	wire _00274_;
	wire _00275_;
	wire _00276_;
	wire _00277_;
	wire _00278_;
	wire _00279_;
	wire _00280_;
	wire _00281_;
	wire _00282_;
	wire _00283_;
	wire _00284_;
	wire _00285_;
	wire _00286_;
	wire _00287_;
	wire _00288_;
	wire _00289_;
	wire _00290_;
	wire _00291_;
	wire _00292_;
	wire _00293_;
	wire _00294_;
	wire _00295_;
	wire _00296_;
	wire _00297_;
	wire _00298_;
	wire _00299_;
	wire _00300_;
	wire _00301_;
	wire _00302_;
	wire _00303_;
	wire _00304_;
	wire _00305_;
	wire _00306_;
	wire _00307_;
	wire _00308_;
	wire _00309_;
	wire _00310_;
	wire _00311_;
	wire _00312_;
	wire _00313_;
	wire _00314_;
	wire _00315_;
	wire _00316_;
	wire _00317_;
	wire _00318_;
	wire _00319_;
	wire _00320_;
	wire _00321_;
	wire _00322_;
	wire _00323_;
	wire _00324_;
	wire _00325_;
	wire _00326_;
	wire _00327_;
	wire _00328_;
	wire _00329_;
	wire _00330_;
	wire _00331_;
	wire _00332_;
	wire _00333_;
	wire _00334_;
	wire _00335_;
	wire _00336_;
	wire _00337_;
	wire _00338_;
	wire _00339_;
	wire _00340_;
	wire _00341_;
	wire _00342_;
	wire _00343_;
	wire _00344_;
	wire _00345_;
	wire _00346_;
	wire _00347_;
	wire _00348_;
	wire _00349_;
	wire _00350_;
	wire _00351_;
	wire _00352_;
	wire _00353_;
	wire _00354_;
	wire _00355_;
	wire _00356_;
	wire _00357_;
	wire _00358_;
	wire _00359_;
	wire _00360_;
	wire _00361_;
	wire _00362_;
	wire _00363_;
	wire _00364_;
	wire _00365_;
	wire _00366_;
	wire _00367_;
	wire _00368_;
	wire _00369_;
	wire _00370_;
	wire _00371_;
	wire _00372_;
	wire _00373_;
	wire _00374_;
	wire _00375_;
	wire _00376_;
	wire _00377_;
	wire _00378_;
	wire _00379_;
	wire _00380_;
	wire _00381_;
	wire _00382_;
	wire _00383_;
	wire _00384_;
	wire _00385_;
	wire _00386_;
	wire _00387_;
	wire _00388_;
	wire _00389_;
	wire _00390_;
	wire _00391_;
	wire _00392_;
	wire _00393_;
	wire _00394_;
	wire _00395_;
	wire _00396_;
	wire _00397_;
	wire _00398_;
	wire _00399_;
	wire _00400_;
	wire _00401_;
	wire _00402_;
	wire _00403_;
	wire _00404_;
	wire _00405_;
	wire _00406_;
	wire _00407_;
	wire _00408_;
	wire _00409_;
	wire _00410_;
	wire _00411_;
	wire _00412_;
	wire _00413_;
	wire _00414_;
	wire _00415_;
	wire _00416_;
	wire _00417_;
	wire _00418_;
	wire _00419_;
	wire _00420_;
	wire _00421_;
	wire _00422_;
	wire _00423_;
	wire _00424_;
	wire _00425_;
	wire _00426_;
	wire _00427_;
	wire _00428_;
	wire _00429_;
	wire _00430_;
	wire _00431_;
	wire _00432_;
	wire _00433_;
	wire _00434_;
	wire _00435_;
	wire _00436_;
	wire _00437_;
	wire _00438_;
	wire _00439_;
	wire _00440_;
	wire _00441_;
	wire _00442_;
	wire _00443_;
	wire _00444_;
	wire _00445_;
	wire _00446_;
	wire _00447_;
	wire _00448_;
	wire _00449_;
	wire _00450_;
	wire _00451_;
	wire _00452_;
	wire _00453_;
	wire _00454_;
	wire _00455_;
	wire _00456_;
	wire _00457_;
	wire _00458_;
	wire _00459_;
	wire _00460_;
	wire _00461_;
	wire _00462_;
	wire _00463_;
	wire _00464_;
	wire _00465_;
	wire _00466_;
	wire _00467_;
	wire _00468_;
	wire _00469_;
	wire _00470_;
	wire _00471_;
	wire _00472_;
	wire _00473_;
	wire _00474_;
	wire _00475_;
	wire _00476_;
	wire _00477_;
	wire _00478_;
	wire _00479_;
	wire _00480_;
	wire _00481_;
	wire _00482_;
	wire _00483_;
	wire _00484_;
	wire _00485_;
	wire _00486_;
	wire _00487_;
	wire _00488_;
	wire _00489_;
	wire _00490_;
	wire _00491_;
	wire _00492_;
	wire _00493_;
	wire _00494_;
	wire _00495_;
	wire _00496_;
	wire _00497_;
	wire _00498_;
	wire _00499_;
	wire _00500_;
	wire _00501_;
	wire _00502_;
	wire _00503_;
	wire _00504_;
	wire _00505_;
	wire _00506_;
	wire _00507_;
	wire _00508_;
	wire _00509_;
	wire _00510_;
	wire _00511_;
	wire _00512_;
	wire _00513_;
	wire _00514_;
	wire _00515_;
	wire _00516_;
	wire _00517_;
	wire _00518_;
	wire _00519_;
	wire _00520_;
	wire _00521_;
	wire _00522_;
	wire _00523_;
	wire _00524_;
	wire _00525_;
	wire _00526_;
	wire _00527_;
	wire _00528_;
	wire _00529_;
	wire _00530_;
	wire _00531_;
	wire _00532_;
	wire _00533_;
	wire _00534_;
	wire _00535_;
	wire _00536_;
	wire _00537_;
	wire _00538_;
	wire _00539_;
	wire _00540_;
	wire _00541_;
	wire _00542_;
	wire _00543_;
	wire _00544_;
	wire _00545_;
	wire _00546_;
	wire _00547_;
	wire _00548_;
	wire _00549_;
	wire _00550_;
	wire _00551_;
	wire _00552_;
	wire _00553_;
	wire _00554_;
	wire _00555_;
	wire _00556_;
	wire _00557_;
	wire _00558_;
	wire _00559_;
	wire _00560_;
	wire _00561_;
	wire _00562_;
	wire _00563_;
	wire _00564_;
	wire _00565_;
	wire _00566_;
	wire _00567_;
	wire _00568_;
	wire _00569_;
	wire _00570_;
	wire _00571_;
	wire _00572_;
	wire _00573_;
	wire _00574_;
	wire _00575_;
	wire _00576_;
	wire _00577_;
	wire _00578_;
	wire _00579_;
	wire _00580_;
	wire _00581_;
	wire _00582_;
	wire _00583_;
	wire _00584_;
	wire _00585_;
	wire _00586_;
	wire _00587_;
	wire _00588_;
	wire _00589_;
	wire _00590_;
	wire _00591_;
	wire _00592_;
	wire _00593_;
	wire _00594_;
	wire _00595_;
	wire _00596_;
	wire _00597_;
	wire _00598_;
	wire _00599_;
	wire _00600_;
	wire _00601_;
	wire _00602_;
	wire _00603_;
	wire _00604_;
	wire _00605_;
	wire _00606_;
	wire _00607_;
	wire _00608_;
	wire _00609_;
	wire _00610_;
	wire _00611_;
	wire _00612_;
	wire _00613_;
	wire _00614_;
	wire _00615_;
	wire _00616_;
	wire _00617_;
	wire _00618_;
	wire _00619_;
	wire _00620_;
	wire _00621_;
	wire _00622_;
	wire _00623_;
	wire _00624_;
	wire _00625_;
	wire _00626_;
	wire _00627_;
	wire _00628_;
	wire _00629_;
	wire _00630_;
	wire _00631_;
	wire _00632_;
	wire _00633_;
	wire _00634_;
	wire _00635_;
	wire _00636_;
	wire _00637_;
	wire _00638_;
	wire _00639_;
	wire _00640_;
	wire _00641_;
	wire _00642_;
	wire _00643_;
	wire _00644_;
	wire _00645_;
	wire _00646_;
	wire _00647_;
	wire _00648_;
	wire _00649_;
	wire _00650_;
	wire _00651_;
	wire _00652_;
	wire _00653_;
	wire _00654_;
	wire _00655_;
	wire _00656_;
	wire _00657_;
	wire _00658_;
	wire _00659_;
	wire _00660_;
	wire _00661_;
	wire _00662_;
	wire _00663_;
	wire _00664_;
	wire _00665_;
	wire _00666_;
	wire _00667_;
	wire _00668_;
	wire _00669_;
	wire _00670_;
	wire _00671_;
	wire _00672_;
	wire _00673_;
	wire _00674_;
	wire _00675_;
	wire _00676_;
	wire _00677_;
	wire _00678_;
	wire _00679_;
	wire _00680_;
	wire _00681_;
	wire _00682_;
	wire _00683_;
	wire _00684_;
	wire _00685_;
	wire _00686_;
	wire _00687_;
	wire _00688_;
	wire _00689_;
	wire _00690_;
	wire _00691_;
	wire _00692_;
	wire _00693_;
	wire _00694_;
	wire _00695_;
	wire _00696_;
	wire _00697_;
	wire _00698_;
	wire _00699_;
	wire _00700_;
	wire _00701_;
	wire _00702_;
	wire _00703_;
	wire _00704_;
	wire _00705_;
	wire _00706_;
	wire _00707_;
	wire _00708_;
	wire _00709_;
	wire _00710_;
	wire _00711_;
	wire _00712_;
	wire _00713_;
	wire _00714_;
	wire _00715_;
	wire _00716_;
	wire _00717_;
	wire _00718_;
	wire _00719_;
	wire _00720_;
	wire _00721_;
	wire _00722_;
	wire _00723_;
	wire _00724_;
	wire _00725_;
	wire _00726_;
	wire _00727_;
	wire _00728_;
	wire _00729_;
	wire _00730_;
	wire _00731_;
	wire _00732_;
	wire _00733_;
	wire _00734_;
	wire _00735_;
	wire _00736_;
	wire _00737_;
	wire _00738_;
	wire _00739_;
	wire _00740_;
	wire _00741_;
	wire _00742_;
	wire _00743_;
	wire _00744_;
	wire _00745_;
	wire _00746_;
	wire _00747_;
	wire _00748_;
	wire _00749_;
	wire _00750_;
	wire _00751_;
	wire _00752_;
	wire _00753_;
	wire _00754_;
	wire _00755_;
	wire _00756_;
	wire _00757_;
	wire _00758_;
	wire _00759_;
	wire _00760_;
	wire _00761_;
	wire _00762_;
	wire _00763_;
	wire _00764_;
	wire _00765_;
	wire _00766_;
	wire _00767_;
	wire _00768_;
	wire _00769_;
	wire _00770_;
	wire _00771_;
	wire _00772_;
	wire _00773_;
	wire _00774_;
	wire _00775_;
	wire _00776_;
	wire _00777_;
	wire _00778_;
	wire _00779_;
	wire _00780_;
	wire _00781_;
	wire _00782_;
	wire _00783_;
	wire _00784_;
	wire _00785_;
	wire _00786_;
	wire _00787_;
	wire _00788_;
	wire _00789_;
	wire _00790_;
	wire _00791_;
	wire _00792_;
	wire _00793_;
	wire _00794_;
	wire _00795_;
	wire _00796_;
	wire _00797_;
	wire _00798_;
	wire _00799_;
	wire _00800_;
	wire _00801_;
	wire _00802_;
	wire _00803_;
	wire _00804_;
	wire _00805_;
	wire _00806_;
	wire _00807_;
	wire _00808_;
	wire _00809_;
	wire _00810_;
	wire _00811_;
	wire _00812_;
	wire _00813_;
	wire _00814_;
	wire _00815_;
	wire _00816_;
	wire _00817_;
	wire _00818_;
	wire _00819_;
	wire _00820_;
	wire _00821_;
	wire _00822_;
	wire _00823_;
	wire _00824_;
	wire _00825_;
	wire _00826_;
	wire _00827_;
	wire _00828_;
	wire _00829_;
	wire _00830_;
	wire _00831_;
	wire _00832_;
	wire _00833_;
	wire _00834_;
	wire _00835_;
	wire _00836_;
	wire _00837_;
	wire _00838_;
	wire _00839_;
	wire _00840_;
	wire _00841_;
	wire _00842_;
	wire _00843_;
	wire _00844_;
	wire _00845_;
	wire _00846_;
	wire _00847_;
	wire _00848_;
	wire _00849_;
	wire _00850_;
	wire _00851_;
	wire _00852_;
	wire _00853_;
	wire _00854_;
	wire _00855_;
	wire _00856_;
	wire _00857_;
	wire _00858_;
	wire _00859_;
	wire _00860_;
	wire _00861_;
	wire _00862_;
	wire _00863_;
	wire _00864_;
	wire _00865_;
	wire _00866_;
	wire _00867_;
	wire _00868_;
	wire _00869_;
	wire _00870_;
	wire _00871_;
	wire _00872_;
	wire _00873_;
	wire _00874_;
	wire _00875_;
	wire _00876_;
	wire _00877_;
	wire _00878_;
	wire _00879_;
	wire _00880_;
	wire _00881_;
	wire _00882_;
	wire _00883_;
	wire _00884_;
	wire _00885_;
	wire _00886_;
	wire _00887_;
	wire _00888_;
	wire _00889_;
	wire _00890_;
	wire _00891_;
	wire _00892_;
	wire _00893_;
	wire _00894_;
	wire _00895_;
	wire _00896_;
	wire _00897_;
	wire _00898_;
	wire _00899_;
	wire _00900_;
	wire _00901_;
	wire _00902_;
	wire _00903_;
	wire _00904_;
	wire _00905_;
	wire _00906_;
	wire _00907_;
	wire _00908_;
	wire _00909_;
	wire _00910_;
	wire _00911_;
	wire _00912_;
	wire _00913_;
	wire _00914_;
	wire _00915_;
	wire _00916_;
	wire _00917_;
	wire _00918_;
	wire _00919_;
	wire _00920_;
	wire _00921_;
	wire _00922_;
	wire _00923_;
	wire _00924_;
	wire _00925_;
	wire _00926_;
	wire _00927_;
	wire _00928_;
	wire _00929_;
	wire _00930_;
	wire _00931_;
	wire _00932_;
	wire _00933_;
	wire _00934_;
	wire _00935_;
	wire _00936_;
	wire _00937_;
	wire _00938_;
	wire _00939_;
	wire _00940_;
	wire _00941_;
	wire _00942_;
	wire _00943_;
	wire _00944_;
	wire _00945_;
	wire _00946_;
	wire _00947_;
	wire _00948_;
	wire _00949_;
	wire _00950_;
	wire _00951_;
	wire _00952_;
	wire _00953_;
	wire _00954_;
	wire _00955_;
	wire _00956_;
	wire _00957_;
	wire _00958_;
	wire _00959_;
	wire _00960_;
	wire _00961_;
	wire _00962_;
	wire _00963_;
	wire _00964_;
	wire _00965_;
	wire _00966_;
	wire _00967_;
	wire _00968_;
	wire _00969_;
	wire _00970_;
	wire _00971_;
	wire _00972_;
	wire _00973_;
	wire _00974_;
	wire _00975_;
	wire _00976_;
	wire _00977_;
	wire _00978_;
	wire _00979_;
	wire _00980_;
	wire _00981_;
	wire _00982_;
	wire _00983_;
	wire _00984_;
	wire _00985_;
	wire _00986_;
	wire _00987_;
	wire _00988_;
	wire _00989_;
	wire _00990_;
	wire _00991_;
	wire _00992_;
	wire _00993_;
	wire _00994_;
	wire _00995_;
	wire _00996_;
	wire _00997_;
	wire _00998_;
	wire _00999_;
	wire _01000_;
	wire _01001_;
	wire _01002_;
	wire _01003_;
	wire _01004_;
	wire _01005_;
	wire _01006_;
	wire _01007_;
	wire _01008_;
	wire _01009_;
	wire _01010_;
	wire _01011_;
	wire _01012_;
	wire _01013_;
	wire _01014_;
	wire _01015_;
	wire _01016_;
	wire _01017_;
	wire _01018_;
	wire _01019_;
	wire _01020_;
	wire _01021_;
	wire _01022_;
	wire _01023_;
	wire _01024_;
	wire _01025_;
	wire _01026_;
	wire _01027_;
	wire _01028_;
	wire _01029_;
	wire _01030_;
	wire _01031_;
	wire _01032_;
	wire _01033_;
	wire _01034_;
	wire _01035_;
	wire _01036_;
	wire _01037_;
	wire _01038_;
	wire _01039_;
	wire _01040_;
	wire _01041_;
	wire _01042_;
	wire _01043_;
	wire _01044_;
	wire _01045_;
	wire _01046_;
	wire _01047_;
	wire _01048_;
	wire _01049_;
	wire _01050_;
	wire _01051_;
	wire _01052_;
	wire _01053_;
	wire _01054_;
	wire _01055_;
	wire _01056_;
	wire _01057_;
	wire _01058_;
	wire _01059_;
	wire _01060_;
	wire _01061_;
	wire _01062_;
	wire _01063_;
	wire _01064_;
	wire _01065_;
	wire _01066_;
	wire _01067_;
	wire _01068_;
	wire _01069_;
	wire _01070_;
	wire _01071_;
	wire _01072_;
	wire _01073_;
	wire _01074_;
	wire _01075_;
	wire _01076_;
	wire _01077_;
	wire _01078_;
	wire _01079_;
	wire _01080_;
	wire _01081_;
	wire _01082_;
	wire _01083_;
	wire _01084_;
	wire _01085_;
	wire _01086_;
	wire _01087_;
	wire _01088_;
	wire _01089_;
	wire _01090_;
	wire _01091_;
	wire _01092_;
	wire _01093_;
	wire _01094_;
	wire _01095_;
	wire _01096_;
	wire _01097_;
	wire _01098_;
	wire _01099_;
	wire _01100_;
	wire _01101_;
	wire _01102_;
	wire _01103_;
	wire _01104_;
	wire _01105_;
	wire _01106_;
	wire _01107_;
	wire _01108_;
	wire _01109_;
	wire _01110_;
	wire _01111_;
	wire _01112_;
	wire _01113_;
	wire _01114_;
	wire _01115_;
	wire _01116_;
	wire _01117_;
	wire _01118_;
	wire _01119_;
	wire _01120_;
	wire _01121_;
	wire _01122_;
	wire _01123_;
	wire _01124_;
	wire _01125_;
	wire _01126_;
	wire _01127_;
	wire _01128_;
	wire _01129_;
	wire _01130_;
	wire _01131_;
	wire _01132_;
	wire _01133_;
	wire _01134_;
	wire _01135_;
	wire _01136_;
	wire _01137_;
	wire _01138_;
	wire _01139_;
	wire _01140_;
	wire _01141_;
	wire _01142_;
	wire _01143_;
	wire _01144_;
	wire _01145_;
	wire _01146_;
	wire _01147_;
	wire _01148_;
	wire _01149_;
	wire _01150_;
	wire _01151_;
	wire _01152_;
	wire _01153_;
	wire _01154_;
	wire _01155_;
	wire _01156_;
	wire _01157_;
	wire _01158_;
	wire _01159_;
	wire _01160_;
	wire _01161_;
	wire _01162_;
	wire _01163_;
	wire _01164_;
	wire _01165_;
	wire _01166_;
	wire _01167_;
	wire _01168_;
	wire _01169_;
	wire _01170_;
	wire _01171_;
	wire _01172_;
	wire _01173_;
	wire _01174_;
	wire _01175_;
	wire _01176_;
	wire _01177_;
	wire _01178_;
	wire _01179_;
	wire _01180_;
	wire _01181_;
	wire _01182_;
	wire _01183_;
	wire _01184_;
	wire _01185_;
	wire _01186_;
	wire _01187_;
	wire _01188_;
	wire _01189_;
	wire _01190_;
	wire _01191_;
	wire _01192_;
	wire _01193_;
	wire _01194_;
	wire _01195_;
	wire _01196_;
	wire _01197_;
	wire _01198_;
	wire _01199_;
	wire _01200_;
	wire _01201_;
	wire _01202_;
	wire _01203_;
	wire _01204_;
	wire _01205_;
	wire _01206_;
	wire _01207_;
	wire _01208_;
	wire _01209_;
	wire _01210_;
	wire _01211_;
	wire _01212_;
	wire _01213_;
	wire _01214_;
	wire _01215_;
	wire _01216_;
	wire _01217_;
	wire _01218_;
	wire _01219_;
	wire _01220_;
	wire _01221_;
	wire _01222_;
	wire _01223_;
	wire _01224_;
	wire _01225_;
	wire _01226_;
	wire _01227_;
	wire _01228_;
	wire _01229_;
	wire _01230_;
	wire _01231_;
	wire _01232_;
	wire _01233_;
	wire _01234_;
	wire _01235_;
	wire _01236_;
	wire _01237_;
	wire _01238_;
	wire _01239_;
	wire _01240_;
	wire _01241_;
	wire _01242_;
	wire _01243_;
	wire _01244_;
	wire _01245_;
	wire _01246_;
	wire _01247_;
	wire _01248_;
	wire _01249_;
	wire _01250_;
	wire _01251_;
	wire _01252_;
	wire _01253_;
	wire _01254_;
	wire _01255_;
	wire _01256_;
	wire _01257_;
	wire _01258_;
	wire _01259_;
	wire _01260_;
	wire _01261_;
	wire _01262_;
	wire _01263_;
	wire _01264_;
	wire _01265_;
	wire _01266_;
	wire _01267_;
	wire _01268_;
	wire _01269_;
	wire _01270_;
	wire _01271_;
	wire _01272_;
	wire _01273_;
	wire _01274_;
	wire _01275_;
	wire _01276_;
	wire _01277_;
	wire _01278_;
	wire _01279_;
	wire _01280_;
	wire _01281_;
	wire _01282_;
	wire _01283_;
	wire _01284_;
	wire _01285_;
	wire _01286_;
	wire _01287_;
	wire _01288_;
	wire _01289_;
	wire _01290_;
	wire _01291_;
	wire _01292_;
	wire _01293_;
	wire _01294_;
	wire _01295_;
	wire _01296_;
	wire _01297_;
	wire _01298_;
	wire _01299_;
	wire _01300_;
	wire _01301_;
	wire _01302_;
	wire _01303_;
	wire _01304_;
	wire _01305_;
	wire _01306_;
	wire _01307_;
	wire _01308_;
	wire _01309_;
	wire _01310_;
	wire _01311_;
	wire _01312_;
	wire _01313_;
	wire _01314_;
	wire _01315_;
	wire _01316_;
	wire _01317_;
	wire _01318_;
	wire _01319_;
	wire _01320_;
	wire _01321_;
	wire _01322_;
	wire _01323_;
	wire _01324_;
	wire _01325_;
	wire _01326_;
	wire _01327_;
	wire _01328_;
	wire _01329_;
	wire _01330_;
	wire _01331_;
	wire _01332_;
	wire _01333_;
	wire _01334_;
	wire _01335_;
	wire _01336_;
	wire _01337_;
	wire _01338_;
	wire _01339_;
	wire _01340_;
	wire _01341_;
	wire _01342_;
	wire _01343_;
	wire _01344_;
	wire _01345_;
	wire _01346_;
	wire _01347_;
	wire _01348_;
	wire _01349_;
	wire _01350_;
	wire _01351_;
	wire _01352_;
	wire _01353_;
	wire _01354_;
	wire _01355_;
	wire _01356_;
	wire _01357_;
	wire _01358_;
	wire _01359_;
	wire _01360_;
	wire _01361_;
	wire _01362_;
	wire _01363_;
	wire _01364_;
	wire _01365_;
	wire _01366_;
	wire _01367_;
	wire _01368_;
	wire _01369_;
	wire _01370_;
	wire _01371_;
	wire _01372_;
	wire _01373_;
	wire _01374_;
	wire _01375_;
	wire _01376_;
	wire _01377_;
	wire _01378_;
	wire _01379_;
	wire _01380_;
	wire _01381_;
	wire _01382_;
	wire _01383_;
	wire _01384_;
	wire _01385_;
	wire _01386_;
	wire _01387_;
	wire _01388_;
	wire _01389_;
	wire _01390_;
	wire _01391_;
	wire _01392_;
	wire _01393_;
	wire _01394_;
	wire _01395_;
	wire _01396_;
	wire _01397_;
	wire _01398_;
	wire _01399_;
	wire _01400_;
	wire _01401_;
	wire _01402_;
	wire _01403_;
	wire _01404_;
	wire _01405_;
	wire _01406_;
	wire _01407_;
	wire _01408_;
	wire _01409_;
	wire _01410_;
	wire _01411_;
	wire _01412_;
	wire _01413_;
	wire _01414_;
	wire _01415_;
	wire _01416_;
	wire _01417_;
	wire _01418_;
	wire _01419_;
	wire _01420_;
	wire _01421_;
	wire _01422_;
	wire _01423_;
	wire _01424_;
	wire _01425_;
	wire _01426_;
	wire _01427_;
	wire _01428_;
	wire _01429_;
	wire _01430_;
	wire _01431_;
	wire _01432_;
	wire _01433_;
	wire _01434_;
	wire _01435_;
	wire _01436_;
	wire _01437_;
	wire _01438_;
	wire _01439_;
	wire _01440_;
	wire _01441_;
	wire _01442_;
	wire _01443_;
	wire _01444_;
	wire _01445_;
	wire _01446_;
	wire _01447_;
	wire _01448_;
	wire _01449_;
	wire _01450_;
	wire _01451_;
	wire _01452_;
	wire _01453_;
	wire _01454_;
	wire _01455_;
	wire _01456_;
	wire _01457_;
	wire _01458_;
	wire _01459_;
	wire _01460_;
	wire _01461_;
	wire _01462_;
	wire _01463_;
	wire _01464_;
	wire _01465_;
	wire _01466_;
	wire _01467_;
	wire _01468_;
	wire _01469_;
	wire _01470_;
	wire _01471_;
	wire _01472_;
	wire _01473_;
	wire _01474_;
	wire _01475_;
	wire _01476_;
	wire _01477_;
	wire _01478_;
	wire _01479_;
	wire _01480_;
	wire _01481_;
	wire _01482_;
	wire _01483_;
	wire _01484_;
	wire _01485_;
	wire _01486_;
	wire _01487_;
	wire _01488_;
	wire _01489_;
	wire _01490_;
	wire _01491_;
	wire _01492_;
	wire _01493_;
	wire _01494_;
	wire _01495_;
	wire _01496_;
	wire _01497_;
	wire _01498_;
	wire _01499_;
	wire _01500_;
	wire _01501_;
	wire _01502_;
	wire _01503_;
	wire _01504_;
	wire _01505_;
	wire _01506_;
	wire _01507_;
	wire _01508_;
	wire _01509_;
	wire _01510_;
	wire _01511_;
	wire _01512_;
	wire _01513_;
	wire _01514_;
	wire _01515_;
	wire _01516_;
	wire _01517_;
	wire _01518_;
	wire _01519_;
	wire _01520_;
	wire _01521_;
	wire _01522_;
	wire _01523_;
	wire _01524_;
	wire _01525_;
	wire _01526_;
	wire _01527_;
	wire _01528_;
	wire _01529_;
	wire _01530_;
	wire _01531_;
	wire _01532_;
	wire _01533_;
	wire _01534_;
	wire _01535_;
	wire _01536_;
	wire _01537_;
	wire _01538_;
	wire _01539_;
	wire _01540_;
	wire _01541_;
	wire _01542_;
	wire _01543_;
	wire _01544_;
	wire _01545_;
	wire _01546_;
	wire _01547_;
	wire _01548_;
	wire _01549_;
	wire _01550_;
	wire _01551_;
	wire _01552_;
	wire _01553_;
	wire _01554_;
	wire _01555_;
	wire _01556_;
	wire _01557_;
	wire _01558_;
	wire _01559_;
	wire _01560_;
	wire _01561_;
	wire _01562_;
	wire _01563_;
	wire _01564_;
	wire _01565_;
	wire _01566_;
	wire _01567_;
	wire _01568_;
	wire _01569_;
	wire _01570_;
	wire _01571_;
	wire _01572_;
	wire _01573_;
	wire _01574_;
	wire _01575_;
	wire _01576_;
	wire _01577_;
	wire _01578_;
	wire _01579_;
	wire _01580_;
	wire _01581_;
	wire _01582_;
	wire _01583_;
	wire _01584_;
	wire _01585_;
	wire _01586_;
	wire _01587_;
	wire _01588_;
	wire _01589_;
	wire _01590_;
	wire _01591_;
	wire _01592_;
	wire _01593_;
	wire _01594_;
	wire _01595_;
	wire _01596_;
	wire _01597_;
	wire _01598_;
	wire _01599_;
	wire _01600_;
	wire _01601_;
	wire _01602_;
	wire _01603_;
	wire _01604_;
	wire _01605_;
	wire _01606_;
	wire _01607_;
	wire _01608_;
	wire _01609_;
	wire _01610_;
	wire _01611_;
	wire _01612_;
	wire _01613_;
	wire _01614_;
	wire _01615_;
	wire _01616_;
	wire _01617_;
	wire _01618_;
	wire _01619_;
	wire _01620_;
	wire _01621_;
	wire _01622_;
	wire _01623_;
	wire _01624_;
	wire _01625_;
	wire _01626_;
	wire _01627_;
	wire _01628_;
	wire _01629_;
	wire _01630_;
	wire _01631_;
	wire _01632_;
	wire _01633_;
	wire _01634_;
	wire _01635_;
	wire _01636_;
	wire _01637_;
	wire _01638_;
	wire _01639_;
	wire _01640_;
	wire _01641_;
	wire _01642_;
	wire _01643_;
	wire _01644_;
	wire _01645_;
	wire _01646_;
	wire _01647_;
	wire _01648_;
	wire _01649_;
	wire _01650_;
	wire _01651_;
	wire _01652_;
	wire _01653_;
	wire _01654_;
	wire _01655_;
	wire _01656_;
	wire _01657_;
	wire _01658_;
	wire _01659_;
	wire _01660_;
	wire _01661_;
	wire _01662_;
	wire _01663_;
	wire _01664_;
	wire _01665_;
	wire _01666_;
	wire _01667_;
	wire _01668_;
	wire _01669_;
	wire _01670_;
	wire _01671_;
	wire _01672_;
	wire _01673_;
	wire _01674_;
	wire _01675_;
	wire _01676_;
	wire _01677_;
	wire _01678_;
	wire _01679_;
	wire _01680_;
	wire _01681_;
	wire _01682_;
	wire _01683_;
	wire _01684_;
	wire _01685_;
	wire _01686_;
	wire _01687_;
	wire _01688_;
	wire _01689_;
	wire _01690_;
	wire _01691_;
	wire _01692_;
	wire _01693_;
	wire _01694_;
	wire _01695_;
	wire _01696_;
	wire _01697_;
	wire _01698_;
	wire _01699_;
	wire _01700_;
	wire _01701_;
	wire _01702_;
	wire _01703_;
	wire _01704_;
	wire _01705_;
	wire _01706_;
	wire _01707_;
	wire _01708_;
	wire _01709_;
	wire _01710_;
	wire _01711_;
	wire _01712_;
	wire _01713_;
	wire _01714_;
	wire _01715_;
	wire _01716_;
	wire _01717_;
	wire _01718_;
	wire _01719_;
	wire _01720_;
	wire _01721_;
	wire _01722_;
	wire _01723_;
	wire _01724_;
	wire _01725_;
	wire _01726_;
	wire _01727_;
	wire _01728_;
	wire _01729_;
	wire _01730_;
	wire _01731_;
	wire _01732_;
	wire _01733_;
	wire _01734_;
	wire _01735_;
	wire _01736_;
	wire _01737_;
	wire _01738_;
	wire _01739_;
	wire _01740_;
	wire _01741_;
	wire _01742_;
	wire _01743_;
	wire _01744_;
	wire _01745_;
	wire _01746_;
	wire _01747_;
	wire _01748_;
	wire _01749_;
	wire _01750_;
	wire _01751_;
	wire _01752_;
	wire _01753_;
	wire _01754_;
	wire _01755_;
	wire _01756_;
	wire _01757_;
	wire _01758_;
	wire _01759_;
	wire _01760_;
	wire _01761_;
	wire _01762_;
	wire _01763_;
	wire _01764_;
	wire _01765_;
	wire _01766_;
	wire _01767_;
	wire _01768_;
	wire _01769_;
	wire _01770_;
	wire _01771_;
	wire _01772_;
	wire _01773_;
	wire _01774_;
	wire _01775_;
	wire _01776_;
	wire _01777_;
	wire _01778_;
	wire _01779_;
	wire _01780_;
	wire _01781_;
	wire _01782_;
	wire _01783_;
	wire _01784_;
	wire _01785_;
	wire _01786_;
	wire _01787_;
	wire _01788_;
	wire _01789_;
	wire _01790_;
	wire _01791_;
	wire _01792_;
	wire _01793_;
	wire _01794_;
	wire _01795_;
	wire _01796_;
	wire _01797_;
	wire _01798_;
	wire _01799_;
	wire _01800_;
	wire _01801_;
	wire _01802_;
	wire _01803_;
	wire _01804_;
	wire _01805_;
	wire _01806_;
	wire _01807_;
	wire _01808_;
	wire _01809_;
	wire _01810_;
	wire _01811_;
	wire _01812_;
	wire _01813_;
	wire _01814_;
	wire _01815_;
	wire _01816_;
	wire _01817_;
	wire _01818_;
	wire _01819_;
	wire _01820_;
	wire _01821_;
	wire _01822_;
	wire _01823_;
	wire _01824_;
	wire _01825_;
	wire _01826_;
	wire _01827_;
	wire _01828_;
	wire _01829_;
	wire _01830_;
	wire _01831_;
	wire _01832_;
	wire _01833_;
	wire _01834_;
	wire _01835_;
	wire _01836_;
	wire _01837_;
	wire _01838_;
	wire _01839_;
	wire _01840_;
	wire _01841_;
	wire _01842_;
	wire _01843_;
	wire _01844_;
	wire _01845_;
	wire _01846_;
	wire _01847_;
	wire _01848_;
	wire _01849_;
	wire _01850_;
	wire _01851_;
	wire _01852_;
	wire _01853_;
	wire _01854_;
	wire _01855_;
	wire _01856_;
	wire _01857_;
	wire _01858_;
	wire _01859_;
	wire _01860_;
	wire _01861_;
	wire _01862_;
	wire _01863_;
	wire _01864_;
	wire _01865_;
	wire _01866_;
	wire _01867_;
	wire _01868_;
	wire _01869_;
	wire _01870_;
	wire _01871_;
	wire _01872_;
	wire _01873_;
	wire _01874_;
	wire _01875_;
	wire _01876_;
	wire _01877_;
	wire _01878_;
	wire _01879_;
	wire _01880_;
	wire _01881_;
	wire _01882_;
	wire _01883_;
	wire _01884_;
	wire _01885_;
	wire _01886_;
	wire _01887_;
	wire _01888_;
	wire _01889_;
	wire _01890_;
	wire _01891_;
	wire _01892_;
	wire _01893_;
	wire _01894_;
	wire _01895_;
	wire _01896_;
	wire _01897_;
	wire _01898_;
	wire _01899_;
	wire _01900_;
	wire _01901_;
	wire _01902_;
	wire _01903_;
	wire _01904_;
	wire _01905_;
	wire _01906_;
	wire _01907_;
	wire _01908_;
	wire _01909_;
	wire _01910_;
	wire _01911_;
	wire _01912_;
	wire _01913_;
	wire _01914_;
	wire _01915_;
	wire _01916_;
	wire _01917_;
	wire _01918_;
	wire _01919_;
	wire _01920_;
	wire _01921_;
	wire _01922_;
	wire _01923_;
	wire _01924_;
	wire _01925_;
	wire _01926_;
	wire _01927_;
	wire _01928_;
	wire _01929_;
	wire _01930_;
	wire _01931_;
	wire _01932_;
	wire _01933_;
	wire _01934_;
	wire _01935_;
	wire _01936_;
	wire _01937_;
	wire _01938_;
	wire _01939_;
	wire _01940_;
	wire _01941_;
	wire _01942_;
	wire _01943_;
	wire _01944_;
	wire _01945_;
	wire _01946_;
	wire _01947_;
	wire _01948_;
	wire _01949_;
	wire _01950_;
	wire _01951_;
	wire _01952_;
	wire _01953_;
	wire _01954_;
	wire _01955_;
	wire _01956_;
	wire _01957_;
	wire _01958_;
	wire _01959_;
	wire _01960_;
	wire _01961_;
	wire _01962_;
	wire _01963_;
	wire _01964_;
	wire _01965_;
	wire _01966_;
	wire _01967_;
	wire _01968_;
	wire _01969_;
	wire _01970_;
	wire _01971_;
	wire _01972_;
	wire _01973_;
	wire _01974_;
	wire _01975_;
	wire _01976_;
	wire _01977_;
	wire _01978_;
	wire _01979_;
	wire _01980_;
	wire _01981_;
	wire _01982_;
	wire _01983_;
	wire _01984_;
	wire _01985_;
	wire _01986_;
	wire _01987_;
	wire _01988_;
	wire _01989_;
	wire _01990_;
	wire _01991_;
	wire _01992_;
	wire _01993_;
	wire _01994_;
	wire _01995_;
	wire _01996_;
	wire _01997_;
	wire _01998_;
	wire _01999_;
	wire _02000_;
	wire _02001_;
	wire _02002_;
	wire _02003_;
	wire _02004_;
	wire _02005_;
	wire _02006_;
	wire _02007_;
	wire _02008_;
	wire _02009_;
	wire _02010_;
	wire _02011_;
	wire _02012_;
	wire _02013_;
	wire _02014_;
	wire _02015_;
	wire _02016_;
	wire _02017_;
	wire _02018_;
	wire _02019_;
	wire _02020_;
	wire _02021_;
	wire _02022_;
	wire _02023_;
	wire _02024_;
	wire _02025_;
	wire _02026_;
	wire _02027_;
	wire _02028_;
	wire _02029_;
	wire _02030_;
	wire _02031_;
	wire _02032_;
	wire _02033_;
	wire _02034_;
	wire _02035_;
	wire _02036_;
	wire _02037_;
	wire _02038_;
	wire _02039_;
	wire _02040_;
	wire _02041_;
	wire _02042_;
	wire _02043_;
	wire _02044_;
	wire _02045_;
	wire _02046_;
	wire _02047_;
	wire _02048_;
	wire _02049_;
	wire _02050_;
	wire _02051_;
	wire _02052_;
	wire _02053_;
	wire _02054_;
	wire _02055_;
	wire _02056_;
	wire _02057_;
	wire _02058_;
	wire _02059_;
	wire _02060_;
	wire _02061_;
	wire _02062_;
	wire _02063_;
	wire _02064_;
	wire _02065_;
	wire _02066_;
	wire _02067_;
	wire _02068_;
	wire _02069_;
	wire _02070_;
	wire _02071_;
	wire _02072_;
	wire _02073_;
	wire _02074_;
	wire _02075_;
	wire _02076_;
	wire _02077_;
	wire _02078_;
	wire _02079_;
	wire _02080_;
	wire _02081_;
	wire _02082_;
	wire _02083_;
	wire _02084_;
	wire _02085_;
	wire _02086_;
	wire _02087_;
	wire _02088_;
	wire _02089_;
	wire _02090_;
	wire _02091_;
	wire _02092_;
	wire _02093_;
	wire _02094_;
	wire _02095_;
	wire _02096_;
	wire _02097_;
	wire _02098_;
	wire _02099_;
	wire _02100_;
	wire _02101_;
	wire _02102_;
	wire _02103_;
	wire _02104_;
	wire _02105_;
	wire _02106_;
	wire _02107_;
	wire _02108_;
	wire _02109_;
	wire _02110_;
	wire _02111_;
	wire _02112_;
	wire _02113_;
	wire _02114_;
	wire _02115_;
	wire _02116_;
	wire _02117_;
	wire _02118_;
	wire _02119_;
	wire _02120_;
	wire _02121_;
	wire _02122_;
	wire _02123_;
	wire _02124_;
	wire _02125_;
	wire _02126_;
	wire _02127_;
	wire _02128_;
	wire _02129_;
	wire _02130_;
	wire _02131_;
	wire _02132_;
	wire _02133_;
	wire _02134_;
	wire _02135_;
	wire _02136_;
	wire _02137_;
	wire _02138_;
	wire _02139_;
	wire _02140_;
	wire _02141_;
	wire _02142_;
	wire _02143_;
	wire _02144_;
	wire _02145_;
	wire _02146_;
	wire _02147_;
	wire _02148_;
	wire _02149_;
	wire _02150_;
	wire _02151_;
	wire _02152_;
	wire _02153_;
	wire _02154_;
	wire _02155_;
	wire _02156_;
	wire _02157_;
	wire _02158_;
	wire _02159_;
	wire _02160_;
	wire _02161_;
	wire _02162_;
	wire _02163_;
	wire _02164_;
	wire _02165_;
	wire _02166_;
	wire _02167_;
	wire _02168_;
	wire _02169_;
	wire _02170_;
	wire _02171_;
	wire _02172_;
	wire _02173_;
	wire _02174_;
	wire _02175_;
	wire _02176_;
	wire _02177_;
	wire _02178_;
	wire _02179_;
	wire _02180_;
	wire _02181_;
	wire _02182_;
	wire _02183_;
	wire _02184_;
	wire _02185_;
	wire _02186_;
	wire _02187_;
	wire _02188_;
	wire _02189_;
	wire _02190_;
	wire _02191_;
	wire _02192_;
	wire _02193_;
	wire _02194_;
	wire _02195_;
	wire _02196_;
	wire _02197_;
	wire _02198_;
	wire _02199_;
	wire _02200_;
	wire _02201_;
	wire _02202_;
	wire _02203_;
	wire _02204_;
	wire _02205_;
	wire _02206_;
	wire _02207_;
	wire _02208_;
	wire _02209_;
	wire _02210_;
	wire _02211_;
	wire _02212_;
	wire _02213_;
	wire _02214_;
	wire _02215_;
	wire _02216_;
	wire _02217_;
	wire _02218_;
	wire _02219_;
	wire _02220_;
	wire _02221_;
	wire _02222_;
	wire _02223_;
	wire _02224_;
	wire _02225_;
	wire _02226_;
	wire _02227_;
	wire _02228_;
	wire _02229_;
	wire _02230_;
	wire _02231_;
	wire _02232_;
	wire _02233_;
	wire _02234_;
	wire _02235_;
	wire _02236_;
	wire _02237_;
	wire _02238_;
	wire _02239_;
	wire _02240_;
	wire _02241_;
	wire _02242_;
	wire _02243_;
	wire _02244_;
	wire _02245_;
	wire _02246_;
	wire _02247_;
	wire _02248_;
	wire _02249_;
	wire _02250_;
	wire _02251_;
	wire _02252_;
	wire _02253_;
	wire _02254_;
	wire _02255_;
	wire _02256_;
	wire _02257_;
	wire _02258_;
	wire _02259_;
	wire _02260_;
	wire _02261_;
	wire _02262_;
	wire _02263_;
	wire _02264_;
	wire _02265_;
	wire _02266_;
	wire _02267_;
	wire _02268_;
	wire _02269_;
	wire _02270_;
	wire _02271_;
	wire _02272_;
	wire _02273_;
	wire _02274_;
	wire _02275_;
	wire _02276_;
	wire _02277_;
	wire _02278_;
	wire _02279_;
	wire _02280_;
	wire _02281_;
	wire _02282_;
	wire _02283_;
	wire _02284_;
	wire _02285_;
	wire _02286_;
	wire _02287_;
	wire _02288_;
	wire _02289_;
	wire _02290_;
	wire _02291_;
	wire _02292_;
	wire _02293_;
	wire _02294_;
	wire _02295_;
	wire _02296_;
	wire _02297_;
	wire _02298_;
	wire _02299_;
	wire _02300_;
	wire _02301_;
	wire _02302_;
	wire _02303_;
	wire _02304_;
	wire _02305_;
	wire _02306_;
	wire _02307_;
	wire _02308_;
	wire _02309_;
	wire _02310_;
	wire _02311_;
	wire _02312_;
	wire _02313_;
	wire _02314_;
	wire _02315_;
	wire _02316_;
	wire _02317_;
	wire _02318_;
	wire _02319_;
	wire _02320_;
	wire _02321_;
	wire _02322_;
	wire _02323_;
	wire _02324_;
	wire _02325_;
	wire _02326_;
	wire _02327_;
	wire _02328_;
	wire _02329_;
	wire _02330_;
	wire _02331_;
	wire _02332_;
	wire _02333_;
	wire _02334_;
	wire _02335_;
	wire _02336_;
	wire _02337_;
	wire _02338_;
	wire _02339_;
	wire _02340_;
	wire _02341_;
	wire _02342_;
	wire _02343_;
	wire _02344_;
	wire _02345_;
	wire _02346_;
	wire _02347_;
	wire _02348_;
	wire _02349_;
	wire _02350_;
	wire _02351_;
	wire _02352_;
	wire _02353_;
	wire _02354_;
	wire _02355_;
	wire _02356_;
	wire _02357_;
	wire _02358_;
	wire _02359_;
	wire _02360_;
	wire _02361_;
	wire _02362_;
	wire _02363_;
	wire _02364_;
	wire _02365_;
	wire _02366_;
	wire _02367_;
	wire _02368_;
	wire _02369_;
	wire _02370_;
	wire _02371_;
	wire _02372_;
	wire _02373_;
	wire _02374_;
	wire _02375_;
	wire _02376_;
	wire _02377_;
	wire _02378_;
	wire _02379_;
	wire _02380_;
	wire _02381_;
	wire _02382_;
	wire _02383_;
	wire _02384_;
	wire _02385_;
	wire _02386_;
	wire _02387_;
	wire _02388_;
	wire _02389_;
	wire _02390_;
	wire _02391_;
	wire _02392_;
	wire _02393_;
	wire _02394_;
	wire _02395_;
	wire _02396_;
	wire _02397_;
	wire _02398_;
	wire _02399_;
	wire _02400_;
	wire _02401_;
	wire _02402_;
	wire _02403_;
	wire _02404_;
	wire _02405_;
	wire _02406_;
	wire _02407_;
	wire _02408_;
	wire _02409_;
	wire _02410_;
	wire _02411_;
	wire _02412_;
	wire _02413_;
	wire _02414_;
	wire _02415_;
	wire _02416_;
	wire _02417_;
	wire _02418_;
	wire _02419_;
	wire _02420_;
	wire _02421_;
	wire _02422_;
	wire _02423_;
	wire _02424_;
	wire _02425_;
	wire _02426_;
	wire _02427_;
	wire _02428_;
	wire _02429_;
	wire _02430_;
	wire _02431_;
	wire _02432_;
	wire _02433_;
	wire _02434_;
	wire _02435_;
	wire _02436_;
	wire _02437_;
	wire _02438_;
	wire _02439_;
	wire _02440_;
	wire _02441_;
	wire _02442_;
	wire _02443_;
	wire _02444_;
	wire _02445_;
	wire _02446_;
	wire _02447_;
	wire _02448_;
	wire _02449_;
	wire _02450_;
	wire _02451_;
	wire _02452_;
	wire _02453_;
	wire _02454_;
	wire _02455_;
	wire _02456_;
	wire _02457_;
	wire _02458_;
	wire _02459_;
	wire _02460_;
	wire _02461_;
	wire _02462_;
	wire _02463_;
	wire _02464_;
	wire _02465_;
	wire _02466_;
	wire _02467_;
	wire _02468_;
	wire _02469_;
	wire _02470_;
	wire _02471_;
	wire _02472_;
	wire _02473_;
	wire _02474_;
	wire _02475_;
	wire _02476_;
	wire _02477_;
	wire _02478_;
	wire _02479_;
	wire _02480_;
	wire _02481_;
	wire _02482_;
	wire _02483_;
	wire _02484_;
	wire _02485_;
	wire _02486_;
	wire _02487_;
	wire _02488_;
	wire _02489_;
	wire _02490_;
	wire _02491_;
	wire _02492_;
	wire _02493_;
	wire _02494_;
	wire _02495_;
	wire _02496_;
	wire _02497_;
	wire _02498_;
	wire _02499_;
	wire _02500_;
	wire _02501_;
	wire _02502_;
	wire _02503_;
	wire _02504_;
	wire _02505_;
	wire _02506_;
	wire _02507_;
	wire _02508_;
	wire _02509_;
	wire _02510_;
	wire _02511_;
	wire _02512_;
	wire _02513_;
	wire _02514_;
	wire _02515_;
	wire _02516_;
	wire _02517_;
	wire _02518_;
	wire _02519_;
	wire _02520_;
	wire _02521_;
	wire _02522_;
	wire _02523_;
	wire _02524_;
	wire _02525_;
	wire _02526_;
	wire _02527_;
	wire _02528_;
	wire _02529_;
	wire _02530_;
	wire _02531_;
	wire _02532_;
	wire _02533_;
	wire _02534_;
	wire _02535_;
	wire _02536_;
	wire _02537_;
	wire _02538_;
	wire _02539_;
	wire _02540_;
	wire _02541_;
	wire _02542_;
	wire _02543_;
	wire _02544_;
	wire _02545_;
	wire _02546_;
	wire _02547_;
	wire _02548_;
	wire _02549_;
	wire _02550_;
	wire _02551_;
	wire _02552_;
	wire _02553_;
	wire _02554_;
	wire _02555_;
	wire _02556_;
	wire _02557_;
	wire _02558_;
	wire _02559_;
	wire _02560_;
	wire _02561_;
	wire _02562_;
	wire _02563_;
	wire _02564_;
	wire _02565_;
	wire _02566_;
	wire _02567_;
	wire _02568_;
	wire _02569_;
	wire _02570_;
	wire _02571_;
	wire _02572_;
	wire _02573_;
	wire _02574_;
	wire _02575_;
	wire _02576_;
	wire _02577_;
	wire _02578_;
	wire _02579_;
	wire _02580_;
	wire _02581_;
	wire _02582_;
	wire _02583_;
	wire _02584_;
	wire _02585_;
	wire _02586_;
	wire _02587_;
	wire _02588_;
	wire _02589_;
	wire _02590_;
	wire _02591_;
	wire _02592_;
	wire _02593_;
	wire _02594_;
	wire _02595_;
	wire _02596_;
	wire _02597_;
	wire _02598_;
	wire _02599_;
	wire _02600_;
	wire _02601_;
	wire _02602_;
	wire _02603_;
	wire _02604_;
	wire _02605_;
	wire _02606_;
	wire _02607_;
	wire _02608_;
	wire _02609_;
	wire _02610_;
	wire _02611_;
	wire _02612_;
	wire _02613_;
	wire _02614_;
	wire _02615_;
	wire _02616_;
	wire _02617_;
	wire _02618_;
	wire _02619_;
	wire _02620_;
	wire _02621_;
	wire _02622_;
	wire _02623_;
	wire _02624_;
	wire _02625_;
	wire _02626_;
	wire _02627_;
	wire _02628_;
	wire _02629_;
	wire _02630_;
	wire _02631_;
	wire _02632_;
	wire _02633_;
	wire _02634_;
	wire _02635_;
	wire _02636_;
	wire _02637_;
	wire _02638_;
	wire _02639_;
	wire _02640_;
	wire _02641_;
	wire _02642_;
	wire _02643_;
	wire _02644_;
	wire _02645_;
	wire _02646_;
	wire _02647_;
	wire _02648_;
	wire _02649_;
	wire _02650_;
	wire _02651_;
	wire _02652_;
	wire _02653_;
	wire _02654_;
	wire _02655_;
	wire _02656_;
	wire _02657_;
	wire _02658_;
	wire _02659_;
	wire _02660_;
	wire _02661_;
	wire _02662_;
	wire _02663_;
	wire _02664_;
	wire _02665_;
	wire _02666_;
	wire _02667_;
	wire _02668_;
	wire _02669_;
	wire _02670_;
	wire _02671_;
	wire _02672_;
	wire _02673_;
	wire _02674_;
	wire _02675_;
	wire _02676_;
	wire _02677_;
	wire _02678_;
	wire _02679_;
	wire _02680_;
	wire _02681_;
	wire _02682_;
	wire _02683_;
	wire _02684_;
	wire _02685_;
	wire _02686_;
	wire _02687_;
	wire _02688_;
	wire _02689_;
	wire _02690_;
	wire _02691_;
	wire _02692_;
	wire _02693_;
	wire _02694_;
	wire _02695_;
	wire _02696_;
	wire _02697_;
	wire _02698_;
	wire _02699_;
	wire _02700_;
	wire _02701_;
	wire _02702_;
	wire _02703_;
	wire _02704_;
	wire _02705_;
	wire _02706_;
	wire _02707_;
	wire _02708_;
	wire _02709_;
	wire _02710_;
	wire _02711_;
	wire _02712_;
	wire _02713_;
	wire _02714_;
	wire _02715_;
	wire _02716_;
	wire _02717_;
	wire _02718_;
	wire _02719_;
	wire _02720_;
	wire _02721_;
	wire _02722_;
	wire _02723_;
	wire _02724_;
	wire _02725_;
	wire _02726_;
	wire _02727_;
	wire _02728_;
	wire _02729_;
	wire _02730_;
	wire _02731_;
	wire _02732_;
	wire _02733_;
	wire _02734_;
	wire _02735_;
	wire _02736_;
	wire _02737_;
	wire _02738_;
	wire _02739_;
	wire _02740_;
	wire _02741_;
	wire _02742_;
	wire _02743_;
	wire _02744_;
	wire _02745_;
	wire _02746_;
	wire _02747_;
	wire _02748_;
	wire _02749_;
	wire _02750_;
	wire _02751_;
	wire _02752_;
	wire _02753_;
	wire _02754_;
	wire _02755_;
	wire _02756_;
	wire _02757_;
	wire _02758_;
	wire _02759_;
	wire _02760_;
	wire _02761_;
	wire _02762_;
	wire _02763_;
	wire _02764_;
	wire _02765_;
	wire _02766_;
	wire _02767_;
	wire _02768_;
	wire _02769_;
	wire _02770_;
	wire _02771_;
	wire _02772_;
	wire _02773_;
	wire _02774_;
	wire _02775_;
	wire _02776_;
	wire _02777_;
	wire _02778_;
	wire _02779_;
	wire _02780_;
	wire _02781_;
	wire _02782_;
	wire _02783_;
	wire _02784_;
	wire _02785_;
	wire _02786_;
	wire _02787_;
	wire _02788_;
	wire _02789_;
	wire _02790_;
	wire _02791_;
	wire _02792_;
	wire _02793_;
	wire _02794_;
	wire _02795_;
	wire _02796_;
	wire _02797_;
	wire _02798_;
	wire _02799_;
	wire _02800_;
	wire _02801_;
	wire _02802_;
	wire _02803_;
	wire _02804_;
	wire _02805_;
	wire _02806_;
	wire _02807_;
	wire _02808_;
	wire _02809_;
	wire _02810_;
	wire _02811_;
	wire _02812_;
	wire _02813_;
	wire _02814_;
	wire _02815_;
	wire _02816_;
	wire _02817_;
	wire _02818_;
	wire _02819_;
	wire _02820_;
	wire _02821_;
	wire _02822_;
	wire _02823_;
	wire _02824_;
	wire _02825_;
	wire _02826_;
	wire _02827_;
	wire _02828_;
	wire _02829_;
	wire _02830_;
	wire _02831_;
	wire _02832_;
	wire _02833_;
	wire _02834_;
	wire _02835_;
	wire _02836_;
	wire _02837_;
	wire _02838_;
	wire _02839_;
	wire _02840_;
	wire _02841_;
	wire _02842_;
	wire _02843_;
	wire _02844_;
	wire _02845_;
	wire _02846_;
	wire _02847_;
	wire _02848_;
	wire _02849_;
	wire _02850_;
	wire _02851_;
	wire _02852_;
	wire _02853_;
	wire _02854_;
	wire _02855_;
	wire _02856_;
	wire _02857_;
	wire _02858_;
	wire _02859_;
	wire _02860_;
	wire _02861_;
	wire _02862_;
	wire _02863_;
	wire _02864_;
	wire _02865_;
	wire _02866_;
	wire _02867_;
	wire _02868_;
	wire _02869_;
	wire _02870_;
	wire _02871_;
	wire _02872_;
	wire _02873_;
	wire _02874_;
	wire _02875_;
	wire _02876_;
	wire _02877_;
	wire _02878_;
	wire _02879_;
	wire _02880_;
	wire _02881_;
	wire _02882_;
	wire _02883_;
	wire _02884_;
	wire _02885_;
	wire _02886_;
	wire _02887_;
	wire _02888_;
	wire _02889_;
	wire _02890_;
	wire _02891_;
	wire _02892_;
	wire _02893_;
	wire _02894_;
	wire _02895_;
	wire _02896_;
	wire _02897_;
	wire _02898_;
	wire _02899_;
	wire _02900_;
	wire _02901_;
	wire _02902_;
	wire _02903_;
	wire _02904_;
	wire _02905_;
	wire _02906_;
	wire _02907_;
	wire _02908_;
	wire _02909_;
	wire _02910_;
	wire _02911_;
	wire _02912_;
	wire _02913_;
	wire _02914_;
	wire _02915_;
	wire _02916_;
	wire _02917_;
	wire _02918_;
	wire _02919_;
	wire _02920_;
	wire _02921_;
	wire _02922_;
	wire _02923_;
	wire _02924_;
	wire _02925_;
	wire _02926_;
	wire _02927_;
	wire _02928_;
	wire _02929_;
	wire _02930_;
	wire _02931_;
	wire _02932_;
	wire _02933_;
	wire _02934_;
	wire _02935_;
	wire _02936_;
	wire _02937_;
	wire _02938_;
	wire _02939_;
	wire _02940_;
	wire _02941_;
	wire _02942_;
	wire _02943_;
	wire _02944_;
	wire _02945_;
	wire _02946_;
	wire _02947_;
	wire _02948_;
	wire _02949_;
	wire _02950_;
	wire _02951_;
	wire _02952_;
	wire _02953_;
	wire _02954_;
	wire _02955_;
	wire _02956_;
	wire _02957_;
	wire _02958_;
	wire _02959_;
	wire _02960_;
	wire _02961_;
	wire _02962_;
	wire _02963_;
	wire _02964_;
	wire _02965_;
	wire _02966_;
	wire _02967_;
	wire _02968_;
	wire _02969_;
	wire _02970_;
	wire _02971_;
	wire _02972_;
	wire _02973_;
	wire _02974_;
	wire _02975_;
	wire _02976_;
	wire _02977_;
	wire _02978_;
	wire _02979_;
	wire _02980_;
	wire _02981_;
	wire _02982_;
	wire _02983_;
	wire _02984_;
	wire _02985_;
	wire _02986_;
	wire _02987_;
	wire _02988_;
	wire _02989_;
	wire _02990_;
	wire _02991_;
	wire _02992_;
	wire _02993_;
	wire _02994_;
	wire _02995_;
	wire _02996_;
	wire _02997_;
	wire _02998_;
	wire _02999_;
	wire _03000_;
	wire _03001_;
	wire _03002_;
	wire _03003_;
	wire _03004_;
	wire _03005_;
	wire _03006_;
	wire _03007_;
	wire _03008_;
	wire _03009_;
	wire _03010_;
	wire _03011_;
	wire _03012_;
	wire _03013_;
	wire _03014_;
	wire _03015_;
	wire _03016_;
	wire _03017_;
	wire _03018_;
	wire _03019_;
	wire _03020_;
	wire _03021_;
	wire _03022_;
	wire _03023_;
	wire _03024_;
	wire _03025_;
	wire _03026_;
	wire _03027_;
	wire _03028_;
	wire _03029_;
	wire _03030_;
	wire _03031_;
	wire _03032_;
	wire _03033_;
	wire _03034_;
	wire _03035_;
	wire _03036_;
	wire _03037_;
	wire _03038_;
	wire _03039_;
	wire _03040_;
	wire _03041_;
	wire _03042_;
	wire _03043_;
	wire _03044_;
	wire _03045_;
	wire _03046_;
	wire _03047_;
	wire _03048_;
	wire _03049_;
	wire _03050_;
	wire _03051_;
	wire _03052_;
	wire _03053_;
	wire _03054_;
	wire _03055_;
	wire _03056_;
	wire _03057_;
	wire _03058_;
	wire _03059_;
	wire _03060_;
	wire _03061_;
	wire _03062_;
	wire _03063_;
	wire _03064_;
	wire _03065_;
	wire _03066_;
	wire _03067_;
	wire _03068_;
	wire _03069_;
	wire _03070_;
	wire _03071_;
	wire _03072_;
	wire _03073_;
	wire _03074_;
	wire _03075_;
	wire _03076_;
	wire _03077_;
	wire _03078_;
	wire _03079_;
	wire _03080_;
	wire _03081_;
	wire _03082_;
	wire _03083_;
	wire _03084_;
	wire _03085_;
	wire _03086_;
	wire _03087_;
	wire _03088_;
	wire _03089_;
	wire _03090_;
	wire _03091_;
	wire _03092_;
	wire _03093_;
	wire _03094_;
	wire _03095_;
	wire _03096_;
	wire _03097_;
	wire _03098_;
	wire _03099_;
	wire _03100_;
	wire _03101_;
	wire _03102_;
	wire _03103_;
	wire _03104_;
	wire _03105_;
	wire _03106_;
	wire _03107_;
	wire _03108_;
	wire _03109_;
	wire _03110_;
	wire _03111_;
	wire _03112_;
	wire _03113_;
	wire _03114_;
	wire _03115_;
	wire _03116_;
	wire _03117_;
	wire _03118_;
	wire _03119_;
	wire _03120_;
	wire _03121_;
	wire _03122_;
	wire _03123_;
	wire _03124_;
	wire _03125_;
	wire _03126_;
	wire _03127_;
	wire _03128_;
	wire _03129_;
	wire _03130_;
	wire _03131_;
	wire _03132_;
	wire _03133_;
	wire _03134_;
	wire _03135_;
	wire _03136_;
	wire _03137_;
	wire _03138_;
	wire _03139_;
	wire _03140_;
	wire _03141_;
	wire _03142_;
	wire _03143_;
	wire _03144_;
	wire _03145_;
	wire _03146_;
	wire _03147_;
	wire _03148_;
	wire _03149_;
	wire _03150_;
	wire _03151_;
	wire _03152_;
	wire _03153_;
	wire _03154_;
	wire _03155_;
	wire _03156_;
	wire _03157_;
	wire _03158_;
	wire _03159_;
	wire _03160_;
	wire _03161_;
	wire _03162_;
	wire _03163_;
	wire _03164_;
	wire _03165_;
	wire _03166_;
	wire _03167_;
	wire _03168_;
	wire _03169_;
	wire _03170_;
	wire _03171_;
	wire _03172_;
	wire _03173_;
	wire _03174_;
	wire _03175_;
	wire _03176_;
	wire _03177_;
	wire _03178_;
	wire _03179_;
	wire _03180_;
	wire _03181_;
	wire _03182_;
	wire _03183_;
	wire _03184_;
	wire _03185_;
	wire _03186_;
	wire _03187_;
	wire _03188_;
	wire _03189_;
	wire _03190_;
	wire _03191_;
	wire _03192_;
	wire _03193_;
	wire _03194_;
	wire _03195_;
	wire _03196_;
	wire _03197_;
	wire _03198_;
	wire _03199_;
	wire _03200_;
	wire _03201_;
	wire _03202_;
	wire _03203_;
	wire _03204_;
	wire _03205_;
	wire _03206_;
	wire _03207_;
	wire _03208_;
	wire _03209_;
	wire _03210_;
	wire _03211_;
	wire _03212_;
	wire _03213_;
	wire _03214_;
	wire _03215_;
	wire _03216_;
	wire _03217_;
	wire _03218_;
	wire _03219_;
	wire _03220_;
	wire _03221_;
	wire _03222_;
	wire _03223_;
	wire _03224_;
	wire _03225_;
	wire _03226_;
	wire _03227_;
	wire _03228_;
	wire _03229_;
	wire _03230_;
	wire _03231_;
	wire _03232_;
	wire _03233_;
	wire _03234_;
	wire _03235_;
	wire _03236_;
	wire _03237_;
	wire _03238_;
	wire _03239_;
	wire _03240_;
	wire _03241_;
	wire _03242_;
	wire _03243_;
	wire _03244_;
	wire _03245_;
	wire _03246_;
	wire _03247_;
	wire _03248_;
	wire _03249_;
	wire _03250_;
	wire _03251_;
	wire _03252_;
	wire _03253_;
	wire _03254_;
	wire _03255_;
	wire _03256_;
	wire _03257_;
	wire _03258_;
	wire _03259_;
	wire _03260_;
	wire _03261_;
	wire _03262_;
	wire _03263_;
	wire _03264_;
	wire _03265_;
	wire _03266_;
	wire _03267_;
	wire _03268_;
	wire _03269_;
	wire _03270_;
	wire _03271_;
	wire _03272_;
	wire _03273_;
	wire _03274_;
	wire _03275_;
	wire _03276_;
	wire _03277_;
	wire _03278_;
	wire _03279_;
	wire _03280_;
	wire _03281_;
	wire _03282_;
	wire _03283_;
	wire _03284_;
	wire _03285_;
	wire _03286_;
	wire _03287_;
	wire _03288_;
	wire _03289_;
	wire _03290_;
	wire _03291_;
	wire _03292_;
	wire _03293_;
	wire _03294_;
	wire _03295_;
	wire _03296_;
	wire _03297_;
	wire _03298_;
	wire _03299_;
	wire _03300_;
	wire _03301_;
	wire _03302_;
	wire _03303_;
	wire _03304_;
	wire _03305_;
	wire _03306_;
	wire _03307_;
	wire _03308_;
	wire _03309_;
	wire _03310_;
	wire _03311_;
	wire _03312_;
	wire _03313_;
	wire _03314_;
	wire _03315_;
	wire _03316_;
	wire _03317_;
	wire _03318_;
	wire _03319_;
	wire _03320_;
	wire _03321_;
	wire _03322_;
	wire _03323_;
	wire _03324_;
	wire _03325_;
	wire _03326_;
	wire _03327_;
	wire _03328_;
	wire _03329_;
	wire _03330_;
	wire _03331_;
	wire _03332_;
	wire _03333_;
	wire _03334_;
	wire _03335_;
	wire _03336_;
	wire _03337_;
	wire _03338_;
	wire _03339_;
	wire _03340_;
	wire _03341_;
	wire _03342_;
	wire _03343_;
	wire _03344_;
	wire _03345_;
	wire _03346_;
	wire _03347_;
	wire _03348_;
	wire _03349_;
	wire _03350_;
	wire _03351_;
	wire _03352_;
	wire _03353_;
	wire _03354_;
	wire _03355_;
	wire _03356_;
	wire _03357_;
	wire _03358_;
	wire _03359_;
	wire _03360_;
	wire _03361_;
	wire _03362_;
	wire _03363_;
	wire _03364_;
	wire _03365_;
	wire _03366_;
	wire _03367_;
	wire _03368_;
	wire _03369_;
	wire _03370_;
	wire _03371_;
	wire _03372_;
	wire _03373_;
	wire _03374_;
	wire _03375_;
	wire _03376_;
	wire _03377_;
	wire _03378_;
	wire _03379_;
	wire _03380_;
	wire _03381_;
	wire _03382_;
	wire _03383_;
	wire _03384_;
	wire _03385_;
	wire _03386_;
	wire _03387_;
	wire _03388_;
	wire _03389_;
	wire _03390_;
	wire _03391_;
	wire _03392_;
	wire _03393_;
	wire _03394_;
	wire _03395_;
	wire _03396_;
	wire _03397_;
	wire _03398_;
	wire _03399_;
	wire _03400_;
	wire _03401_;
	wire _03402_;
	wire _03403_;
	wire _03404_;
	wire _03405_;
	wire _03406_;
	wire _03407_;
	wire _03408_;
	wire _03409_;
	wire _03410_;
	wire _03411_;
	wire _03412_;
	wire _03413_;
	wire _03414_;
	wire _03415_;
	wire _03416_;
	wire _03417_;
	wire _03418_;
	wire _03419_;
	wire _03420_;
	wire _03421_;
	wire _03422_;
	wire _03423_;
	wire _03424_;
	wire _03425_;
	wire _03426_;
	wire _03427_;
	wire _03428_;
	wire _03429_;
	wire _03430_;
	wire _03431_;
	wire _03432_;
	wire _03433_;
	wire _03434_;
	wire _03435_;
	wire _03436_;
	wire _03437_;
	wire _03438_;
	wire _03439_;
	wire _03440_;
	wire _03441_;
	wire _03442_;
	wire _03443_;
	wire _03444_;
	wire _03445_;
	wire _03446_;
	wire _03447_;
	wire _03448_;
	wire _03449_;
	wire _03450_;
	wire _03451_;
	wire _03452_;
	wire _03453_;
	wire _03454_;
	wire _03455_;
	wire _03456_;
	wire _03457_;
	wire _03458_;
	wire _03459_;
	wire _03460_;
	wire _03461_;
	wire _03462_;
	wire _03463_;
	wire _03464_;
	wire _03465_;
	wire _03466_;
	wire _03467_;
	wire _03468_;
	wire _03469_;
	wire _03470_;
	wire _03471_;
	wire _03472_;
	wire _03473_;
	wire _03474_;
	wire _03475_;
	wire _03476_;
	wire _03477_;
	wire _03478_;
	wire _03479_;
	wire _03480_;
	wire _03481_;
	wire _03482_;
	wire _03483_;
	wire _03484_;
	wire _03485_;
	wire _03486_;
	wire _03487_;
	wire _03488_;
	wire _03489_;
	wire _03490_;
	wire _03491_;
	wire _03492_;
	wire _03493_;
	wire _03494_;
	wire _03495_;
	wire _03496_;
	wire _03497_;
	wire _03498_;
	wire _03499_;
	wire _03500_;
	wire _03501_;
	wire _03502_;
	wire _03503_;
	wire _03504_;
	wire _03505_;
	wire _03506_;
	wire _03507_;
	wire _03508_;
	wire _03509_;
	wire _03510_;
	wire _03511_;
	wire _03512_;
	wire _03513_;
	wire _03514_;
	wire _03515_;
	wire _03516_;
	wire _03517_;
	wire _03518_;
	wire _03519_;
	wire _03520_;
	wire _03521_;
	wire _03522_;
	wire _03523_;
	wire _03524_;
	wire _03525_;
	wire _03526_;
	wire _03527_;
	wire _03528_;
	wire _03529_;
	wire _03530_;
	wire _03531_;
	wire _03532_;
	wire _03533_;
	wire _03534_;
	wire _03535_;
	wire _03536_;
	wire _03537_;
	wire _03538_;
	wire _03539_;
	wire _03540_;
	wire _03541_;
	wire _03542_;
	wire _03543_;
	wire _03544_;
	wire _03545_;
	wire _03546_;
	wire _03547_;
	wire _03548_;
	wire _03549_;
	wire _03550_;
	wire _03551_;
	wire _03552_;
	wire _03553_;
	wire _03554_;
	wire _03555_;
	wire _03556_;
	wire _03557_;
	wire _03558_;
	wire _03559_;
	wire _03560_;
	wire _03561_;
	wire _03562_;
	wire _03563_;
	wire _03564_;
	wire _03565_;
	wire _03566_;
	wire _03567_;
	wire _03568_;
	wire _03569_;
	wire _03570_;
	wire _03571_;
	wire _03572_;
	wire _03573_;
	wire _03574_;
	wire _03575_;
	wire _03576_;
	wire _03577_;
	wire _03578_;
	wire _03579_;
	wire _03580_;
	wire _03581_;
	wire _03582_;
	wire _03583_;
	wire _03584_;
	wire _03585_;
	wire _03586_;
	wire _03587_;
	wire _03588_;
	wire _03589_;
	wire _03590_;
	wire _03591_;
	wire _03592_;
	wire _03593_;
	wire _03594_;
	wire _03595_;
	wire _03596_;
	wire _03597_;
	wire _03598_;
	wire _03599_;
	wire _03600_;
	wire _03601_;
	wire _03602_;
	wire _03603_;
	wire _03604_;
	wire _03605_;
	wire _03606_;
	wire _03607_;
	wire _03608_;
	wire _03609_;
	wire _03610_;
	wire _03611_;
	wire _03612_;
	wire _03613_;
	wire _03614_;
	wire _03615_;
	wire _03616_;
	wire _03617_;
	wire _03618_;
	wire _03619_;
	wire _03620_;
	wire _03621_;
	wire _03622_;
	wire _03623_;
	wire _03624_;
	wire _03625_;
	wire _03626_;
	wire _03627_;
	wire _03628_;
	wire _03629_;
	wire _03630_;
	wire _03631_;
	wire _03632_;
	wire _03633_;
	wire _03634_;
	wire _03635_;
	wire _03636_;
	wire _03637_;
	wire _03638_;
	wire _03639_;
	wire _03640_;
	wire _03641_;
	wire _03642_;
	wire _03643_;
	wire _03644_;
	wire _03645_;
	wire _03646_;
	wire _03647_;
	wire _03648_;
	wire _03649_;
	wire _03650_;
	wire _03651_;
	wire _03652_;
	wire _03653_;
	wire _03654_;
	wire _03655_;
	wire _03656_;
	wire _03657_;
	wire _03658_;
	wire _03659_;
	wire _03660_;
	wire _03661_;
	wire _03662_;
	wire _03663_;
	wire _03664_;
	wire _03665_;
	wire _03666_;
	wire _03667_;
	wire _03668_;
	wire _03669_;
	wire _03670_;
	wire _03671_;
	wire _03672_;
	wire _03673_;
	wire _03674_;
	wire _03675_;
	wire _03676_;
	wire _03677_;
	wire _03678_;
	wire _03679_;
	wire _03680_;
	wire _03681_;
	wire _03682_;
	wire _03683_;
	wire _03684_;
	wire _03685_;
	wire _03686_;
	wire _03687_;
	wire _03688_;
	wire _03689_;
	wire _03690_;
	wire _03691_;
	wire _03692_;
	wire _03693_;
	wire _03694_;
	wire _03695_;
	wire _03696_;
	wire _03697_;
	wire _03698_;
	wire _03699_;
	wire _03700_;
	wire _03701_;
	wire _03702_;
	wire _03703_;
	wire _03704_;
	wire _03705_;
	wire _03706_;
	wire _03707_;
	wire _03708_;
	wire _03709_;
	wire _03710_;
	wire _03711_;
	wire _03712_;
	wire _03713_;
	wire _03714_;
	wire _03715_;
	wire _03716_;
	wire _03717_;
	wire _03718_;
	wire _03719_;
	wire _03720_;
	wire _03721_;
	wire _03722_;
	wire _03723_;
	wire _03724_;
	wire _03725_;
	wire _03726_;
	wire _03727_;
	wire _03728_;
	wire _03729_;
	wire _03730_;
	wire _03731_;
	wire _03732_;
	wire _03733_;
	wire _03734_;
	wire _03735_;
	wire _03736_;
	wire _03737_;
	wire _03738_;
	wire _03739_;
	wire _03740_;
	wire _03741_;
	wire _03742_;
	wire _03743_;
	wire _03744_;
	wire _03745_;
	wire _03746_;
	wire _03747_;
	wire _03748_;
	wire _03749_;
	wire _03750_;
	wire _03751_;
	wire _03752_;
	wire _03753_;
	wire _03754_;
	wire _03755_;
	wire _03756_;
	wire _03757_;
	wire _03758_;
	wire _03759_;
	wire _03760_;
	wire _03761_;
	wire _03762_;
	wire _03763_;
	wire _03764_;
	wire _03765_;
	wire _03766_;
	wire _03767_;
	wire _03768_;
	wire _03769_;
	wire _03770_;
	wire _03771_;
	wire _03772_;
	wire _03773_;
	wire _03774_;
	wire _03775_;
	wire _03776_;
	wire _03777_;
	wire _03778_;
	wire _03779_;
	wire _03780_;
	wire _03781_;
	wire _03782_;
	wire _03783_;
	wire _03784_;
	wire _03785_;
	wire _03786_;
	wire _03787_;
	wire _03788_;
	wire _03789_;
	wire _03790_;
	wire _03791_;
	wire _03792_;
	wire _03793_;
	wire _03794_;
	wire _03795_;
	wire _03796_;
	wire _03797_;
	wire _03798_;
	wire _03799_;
	wire _03800_;
	wire _03801_;
	wire _03802_;
	wire _03803_;
	wire _03804_;
	wire _03805_;
	wire _03806_;
	wire _03807_;
	wire _03808_;
	wire _03809_;
	wire _03810_;
	wire _03811_;
	wire _03812_;
	wire _03813_;
	wire _03814_;
	wire _03815_;
	wire _03816_;
	wire _03817_;
	wire _03818_;
	wire _03819_;
	wire _03820_;
	wire _03821_;
	wire _03822_;
	wire _03823_;
	wire _03824_;
	wire _03825_;
	wire _03826_;
	wire _03827_;
	wire _03828_;
	wire _03829_;
	wire _03830_;
	wire _03831_;
	wire _03832_;
	wire _03833_;
	wire _03834_;
	wire _03835_;
	wire _03836_;
	wire _03837_;
	wire _03838_;
	wire _03839_;
	wire _03840_;
	wire _03841_;
	wire _03842_;
	wire _03843_;
	wire _03844_;
	wire _03845_;
	wire _03846_;
	wire _03847_;
	wire _03848_;
	wire _03849_;
	wire _03850_;
	wire _03851_;
	wire _03852_;
	wire _03853_;
	wire _03854_;
	wire _03855_;
	wire _03856_;
	wire _03857_;
	wire _03858_;
	wire _03859_;
	wire _03860_;
	wire _03861_;
	wire _03862_;
	wire _03863_;
	wire _03864_;
	wire _03865_;
	wire _03866_;
	wire _03867_;
	wire _03868_;
	wire _03869_;
	wire _03870_;
	wire _03871_;
	wire _03872_;
	wire _03873_;
	wire _03874_;
	wire _03875_;
	wire _03876_;
	wire _03877_;
	wire _03878_;
	wire _03879_;
	wire _03880_;
	wire _03881_;
	wire _03882_;
	wire _03883_;
	wire _03884_;
	wire _03885_;
	wire _03886_;
	wire _03887_;
	wire _03888_;
	wire _03889_;
	wire _03890_;
	wire _03891_;
	wire _03892_;
	wire _03893_;
	wire _03894_;
	wire _03895_;
	wire _03896_;
	wire _03897_;
	wire _03898_;
	wire _03899_;
	wire _03900_;
	wire _03901_;
	wire _03902_;
	wire _03903_;
	wire _03904_;
	wire _03905_;
	wire _03906_;
	wire _03907_;
	wire _03908_;
	wire _03909_;
	wire _03910_;
	wire _03911_;
	wire _03912_;
	wire _03913_;
	wire _03914_;
	wire _03915_;
	wire _03916_;
	wire _03917_;
	wire _03918_;
	wire _03919_;
	wire _03920_;
	wire _03921_;
	wire _03922_;
	wire _03923_;
	wire _03924_;
	wire _03925_;
	wire _03926_;
	wire _03927_;
	wire _03928_;
	wire _03929_;
	wire _03930_;
	wire _03931_;
	wire _03932_;
	wire _03933_;
	wire _03934_;
	wire _03935_;
	wire _03936_;
	wire _03937_;
	wire _03938_;
	wire _03939_;
	wire _03940_;
	wire _03941_;
	wire _03942_;
	wire _03943_;
	wire _03944_;
	wire _03945_;
	wire _03946_;
	wire _03947_;
	wire _03948_;
	wire _03949_;
	wire _03950_;
	wire _03951_;
	wire _03952_;
	wire _03953_;
	wire _03954_;
	wire _03955_;
	wire _03956_;
	wire _03957_;
	wire _03958_;
	wire _03959_;
	wire _03960_;
	wire _03961_;
	wire _03962_;
	wire _03963_;
	wire _03964_;
	wire _03965_;
	wire _03966_;
	wire _03967_;
	wire _03968_;
	wire _03969_;
	wire _03970_;
	wire _03971_;
	wire _03972_;
	wire _03973_;
	wire _03974_;
	wire _03975_;
	wire _03976_;
	wire _03977_;
	wire _03978_;
	wire _03979_;
	wire _03980_;
	wire _03981_;
	wire _03982_;
	wire _03983_;
	wire _03984_;
	wire _03985_;
	wire _03986_;
	wire _03987_;
	wire _03988_;
	wire _03989_;
	wire _03990_;
	wire _03991_;
	wire _03992_;
	wire _03993_;
	wire _03994_;
	wire _03995_;
	wire _03996_;
	wire _03997_;
	wire _03998_;
	wire _03999_;
	wire _04000_;
	wire _04001_;
	wire _04002_;
	wire _04003_;
	wire _04004_;
	wire _04005_;
	wire _04006_;
	wire _04007_;
	wire _04008_;
	wire _04009_;
	wire _04010_;
	wire _04011_;
	wire _04012_;
	wire _04013_;
	wire _04014_;
	wire _04015_;
	wire _04016_;
	wire _04017_;
	wire _04018_;
	wire _04019_;
	wire _04020_;
	wire _04021_;
	wire _04022_;
	wire _04023_;
	wire _04024_;
	wire _04025_;
	wire _04026_;
	wire _04027_;
	wire _04028_;
	wire _04029_;
	wire _04030_;
	wire _04031_;
	wire _04032_;
	wire _04033_;
	wire _04034_;
	wire _04035_;
	wire _04036_;
	wire _04037_;
	wire _04038_;
	wire _04039_;
	wire _04040_;
	wire _04041_;
	wire _04042_;
	wire _04043_;
	wire _04044_;
	wire _04045_;
	wire _04046_;
	wire _04047_;
	wire _04048_;
	wire _04049_;
	wire _04050_;
	wire _04051_;
	wire _04052_;
	wire _04053_;
	wire _04054_;
	wire _04055_;
	wire _04056_;
	wire _04057_;
	wire _04058_;
	wire _04059_;
	wire _04060_;
	wire _04061_;
	wire _04062_;
	wire _04063_;
	wire _04064_;
	wire _04065_;
	wire _04066_;
	wire _04067_;
	wire _04068_;
	wire _04069_;
	wire _04070_;
	wire _04071_;
	wire _04072_;
	wire _04073_;
	wire _04074_;
	wire _04075_;
	wire _04076_;
	wire _04077_;
	wire _04078_;
	wire _04079_;
	wire _04080_;
	wire _04081_;
	wire _04082_;
	wire _04083_;
	wire _04084_;
	wire _04085_;
	wire _04086_;
	wire _04087_;
	wire _04088_;
	wire _04089_;
	wire _04090_;
	wire _04091_;
	wire _04092_;
	wire _04093_;
	wire _04094_;
	wire _04095_;
	wire _04096_;
	wire _04097_;
	wire _04098_;
	wire _04099_;
	wire _04100_;
	wire _04101_;
	wire _04102_;
	wire _04103_;
	wire _04104_;
	wire _04105_;
	wire _04106_;
	wire _04107_;
	wire _04108_;
	wire _04109_;
	wire _04110_;
	wire _04111_;
	wire _04112_;
	wire _04113_;
	wire _04114_;
	wire _04115_;
	wire _04116_;
	wire _04117_;
	wire _04118_;
	wire _04119_;
	wire _04120_;
	wire _04121_;
	wire _04122_;
	wire _04123_;
	wire _04124_;
	wire _04125_;
	wire _04126_;
	wire _04127_;
	wire _04128_;
	wire _04129_;
	wire _04130_;
	wire _04131_;
	wire _04132_;
	wire _04133_;
	wire _04134_;
	wire _04135_;
	wire _04136_;
	wire _04137_;
	wire _04138_;
	wire _04139_;
	wire _04140_;
	wire _04141_;
	wire _04142_;
	wire _04143_;
	wire _04144_;
	wire _04145_;
	wire _04146_;
	wire _04147_;
	wire _04148_;
	wire _04149_;
	wire _04150_;
	wire _04151_;
	wire _04152_;
	wire _04153_;
	wire _04154_;
	wire _04155_;
	wire _04156_;
	wire _04157_;
	wire _04158_;
	wire _04159_;
	wire _04160_;
	wire _04161_;
	wire _04162_;
	wire _04163_;
	wire _04164_;
	wire _04165_;
	wire _04166_;
	wire _04167_;
	wire _04168_;
	wire _04169_;
	wire _04170_;
	wire _04171_;
	wire _04172_;
	wire _04173_;
	wire _04174_;
	wire _04175_;
	wire _04176_;
	wire _04177_;
	wire _04178_;
	wire _04179_;
	wire _04180_;
	wire _04181_;
	wire _04182_;
	wire _04183_;
	wire _04184_;
	wire _04185_;
	wire _04186_;
	wire _04187_;
	wire _04188_;
	wire _04189_;
	wire _04190_;
	wire _04191_;
	wire _04192_;
	wire _04193_;
	wire _04194_;
	wire _04195_;
	wire _04196_;
	wire _04197_;
	wire _04198_;
	wire _04199_;
	wire _04200_;
	wire _04201_;
	wire _04202_;
	wire _04203_;
	wire _04204_;
	wire _04205_;
	wire _04206_;
	wire _04207_;
	wire _04208_;
	wire _04209_;
	wire _04210_;
	wire _04211_;
	wire _04212_;
	wire _04213_;
	wire _04214_;
	wire _04215_;
	wire _04216_;
	wire _04217_;
	wire _04218_;
	wire _04219_;
	wire _04220_;
	wire _04221_;
	wire _04222_;
	wire _04223_;
	wire _04224_;
	wire _04225_;
	wire _04226_;
	wire _04227_;
	wire _04228_;
	wire _04229_;
	wire _04230_;
	wire _04231_;
	wire _04232_;
	wire _04233_;
	wire _04234_;
	wire _04235_;
	wire _04236_;
	wire _04237_;
	wire _04238_;
	wire _04239_;
	wire _04240_;
	wire _04241_;
	wire _04242_;
	wire _04243_;
	wire _04244_;
	wire _04245_;
	wire _04246_;
	wire _04247_;
	wire _04248_;
	wire _04249_;
	wire _04250_;
	wire _04251_;
	wire _04252_;
	wire _04253_;
	wire _04254_;
	wire _04255_;
	wire _04256_;
	wire _04257_;
	wire _04258_;
	wire _04259_;
	wire _04260_;
	wire _04261_;
	wire _04262_;
	wire _04263_;
	wire _04264_;
	wire _04265_;
	wire _04266_;
	wire _04267_;
	wire _04268_;
	wire _04269_;
	wire _04270_;
	wire _04271_;
	wire _04272_;
	wire _04273_;
	wire _04274_;
	wire _04275_;
	wire _04276_;
	wire _04277_;
	wire _04278_;
	wire _04279_;
	wire _04280_;
	wire _04281_;
	wire _04282_;
	wire _04283_;
	wire _04284_;
	wire _04285_;
	wire _04286_;
	wire _04287_;
	wire _04288_;
	wire _04289_;
	wire _04290_;
	wire _04291_;
	wire _04292_;
	wire _04293_;
	wire _04294_;
	wire _04295_;
	wire _04296_;
	wire _04297_;
	wire _04298_;
	wire _04299_;
	wire _04300_;
	wire _04301_;
	wire _04302_;
	wire _04303_;
	wire _04304_;
	wire _04305_;
	wire _04306_;
	wire _04307_;
	wire _04308_;
	wire _04309_;
	wire _04310_;
	wire _04311_;
	wire _04312_;
	wire _04313_;
	wire _04314_;
	wire _04315_;
	wire _04316_;
	wire _04317_;
	wire _04318_;
	wire _04319_;
	wire _04320_;
	wire _04321_;
	wire _04322_;
	wire _04323_;
	wire _04324_;
	wire _04325_;
	wire _04326_;
	wire _04327_;
	wire _04328_;
	wire _04329_;
	wire _04330_;
	wire _04331_;
	wire _04332_;
	wire _04333_;
	wire _04334_;
	wire _04335_;
	wire _04336_;
	wire _04337_;
	wire _04338_;
	wire _04339_;
	wire _04340_;
	wire _04341_;
	wire _04342_;
	wire _04343_;
	wire _04344_;
	wire _04345_;
	wire _04346_;
	wire _04347_;
	wire _04348_;
	wire _04349_;
	wire _04350_;
	wire _04351_;
	wire _04352_;
	wire _04353_;
	wire _04354_;
	wire _04355_;
	wire _04356_;
	wire _04357_;
	wire _04358_;
	wire _04359_;
	wire _04360_;
	wire _04361_;
	wire _04362_;
	wire _04363_;
	wire _04364_;
	wire _04365_;
	wire _04366_;
	wire _04367_;
	wire _04368_;
	wire _04369_;
	wire _04370_;
	wire _04371_;
	wire _04372_;
	wire _04373_;
	wire _04374_;
	wire _04375_;
	wire _04376_;
	wire _04377_;
	wire _04378_;
	wire _04379_;
	wire _04380_;
	wire _04381_;
	wire _04382_;
	wire _04383_;
	wire _04384_;
	wire _04385_;
	wire _04386_;
	wire _04387_;
	wire _04388_;
	wire _04389_;
	wire _04390_;
	wire _04391_;
	wire _04392_;
	wire _04393_;
	wire _04394_;
	wire _04395_;
	wire _04396_;
	wire _04397_;
	wire _04398_;
	wire _04399_;
	wire _04400_;
	wire _04401_;
	wire _04402_;
	wire _04403_;
	wire _04404_;
	wire _04405_;
	wire _04406_;
	wire _04407_;
	wire _04408_;
	wire _04409_;
	wire _04410_;
	wire _04411_;
	wire _04412_;
	wire _04413_;
	wire _04414_;
	wire _04415_;
	wire _04416_;
	wire _04417_;
	wire _04418_;
	wire _04419_;
	wire _04420_;
	wire _04421_;
	wire _04422_;
	wire _04423_;
	wire _04424_;
	wire _04425_;
	wire _04426_;
	wire _04427_;
	wire _04428_;
	wire _04429_;
	wire _04430_;
	wire _04431_;
	wire _04432_;
	wire _04433_;
	wire _04434_;
	wire _04435_;
	wire _04436_;
	wire _04437_;
	wire _04438_;
	wire _04439_;
	wire _04440_;
	wire _04441_;
	wire _04442_;
	wire _04443_;
	wire _04444_;
	wire _04445_;
	wire _04446_;
	wire _04447_;
	wire _04448_;
	wire _04449_;
	wire _04450_;
	wire _04451_;
	wire _04452_;
	wire _04453_;
	wire _04454_;
	wire _04455_;
	wire _04456_;
	wire _04457_;
	wire _04458_;
	wire _04459_;
	wire _04460_;
	wire _04461_;
	wire _04462_;
	wire _04463_;
	wire _04464_;
	wire _04465_;
	wire _04466_;
	wire _04467_;
	wire _04468_;
	wire _04469_;
	wire _04470_;
	wire _04471_;
	wire _04472_;
	wire _04473_;
	wire _04474_;
	wire _04475_;
	wire _04476_;
	wire _04477_;
	wire _04478_;
	wire _04479_;
	wire _04480_;
	wire _04481_;
	wire _04482_;
	wire _04483_;
	wire _04484_;
	wire _04485_;
	wire _04486_;
	wire _04487_;
	wire _04488_;
	wire _04489_;
	wire _04490_;
	wire _04491_;
	wire _04492_;
	wire _04493_;
	wire _04494_;
	wire _04495_;
	wire _04496_;
	wire _04497_;
	wire _04498_;
	wire _04499_;
	wire _04500_;
	wire _04501_;
	wire _04502_;
	wire _04503_;
	wire _04504_;
	wire _04505_;
	wire _04506_;
	wire _04507_;
	wire _04508_;
	wire _04509_;
	wire _04510_;
	wire _04511_;
	wire _04512_;
	wire _04513_;
	wire _04514_;
	wire _04515_;
	wire _04516_;
	wire _04517_;
	wire _04518_;
	wire _04519_;
	wire _04520_;
	wire _04521_;
	wire _04522_;
	wire _04523_;
	wire _04524_;
	wire _04525_;
	wire _04526_;
	wire _04527_;
	wire _04528_;
	wire _04529_;
	wire _04530_;
	wire _04531_;
	wire _04532_;
	wire _04533_;
	wire _04534_;
	wire _04535_;
	wire _04536_;
	wire _04537_;
	wire _04538_;
	wire _04539_;
	wire _04540_;
	wire _04541_;
	wire _04542_;
	wire _04543_;
	wire _04544_;
	wire _04545_;
	wire _04546_;
	wire _04547_;
	wire _04548_;
	wire _04549_;
	wire _04550_;
	wire _04551_;
	wire _04552_;
	wire _04553_;
	wire _04554_;
	wire _04555_;
	wire _04556_;
	wire _04557_;
	wire _04558_;
	wire _04559_;
	wire _04560_;
	wire _04561_;
	wire _04562_;
	wire _04563_;
	wire _04564_;
	wire _04565_;
	wire _04566_;
	wire _04567_;
	wire _04568_;
	wire _04569_;
	wire _04570_;
	wire _04571_;
	wire _04572_;
	wire _04573_;
	wire _04574_;
	wire _04575_;
	wire _04576_;
	wire _04577_;
	wire _04578_;
	wire _04579_;
	wire _04580_;
	wire _04581_;
	wire _04582_;
	wire _04583_;
	wire _04584_;
	wire _04585_;
	wire _04586_;
	wire _04587_;
	wire _04588_;
	wire _04589_;
	wire _04590_;
	wire _04591_;
	wire _04592_;
	wire _04593_;
	wire _04594_;
	wire _04595_;
	wire _04596_;
	wire _04597_;
	wire _04598_;
	wire _04599_;
	wire _04600_;
	wire _04601_;
	wire _04602_;
	wire _04603_;
	wire _04604_;
	wire _04605_;
	wire _04606_;
	wire _04607_;
	wire _04608_;
	wire _04609_;
	wire _04610_;
	wire _04611_;
	wire _04612_;
	wire _04613_;
	wire _04614_;
	wire _04615_;
	wire _04616_;
	wire _04617_;
	wire _04618_;
	wire _04619_;
	wire _04620_;
	wire _04621_;
	wire _04622_;
	wire _04623_;
	wire _04624_;
	wire _04625_;
	wire _04626_;
	wire _04627_;
	wire _04628_;
	wire _04629_;
	wire _04630_;
	wire _04631_;
	wire _04632_;
	wire _04633_;
	wire _04634_;
	wire _04635_;
	wire _04636_;
	wire _04637_;
	wire _04638_;
	wire _04639_;
	wire _04640_;
	wire _04641_;
	wire _04642_;
	wire _04643_;
	wire _04644_;
	wire _04645_;
	wire _04646_;
	wire _04647_;
	wire _04648_;
	wire _04649_;
	wire _04650_;
	wire _04651_;
	wire _04652_;
	wire _04653_;
	wire _04654_;
	wire _04655_;
	wire _04656_;
	wire _04657_;
	wire _04658_;
	wire _04659_;
	wire _04660_;
	wire _04661_;
	wire _04662_;
	wire _04663_;
	wire _04664_;
	wire _04665_;
	wire _04666_;
	wire _04667_;
	wire _04668_;
	wire _04669_;
	wire _04670_;
	wire _04671_;
	wire _04672_;
	wire _04673_;
	wire _04674_;
	wire _04675_;
	wire _04676_;
	wire _04677_;
	wire _04678_;
	wire _04679_;
	wire _04680_;
	wire _04681_;
	wire _04682_;
	wire _04683_;
	wire _04684_;
	wire _04685_;
	wire _04686_;
	wire _04687_;
	wire _04688_;
	wire _04689_;
	wire _04690_;
	wire _04691_;
	wire _04692_;
	wire _04693_;
	wire _04694_;
	wire _04695_;
	wire _04696_;
	wire _04697_;
	wire _04698_;
	wire _04699_;
	wire _04700_;
	wire _04701_;
	wire _04702_;
	wire _04703_;
	wire _04704_;
	wire _04705_;
	wire _04706_;
	wire _04707_;
	wire _04708_;
	wire _04709_;
	wire _04710_;
	wire _04711_;
	wire _04712_;
	wire _04713_;
	wire _04714_;
	wire _04715_;
	wire _04716_;
	wire _04717_;
	wire _04718_;
	wire _04719_;
	wire _04720_;
	wire _04721_;
	wire _04722_;
	wire _04723_;
	wire _04724_;
	wire _04725_;
	wire _04726_;
	wire _04727_;
	wire _04728_;
	wire _04729_;
	wire _04730_;
	wire _04731_;
	wire _04732_;
	wire _04733_;
	wire _04734_;
	wire _04735_;
	wire _04736_;
	wire _04737_;
	wire _04738_;
	wire _04739_;
	wire _04740_;
	wire _04741_;
	wire _04742_;
	wire _04743_;
	wire _04744_;
	wire _04745_;
	wire _04746_;
	wire _04747_;
	wire _04748_;
	wire _04749_;
	wire _04750_;
	wire _04751_;
	wire _04752_;
	wire _04753_;
	wire _04754_;
	wire _04755_;
	wire _04756_;
	wire _04757_;
	wire _04758_;
	wire _04759_;
	wire _04760_;
	wire _04761_;
	wire _04762_;
	wire _04763_;
	wire _04764_;
	wire _04765_;
	wire _04766_;
	wire _04767_;
	wire _04768_;
	wire _04769_;
	wire _04770_;
	wire _04771_;
	wire _04772_;
	wire _04773_;
	wire _04774_;
	wire _04775_;
	wire _04776_;
	wire _04777_;
	wire _04778_;
	wire _04779_;
	wire _04780_;
	wire _04781_;
	wire _04782_;
	wire _04783_;
	wire _04784_;
	wire _04785_;
	wire _04786_;
	wire _04787_;
	wire _04788_;
	wire _04789_;
	wire _04790_;
	wire _04791_;
	wire _04792_;
	wire _04793_;
	wire _04794_;
	wire _04795_;
	wire _04796_;
	wire _04797_;
	wire _04798_;
	wire _04799_;
	wire _04800_;
	wire _04801_;
	wire _04802_;
	wire _04803_;
	wire _04804_;
	wire _04805_;
	wire _04806_;
	wire _04807_;
	wire _04808_;
	wire _04809_;
	wire _04810_;
	wire _04811_;
	wire _04812_;
	wire _04813_;
	wire _04814_;
	wire _04815_;
	wire _04816_;
	wire _04817_;
	wire _04818_;
	wire _04819_;
	wire _04820_;
	wire _04821_;
	wire _04822_;
	wire _04823_;
	wire _04824_;
	wire _04825_;
	wire _04826_;
	wire _04827_;
	wire _04828_;
	wire _04829_;
	wire _04830_;
	wire _04831_;
	wire _04832_;
	wire _04833_;
	wire _04834_;
	wire _04835_;
	wire _04836_;
	wire _04837_;
	wire _04838_;
	wire _04839_;
	wire _04840_;
	wire _04841_;
	wire _04842_;
	wire _04843_;
	wire _04844_;
	wire _04845_;
	wire _04846_;
	wire _04847_;
	wire _04848_;
	wire _04849_;
	wire _04850_;
	wire _04851_;
	wire _04852_;
	wire _04853_;
	wire _04854_;
	wire _04855_;
	wire _04856_;
	wire _04857_;
	wire _04858_;
	wire _04859_;
	wire _04860_;
	wire _04861_;
	wire _04862_;
	wire _04863_;
	wire _04864_;
	wire _04865_;
	wire _04866_;
	wire _04867_;
	wire _04868_;
	wire _04869_;
	wire _04870_;
	wire _04871_;
	wire _04872_;
	wire _04873_;
	wire _04874_;
	wire _04875_;
	wire _04876_;
	wire _04877_;
	wire _04878_;
	wire _04879_;
	wire _04880_;
	wire _04881_;
	wire _04882_;
	wire _04883_;
	wire _04884_;
	wire _04885_;
	wire _04886_;
	wire _04887_;
	wire _04888_;
	wire _04889_;
	wire _04890_;
	wire _04891_;
	wire _04892_;
	wire _04893_;
	wire _04894_;
	wire _04895_;
	wire _04896_;
	wire _04897_;
	wire _04898_;
	wire _04899_;
	wire _04900_;
	wire _04901_;
	wire _04902_;
	wire _04903_;
	wire _04904_;
	wire _04905_;
	wire _04906_;
	wire _04907_;
	wire _04908_;
	wire _04909_;
	wire _04910_;
	wire _04911_;
	wire _04912_;
	wire _04913_;
	wire _04914_;
	wire _04915_;
	wire _04916_;
	wire _04917_;
	wire _04918_;
	wire _04919_;
	wire _04920_;
	wire _04921_;
	wire _04922_;
	wire _04923_;
	wire _04924_;
	wire _04925_;
	wire _04926_;
	wire _04927_;
	wire _04928_;
	wire _04929_;
	wire _04930_;
	wire _04931_;
	wire _04932_;
	wire _04933_;
	wire _04934_;
	wire _04935_;
	wire _04936_;
	wire _04937_;
	wire _04938_;
	wire _04939_;
	wire _04940_;
	wire _04941_;
	wire _04942_;
	wire _04943_;
	wire _04944_;
	wire _04945_;
	wire _04946_;
	wire _04947_;
	wire _04948_;
	wire _04949_;
	wire _04950_;
	wire _04951_;
	wire _04952_;
	wire _04953_;
	wire _04954_;
	wire _04955_;
	wire _04956_;
	wire _04957_;
	wire _04958_;
	wire _04959_;
	wire _04960_;
	wire _04961_;
	wire _04962_;
	wire _04963_;
	wire _04964_;
	wire _04965_;
	wire _04966_;
	wire _04967_;
	wire _04968_;
	wire _04969_;
	wire _04970_;
	wire _04971_;
	wire _04972_;
	wire _04973_;
	wire _04974_;
	wire _04975_;
	wire _04976_;
	wire _04977_;
	wire _04978_;
	wire _04979_;
	wire _04980_;
	wire _04981_;
	wire _04982_;
	wire _04983_;
	wire _04984_;
	wire _04985_;
	wire _04986_;
	wire _04987_;
	wire _04988_;
	wire _04989_;
	wire _04990_;
	wire _04991_;
	wire _04992_;
	wire _04993_;
	wire _04994_;
	wire _04995_;
	wire _04996_;
	wire _04997_;
	wire _04998_;
	wire _04999_;
	wire _05000_;
	wire _05001_;
	wire _05002_;
	wire _05003_;
	wire _05004_;
	wire _05005_;
	wire _05006_;
	wire _05007_;
	wire _05008_;
	wire _05009_;
	wire _05010_;
	wire _05011_;
	wire _05012_;
	wire _05013_;
	wire _05014_;
	wire _05015_;
	wire _05016_;
	wire _05017_;
	wire _05018_;
	wire _05019_;
	wire _05020_;
	wire _05021_;
	wire _05022_;
	wire _05023_;
	wire _05024_;
	wire _05025_;
	wire _05026_;
	wire _05027_;
	wire _05028_;
	wire _05029_;
	wire _05030_;
	wire _05031_;
	wire _05032_;
	wire _05033_;
	wire _05034_;
	wire _05035_;
	wire _05036_;
	wire _05037_;
	wire _05038_;
	wire _05039_;
	wire _05040_;
	wire _05041_;
	wire _05042_;
	wire _05043_;
	wire _05044_;
	wire _05045_;
	wire _05046_;
	wire _05047_;
	wire _05048_;
	wire _05049_;
	wire _05050_;
	wire _05051_;
	wire _05052_;
	wire _05053_;
	wire _05054_;
	wire _05055_;
	wire _05056_;
	wire _05057_;
	wire _05058_;
	wire _05059_;
	wire _05060_;
	wire _05061_;
	wire _05062_;
	wire _05063_;
	wire _05064_;
	wire _05065_;
	wire _05066_;
	wire _05067_;
	wire _05068_;
	wire _05069_;
	wire _05070_;
	wire _05071_;
	wire _05072_;
	wire _05073_;
	wire _05074_;
	wire _05075_;
	wire _05076_;
	wire _05077_;
	wire _05078_;
	wire _05079_;
	wire _05080_;
	wire _05081_;
	wire _05082_;
	wire _05083_;
	wire _05084_;
	wire _05085_;
	wire _05086_;
	wire _05087_;
	wire _05088_;
	wire _05089_;
	wire _05090_;
	wire _05091_;
	wire _05092_;
	wire _05093_;
	wire _05094_;
	wire _05095_;
	wire _05096_;
	wire _05097_;
	wire _05098_;
	wire _05099_;
	wire _05100_;
	wire _05101_;
	wire _05102_;
	wire _05103_;
	wire _05104_;
	wire _05105_;
	wire _05106_;
	wire _05107_;
	wire _05108_;
	wire _05109_;
	wire _05110_;
	wire _05111_;
	wire _05112_;
	wire _05113_;
	wire _05114_;
	wire _05115_;
	wire _05116_;
	wire _05117_;
	wire _05118_;
	wire _05119_;
	wire _05120_;
	wire _05121_;
	wire _05122_;
	wire _05123_;
	wire _05124_;
	wire _05125_;
	wire _05126_;
	wire _05127_;
	wire _05128_;
	wire _05129_;
	wire _05130_;
	wire _05131_;
	wire _05132_;
	wire _05133_;
	wire _05134_;
	wire _05135_;
	wire _05136_;
	wire _05137_;
	wire _05138_;
	wire _05139_;
	wire _05140_;
	wire _05141_;
	wire _05142_;
	wire _05143_;
	wire _05144_;
	wire _05145_;
	wire _05146_;
	wire _05147_;
	wire _05148_;
	wire _05149_;
	wire _05150_;
	wire _05151_;
	wire _05152_;
	wire _05153_;
	wire _05154_;
	wire _05155_;
	wire _05156_;
	wire _05157_;
	wire _05158_;
	wire _05159_;
	wire _05160_;
	wire _05161_;
	wire _05162_;
	wire _05163_;
	wire _05164_;
	wire _05165_;
	wire _05166_;
	wire _05167_;
	wire _05168_;
	wire _05169_;
	wire _05170_;
	wire _05171_;
	wire _05172_;
	wire _05173_;
	wire _05174_;
	wire _05175_;
	wire _05176_;
	wire _05177_;
	wire _05178_;
	wire _05179_;
	wire _05180_;
	wire _05181_;
	wire _05182_;
	wire _05183_;
	wire _05184_;
	wire _05185_;
	wire _05186_;
	wire _05187_;
	wire _05188_;
	wire _05189_;
	wire _05190_;
	wire _05191_;
	wire _05192_;
	wire _05193_;
	wire _05194_;
	wire _05195_;
	wire _05196_;
	wire _05197_;
	wire _05198_;
	wire _05199_;
	wire _05200_;
	wire _05201_;
	wire _05202_;
	wire _05203_;
	wire _05204_;
	wire _05205_;
	wire _05206_;
	wire _05207_;
	wire _05208_;
	wire _05209_;
	wire _05210_;
	wire _05211_;
	wire _05212_;
	wire _05213_;
	wire _05214_;
	wire _05215_;
	wire _05216_;
	wire _05217_;
	wire _05218_;
	wire _05219_;
	wire _05220_;
	wire _05221_;
	wire _05222_;
	wire _05223_;
	wire _05224_;
	wire _05225_;
	wire _05226_;
	wire _05227_;
	wire _05228_;
	wire _05229_;
	wire _05230_;
	wire _05231_;
	wire _05232_;
	wire _05233_;
	wire _05234_;
	wire _05235_;
	wire _05236_;
	wire _05237_;
	wire _05238_;
	wire _05239_;
	wire _05240_;
	wire _05241_;
	wire _05242_;
	wire _05243_;
	wire _05244_;
	wire _05245_;
	wire _05246_;
	wire _05247_;
	wire _05248_;
	wire _05249_;
	wire _05250_;
	wire _05251_;
	wire _05252_;
	wire _05253_;
	wire _05254_;
	wire _05255_;
	wire _05256_;
	wire _05257_;
	wire _05258_;
	wire _05259_;
	wire _05260_;
	wire _05261_;
	wire _05262_;
	wire _05263_;
	wire _05264_;
	wire _05265_;
	wire _05266_;
	wire _05267_;
	wire _05268_;
	wire _05269_;
	wire _05270_;
	wire _05271_;
	wire _05272_;
	wire _05273_;
	wire _05274_;
	wire _05275_;
	wire _05276_;
	wire _05277_;
	wire _05278_;
	wire _05279_;
	wire _05280_;
	wire _05281_;
	wire _05282_;
	wire _05283_;
	wire _05284_;
	wire _05285_;
	wire _05286_;
	wire _05287_;
	wire _05288_;
	wire _05289_;
	wire _05290_;
	wire _05291_;
	wire _05292_;
	wire _05293_;
	wire _05294_;
	wire _05295_;
	wire _05296_;
	wire _05297_;
	wire _05298_;
	wire _05299_;
	wire _05300_;
	wire _05301_;
	wire _05302_;
	wire _05303_;
	wire _05304_;
	wire _05305_;
	wire _05306_;
	wire _05307_;
	wire _05308_;
	wire _05309_;
	wire _05310_;
	wire _05311_;
	wire _05312_;
	wire _05313_;
	wire _05314_;
	wire _05315_;
	wire _05316_;
	wire _05317_;
	wire _05318_;
	wire _05319_;
	wire _05320_;
	wire _05321_;
	wire _05322_;
	wire _05323_;
	wire _05324_;
	wire _05325_;
	wire _05326_;
	wire _05327_;
	wire _05328_;
	wire _05329_;
	wire _05330_;
	wire _05331_;
	wire _05332_;
	wire _05333_;
	wire _05334_;
	wire _05335_;
	wire _05336_;
	wire _05337_;
	wire _05338_;
	wire _05339_;
	wire _05340_;
	wire _05341_;
	wire _05342_;
	wire _05343_;
	wire _05344_;
	wire _05345_;
	wire _05346_;
	wire _05347_;
	wire _05348_;
	wire _05349_;
	wire _05350_;
	wire _05351_;
	wire _05352_;
	wire _05353_;
	wire _05354_;
	wire _05355_;
	wire _05356_;
	wire _05357_;
	wire _05358_;
	wire _05359_;
	wire _05360_;
	wire _05361_;
	wire _05362_;
	wire _05363_;
	wire _05364_;
	wire _05365_;
	wire _05366_;
	wire _05367_;
	wire _05368_;
	wire _05369_;
	wire _05370_;
	wire _05371_;
	wire _05372_;
	wire _05373_;
	wire _05374_;
	wire _05375_;
	wire _05376_;
	wire _05377_;
	wire _05378_;
	wire _05379_;
	wire _05380_;
	wire _05381_;
	wire _05382_;
	wire _05383_;
	wire _05384_;
	wire _05385_;
	wire _05386_;
	wire _05387_;
	wire _05388_;
	wire _05389_;
	wire _05390_;
	wire _05391_;
	wire _05392_;
	wire _05393_;
	wire _05394_;
	wire _05395_;
	wire _05396_;
	wire _05397_;
	wire _05398_;
	wire _05399_;
	wire _05400_;
	wire _05401_;
	wire _05402_;
	wire _05403_;
	wire _05404_;
	wire _05405_;
	wire _05406_;
	wire _05407_;
	wire _05408_;
	wire _05409_;
	wire _05410_;
	wire _05411_;
	wire _05412_;
	wire _05413_;
	wire _05414_;
	wire _05415_;
	wire _05416_;
	wire _05417_;
	wire _05418_;
	wire _05419_;
	wire _05420_;
	wire _05421_;
	wire _05422_;
	wire _05423_;
	wire _05424_;
	wire _05425_;
	wire _05426_;
	wire _05427_;
	wire _05428_;
	wire _05429_;
	wire _05430_;
	wire _05431_;
	wire _05432_;
	wire _05433_;
	wire _05434_;
	wire _05435_;
	wire _05436_;
	wire _05437_;
	wire _05438_;
	wire _05439_;
	wire _05440_;
	wire _05441_;
	wire _05442_;
	wire _05443_;
	wire _05444_;
	wire _05445_;
	wire _05446_;
	wire _05447_;
	wire _05448_;
	wire _05449_;
	wire _05450_;
	wire _05451_;
	wire _05452_;
	wire _05453_;
	wire _05454_;
	wire _05455_;
	wire _05456_;
	wire _05457_;
	wire _05458_;
	wire _05459_;
	wire _05460_;
	wire _05461_;
	wire _05462_;
	wire _05463_;
	wire _05464_;
	wire _05465_;
	wire _05466_;
	wire _05467_;
	wire _05468_;
	wire _05469_;
	wire _05470_;
	wire _05471_;
	wire _05472_;
	wire _05473_;
	wire _05474_;
	wire _05475_;
	wire _05476_;
	wire _05477_;
	wire _05478_;
	wire _05479_;
	wire _05480_;
	wire _05481_;
	wire _05482_;
	wire _05483_;
	wire _05484_;
	wire _05485_;
	wire _05486_;
	wire _05487_;
	wire _05488_;
	wire _05489_;
	wire _05490_;
	wire _05491_;
	wire _05492_;
	wire _05493_;
	wire _05494_;
	wire _05495_;
	wire _05496_;
	wire _05497_;
	wire _05498_;
	wire _05499_;
	wire _05500_;
	wire _05501_;
	wire _05502_;
	wire _05503_;
	wire _05504_;
	wire _05505_;
	wire _05506_;
	wire _05507_;
	wire _05508_;
	wire _05509_;
	wire _05510_;
	wire _05511_;
	wire _05512_;
	wire _05513_;
	wire _05514_;
	wire _05515_;
	wire _05516_;
	wire _05517_;
	wire _05518_;
	wire _05519_;
	wire _05520_;
	wire _05521_;
	wire _05522_;
	wire _05523_;
	wire _05524_;
	wire _05525_;
	wire _05526_;
	wire _05527_;
	wire _05528_;
	wire _05529_;
	wire _05530_;
	wire _05531_;
	wire _05532_;
	wire _05533_;
	wire _05534_;
	wire _05535_;
	wire _05536_;
	wire _05537_;
	wire _05538_;
	wire _05539_;
	wire _05540_;
	wire _05541_;
	wire _05542_;
	wire _05543_;
	wire _05544_;
	wire _05545_;
	wire _05546_;
	wire _05547_;
	wire _05548_;
	wire _05549_;
	wire _05550_;
	wire _05551_;
	wire _05552_;
	wire _05553_;
	wire _05554_;
	wire _05555_;
	wire _05556_;
	wire _05557_;
	wire _05558_;
	wire _05559_;
	wire _05560_;
	wire _05561_;
	wire _05562_;
	wire _05563_;
	wire _05564_;
	wire _05565_;
	wire _05566_;
	wire _05567_;
	wire _05568_;
	wire _05569_;
	wire _05570_;
	wire _05571_;
	wire _05572_;
	wire _05573_;
	wire _05574_;
	wire _05575_;
	wire _05576_;
	wire _05577_;
	wire _05578_;
	wire _05579_;
	wire _05580_;
	wire _05581_;
	wire _05582_;
	wire _05583_;
	wire _05584_;
	wire _05585_;
	wire _05586_;
	wire _05587_;
	wire _05588_;
	wire _05589_;
	wire _05590_;
	wire _05591_;
	wire _05592_;
	wire _05593_;
	wire _05594_;
	wire _05595_;
	wire _05596_;
	wire _05597_;
	wire _05598_;
	wire _05599_;
	wire _05600_;
	wire _05601_;
	wire _05602_;
	wire _05603_;
	wire _05604_;
	wire _05605_;
	wire _05606_;
	wire _05607_;
	wire _05608_;
	wire _05609_;
	wire _05610_;
	wire _05611_;
	wire _05612_;
	wire _05613_;
	wire _05614_;
	wire _05615_;
	wire _05616_;
	wire _05617_;
	wire _05618_;
	wire _05619_;
	wire _05620_;
	wire _05621_;
	wire _05622_;
	wire _05623_;
	wire _05624_;
	wire _05625_;
	wire _05626_;
	wire _05627_;
	wire _05628_;
	wire _05629_;
	wire _05630_;
	wire _05631_;
	wire _05632_;
	wire _05633_;
	wire _05634_;
	wire _05635_;
	wire _05636_;
	wire _05637_;
	wire _05638_;
	wire _05639_;
	wire _05640_;
	wire _05641_;
	wire _05642_;
	wire _05643_;
	wire _05644_;
	wire _05645_;
	wire _05646_;
	wire _05647_;
	wire _05648_;
	wire _05649_;
	wire _05650_;
	wire _05651_;
	wire _05652_;
	wire _05653_;
	wire _05654_;
	wire _05655_;
	wire _05656_;
	wire _05657_;
	wire _05658_;
	wire _05659_;
	wire _05660_;
	wire _05661_;
	wire _05662_;
	wire _05663_;
	wire _05664_;
	wire _05665_;
	wire _05666_;
	wire _05667_;
	wire _05668_;
	wire _05669_;
	wire _05670_;
	wire _05671_;
	wire _05672_;
	wire _05673_;
	wire _05674_;
	wire _05675_;
	wire _05676_;
	wire _05677_;
	wire _05678_;
	wire _05679_;
	wire _05680_;
	wire _05681_;
	wire _05682_;
	wire _05683_;
	wire _05684_;
	wire _05685_;
	wire _05686_;
	wire _05687_;
	wire _05688_;
	wire _05689_;
	wire _05690_;
	wire _05691_;
	wire _05692_;
	wire _05693_;
	wire _05694_;
	wire _05695_;
	wire _05696_;
	wire _05697_;
	wire _05698_;
	wire _05699_;
	wire _05700_;
	wire _05701_;
	wire _05702_;
	wire _05703_;
	wire _05704_;
	wire _05705_;
	wire _05706_;
	wire _05707_;
	wire _05708_;
	wire _05709_;
	wire _05710_;
	wire _05711_;
	wire _05712_;
	wire _05713_;
	wire _05714_;
	wire _05715_;
	wire _05716_;
	wire _05717_;
	wire _05718_;
	wire _05719_;
	wire _05720_;
	wire _05721_;
	wire _05722_;
	wire _05723_;
	wire _05724_;
	wire _05725_;
	wire _05726_;
	wire _05727_;
	wire _05728_;
	wire _05729_;
	wire _05730_;
	wire _05731_;
	wire _05732_;
	wire _05733_;
	wire _05734_;
	wire _05735_;
	wire _05736_;
	wire _05737_;
	wire _05738_;
	wire _05739_;
	wire _05740_;
	wire _05741_;
	wire _05742_;
	wire _05743_;
	wire _05744_;
	wire _05745_;
	wire _05746_;
	wire _05747_;
	wire _05748_;
	wire _05749_;
	wire _05750_;
	wire _05751_;
	wire _05752_;
	wire _05753_;
	wire _05754_;
	wire _05755_;
	wire _05756_;
	wire _05757_;
	wire _05758_;
	wire _05759_;
	wire _05760_;
	wire _05761_;
	wire _05762_;
	wire _05763_;
	wire _05764_;
	wire _05765_;
	wire _05766_;
	wire _05767_;
	wire _05768_;
	wire _05769_;
	wire _05770_;
	wire _05771_;
	wire _05772_;
	wire _05773_;
	wire _05774_;
	wire _05775_;
	wire _05776_;
	wire _05777_;
	wire _05778_;
	wire _05779_;
	wire _05780_;
	wire _05781_;
	wire _05782_;
	wire _05783_;
	wire _05784_;
	wire _05785_;
	wire _05786_;
	wire _05787_;
	wire _05788_;
	wire _05789_;
	wire _05790_;
	wire _05791_;
	wire _05792_;
	wire _05793_;
	wire _05794_;
	wire _05795_;
	wire _05796_;
	wire _05797_;
	wire _05798_;
	wire _05799_;
	wire _05800_;
	wire _05801_;
	wire _05802_;
	wire _05803_;
	wire _05804_;
	wire _05805_;
	wire _05806_;
	wire _05807_;
	wire _05808_;
	wire _05809_;
	wire _05810_;
	wire _05811_;
	wire _05812_;
	wire _05813_;
	wire _05814_;
	wire _05815_;
	wire _05816_;
	wire _05817_;
	wire _05818_;
	wire _05819_;
	wire _05820_;
	wire _05821_;
	wire _05822_;
	wire _05823_;
	wire _05824_;
	wire _05825_;
	wire _05826_;
	wire _05827_;
	wire _05828_;
	wire _05829_;
	wire _05830_;
	wire _05831_;
	wire _05832_;
	wire _05833_;
	wire _05834_;
	wire _05835_;
	wire _05836_;
	wire _05837_;
	wire _05838_;
	wire _05839_;
	wire _05840_;
	wire _05841_;
	wire _05842_;
	wire _05843_;
	wire _05844_;
	wire _05845_;
	wire _05846_;
	wire _05847_;
	wire _05848_;
	wire _05849_;
	wire _05850_;
	wire _05851_;
	wire _05852_;
	wire _05853_;
	wire _05854_;
	wire _05855_;
	wire _05856_;
	wire _05857_;
	wire _05858_;
	wire _05859_;
	wire _05860_;
	wire _05861_;
	wire _05862_;
	wire _05863_;
	wire _05864_;
	wire _05865_;
	wire _05866_;
	wire _05867_;
	wire _05868_;
	wire _05869_;
	wire _05870_;
	wire _05871_;
	wire _05872_;
	wire _05873_;
	wire _05874_;
	wire _05875_;
	wire _05876_;
	wire _05877_;
	wire _05878_;
	wire _05879_;
	wire _05880_;
	wire _05881_;
	wire _05882_;
	wire _05883_;
	wire _05884_;
	wire _05885_;
	wire _05886_;
	wire _05887_;
	wire _05888_;
	wire _05889_;
	wire _05890_;
	wire _05891_;
	wire _05892_;
	wire _05893_;
	wire _05894_;
	wire _05895_;
	wire _05896_;
	wire _05897_;
	wire _05898_;
	wire _05899_;
	wire _05900_;
	wire _05901_;
	wire _05902_;
	wire _05903_;
	wire _05904_;
	wire _05905_;
	wire _05906_;
	wire _05907_;
	wire _05908_;
	wire _05909_;
	wire _05910_;
	wire _05911_;
	wire _05912_;
	wire _05913_;
	wire _05914_;
	wire _05915_;
	wire _05916_;
	wire _05917_;
	wire _05918_;
	wire _05919_;
	wire _05920_;
	wire _05921_;
	wire _05922_;
	wire _05923_;
	wire _05924_;
	wire _05925_;
	wire _05926_;
	wire _05927_;
	wire _05928_;
	wire _05929_;
	wire _05930_;
	wire _05931_;
	wire _05932_;
	wire _05933_;
	wire _05934_;
	wire _05935_;
	wire _05936_;
	wire _05937_;
	wire _05938_;
	wire _05939_;
	wire _05940_;
	wire _05941_;
	wire _05942_;
	wire _05943_;
	wire _05944_;
	wire _05945_;
	wire _05946_;
	wire _05947_;
	wire _05948_;
	wire _05949_;
	wire _05950_;
	wire _05951_;
	wire _05952_;
	wire _05953_;
	wire _05954_;
	wire _05955_;
	wire _05956_;
	wire _05957_;
	wire _05958_;
	wire _05959_;
	wire _05960_;
	wire _05961_;
	wire _05962_;
	wire _05963_;
	wire _05964_;
	wire _05965_;
	wire _05966_;
	wire _05967_;
	wire _05968_;
	wire _05969_;
	wire _05970_;
	wire _05971_;
	wire _05972_;
	wire _05973_;
	wire _05974_;
	wire _05975_;
	wire _05976_;
	wire _05977_;
	wire _05978_;
	wire _05979_;
	wire _05980_;
	wire _05981_;
	wire _05982_;
	wire _05983_;
	wire _05984_;
	wire _05985_;
	wire _05986_;
	wire _05987_;
	wire _05988_;
	wire _05989_;
	wire _05990_;
	wire _05991_;
	wire _05992_;
	wire _05993_;
	wire _05994_;
	wire _05995_;
	wire _05996_;
	wire _05997_;
	wire _05998_;
	wire _05999_;
	wire _06000_;
	wire _06001_;
	wire _06002_;
	wire _06003_;
	wire _06004_;
	wire _06005_;
	wire _06006_;
	wire _06007_;
	wire _06008_;
	wire _06009_;
	wire _06010_;
	wire _06011_;
	wire _06012_;
	wire _06013_;
	wire _06014_;
	wire _06015_;
	wire _06016_;
	wire _06017_;
	wire _06018_;
	wire _06019_;
	wire _06020_;
	wire _06021_;
	wire _06022_;
	wire _06023_;
	wire _06024_;
	wire _06025_;
	wire _06026_;
	wire _06027_;
	wire _06028_;
	wire _06029_;
	wire _06030_;
	wire _06031_;
	wire _06032_;
	wire _06033_;
	wire _06034_;
	wire _06035_;
	wire _06036_;
	wire _06037_;
	wire _06038_;
	wire _06039_;
	wire _06040_;
	wire _06041_;
	wire _06042_;
	wire _06043_;
	wire _06044_;
	wire _06045_;
	wire _06046_;
	wire _06047_;
	wire _06048_;
	wire _06049_;
	wire _06050_;
	wire _06051_;
	wire _06052_;
	wire _06053_;
	wire _06054_;
	wire _06055_;
	wire _06056_;
	wire _06057_;
	wire _06058_;
	wire _06059_;
	wire _06060_;
	wire _06061_;
	wire _06062_;
	wire _06063_;
	wire _06064_;
	wire _06065_;
	wire _06066_;
	wire _06067_;
	wire _06068_;
	wire _06069_;
	wire _06070_;
	wire _06071_;
	wire _06072_;
	wire _06073_;
	wire _06074_;
	wire _06075_;
	wire _06076_;
	wire _06077_;
	wire _06078_;
	wire _06079_;
	wire _06080_;
	wire _06081_;
	wire _06082_;
	wire _06083_;
	wire _06084_;
	wire _06085_;
	wire _06086_;
	wire _06087_;
	wire _06088_;
	wire _06089_;
	wire _06090_;
	wire _06091_;
	wire _06092_;
	wire _06093_;
	wire _06094_;
	wire _06095_;
	wire _06096_;
	wire _06097_;
	wire _06098_;
	wire _06099_;
	wire _06100_;
	wire _06101_;
	wire _06102_;
	wire _06103_;
	wire _06104_;
	wire _06105_;
	wire _06106_;
	wire _06107_;
	wire _06108_;
	wire _06109_;
	wire _06110_;
	wire _06111_;
	wire _06112_;
	wire _06113_;
	wire _06114_;
	wire _06115_;
	wire _06116_;
	wire _06117_;
	wire _06118_;
	wire _06119_;
	wire _06120_;
	wire _06121_;
	wire _06122_;
	wire _06123_;
	wire _06124_;
	wire _06125_;
	wire _06126_;
	wire _06127_;
	wire _06128_;
	wire _06129_;
	wire _06130_;
	wire _06131_;
	wire _06132_;
	wire _06133_;
	wire _06134_;
	wire _06135_;
	wire _06136_;
	wire _06137_;
	wire _06138_;
	wire _06139_;
	wire _06140_;
	wire _06141_;
	wire _06142_;
	wire _06143_;
	wire _06144_;
	wire _06145_;
	wire _06146_;
	wire _06147_;
	wire _06148_;
	wire _06149_;
	wire _06150_;
	wire _06151_;
	wire _06152_;
	wire _06153_;
	wire _06154_;
	wire _06155_;
	wire _06156_;
	wire _06157_;
	wire _06158_;
	wire _06159_;
	wire _06160_;
	wire _06161_;
	wire _06162_;
	wire _06163_;
	wire _06164_;
	wire _06165_;
	wire _06166_;
	wire _06167_;
	wire _06168_;
	wire _06169_;
	wire _06170_;
	wire _06171_;
	wire _06172_;
	wire _06173_;
	wire _06174_;
	wire _06175_;
	wire _06176_;
	wire _06177_;
	wire _06178_;
	wire _06179_;
	wire _06180_;
	wire _06181_;
	wire _06182_;
	wire _06183_;
	wire _06184_;
	wire _06185_;
	wire _06186_;
	wire _06187_;
	wire _06188_;
	wire _06189_;
	wire _06190_;
	wire _06191_;
	wire _06192_;
	wire _06193_;
	wire _06194_;
	wire _06195_;
	wire _06196_;
	wire _06197_;
	wire _06198_;
	wire _06199_;
	wire _06200_;
	wire _06201_;
	wire _06202_;
	wire _06203_;
	wire _06204_;
	wire _06205_;
	wire _06206_;
	wire _06207_;
	wire _06208_;
	wire _06209_;
	wire _06210_;
	wire _06211_;
	wire _06212_;
	wire _06213_;
	wire _06214_;
	wire _06215_;
	wire _06216_;
	wire _06217_;
	wire _06218_;
	wire _06219_;
	wire _06220_;
	wire _06221_;
	wire _06222_;
	wire _06223_;
	wire _06224_;
	wire _06225_;
	wire _06226_;
	wire _06227_;
	wire _06228_;
	wire _06229_;
	wire _06230_;
	wire _06231_;
	wire _06232_;
	wire _06233_;
	wire _06234_;
	wire _06235_;
	wire _06236_;
	wire _06237_;
	wire _06238_;
	wire _06239_;
	wire _06240_;
	wire _06241_;
	wire _06242_;
	wire _06243_;
	wire _06244_;
	wire _06245_;
	wire _06246_;
	wire _06247_;
	wire _06248_;
	wire _06249_;
	wire _06250_;
	wire _06251_;
	wire _06252_;
	wire _06253_;
	wire _06254_;
	wire _06255_;
	wire _06256_;
	wire _06257_;
	wire _06258_;
	wire _06259_;
	wire _06260_;
	wire _06261_;
	wire _06262_;
	wire _06263_;
	wire _06264_;
	wire _06265_;
	wire _06266_;
	wire _06267_;
	wire _06268_;
	wire _06269_;
	wire _06270_;
	wire _06271_;
	wire _06272_;
	wire _06273_;
	wire _06274_;
	wire _06275_;
	wire _06276_;
	wire _06277_;
	wire _06278_;
	wire _06279_;
	wire _06280_;
	wire _06281_;
	wire _06282_;
	wire _06283_;
	wire _06284_;
	wire _06285_;
	wire _06286_;
	wire _06287_;
	wire _06288_;
	wire _06289_;
	wire _06290_;
	wire _06291_;
	wire _06292_;
	wire _06293_;
	wire _06294_;
	wire _06295_;
	wire _06296_;
	wire _06297_;
	wire _06298_;
	wire _06299_;
	wire _06300_;
	wire _06301_;
	wire _06302_;
	wire _06303_;
	wire _06304_;
	wire _06305_;
	wire _06306_;
	wire _06307_;
	wire _06308_;
	wire _06309_;
	wire _06310_;
	wire _06311_;
	wire _06312_;
	wire _06313_;
	wire _06314_;
	wire _06315_;
	wire _06316_;
	wire _06317_;
	wire _06318_;
	wire _06319_;
	wire _06320_;
	wire _06321_;
	wire _06322_;
	wire _06323_;
	wire _06324_;
	wire _06325_;
	wire _06326_;
	wire _06327_;
	wire _06328_;
	wire _06329_;
	wire _06330_;
	wire _06331_;
	wire _06332_;
	wire _06333_;
	wire _06334_;
	wire _06335_;
	wire _06336_;
	wire _06337_;
	wire _06338_;
	wire _06339_;
	wire _06340_;
	wire _06341_;
	wire _06342_;
	wire _06343_;
	wire _06344_;
	wire _06345_;
	wire _06346_;
	wire _06347_;
	wire _06348_;
	wire _06349_;
	wire _06350_;
	wire _06351_;
	wire _06352_;
	wire _06353_;
	wire _06354_;
	wire _06355_;
	wire _06356_;
	wire _06357_;
	wire _06358_;
	wire _06359_;
	wire _06360_;
	wire _06361_;
	wire _06362_;
	wire _06363_;
	wire _06364_;
	wire _06365_;
	wire _06366_;
	wire _06367_;
	wire _06368_;
	wire _06369_;
	wire _06370_;
	wire _06371_;
	wire _06372_;
	wire _06373_;
	wire _06374_;
	wire _06375_;
	wire _06376_;
	wire _06377_;
	wire _06378_;
	wire _06379_;
	wire _06380_;
	wire _06381_;
	wire _06382_;
	wire _06383_;
	wire _06384_;
	wire _06385_;
	wire _06386_;
	wire _06387_;
	wire _06388_;
	wire _06389_;
	wire _06390_;
	wire _06391_;
	wire _06392_;
	wire _06393_;
	wire _06394_;
	wire _06395_;
	wire _06396_;
	wire _06397_;
	wire _06398_;
	wire _06399_;
	wire _06400_;
	wire _06401_;
	wire _06402_;
	wire _06403_;
	wire _06404_;
	wire _06405_;
	wire _06406_;
	wire _06407_;
	wire _06408_;
	wire _06409_;
	wire _06410_;
	wire _06411_;
	wire _06412_;
	wire _06413_;
	wire _06414_;
	wire _06415_;
	wire _06416_;
	wire _06417_;
	wire _06418_;
	wire _06419_;
	wire _06420_;
	wire _06421_;
	wire _06422_;
	wire _06423_;
	wire _06424_;
	wire _06425_;
	wire _06426_;
	wire _06427_;
	wire _06428_;
	wire _06429_;
	wire _06430_;
	wire _06431_;
	wire _06432_;
	wire _06433_;
	wire _06434_;
	wire _06435_;
	wire _06436_;
	wire _06437_;
	wire _06438_;
	wire _06439_;
	wire _06440_;
	wire _06441_;
	wire _06442_;
	wire _06443_;
	wire _06444_;
	wire _06445_;
	wire _06446_;
	wire _06447_;
	wire _06448_;
	wire _06449_;
	wire _06450_;
	wire _06451_;
	wire _06452_;
	wire _06453_;
	wire _06454_;
	wire _06455_;
	wire _06456_;
	wire _06457_;
	wire _06458_;
	wire _06459_;
	wire _06460_;
	wire _06461_;
	wire _06462_;
	wire _06463_;
	wire _06464_;
	wire _06465_;
	wire _06466_;
	wire _06467_;
	wire _06468_;
	wire _06469_;
	wire _06470_;
	wire _06471_;
	wire _06472_;
	wire _06473_;
	wire _06474_;
	wire _06475_;
	wire _06476_;
	wire _06477_;
	wire _06478_;
	wire _06479_;
	wire _06480_;
	wire _06481_;
	wire _06482_;
	wire _06483_;
	wire _06484_;
	wire _06485_;
	wire _06486_;
	wire _06487_;
	wire _06488_;
	wire _06489_;
	wire _06490_;
	wire _06491_;
	wire _06492_;
	wire _06493_;
	wire _06494_;
	wire _06495_;
	wire _06496_;
	wire _06497_;
	wire _06498_;
	wire _06499_;
	wire _06500_;
	wire _06501_;
	wire _06502_;
	wire _06503_;
	wire _06504_;
	wire _06505_;
	wire _06506_;
	wire _06507_;
	wire _06508_;
	wire _06509_;
	wire _06510_;
	wire _06511_;
	wire _06512_;
	wire _06513_;
	wire _06514_;
	wire _06515_;
	wire _06516_;
	wire _06517_;
	wire _06518_;
	wire _06519_;
	wire _06520_;
	wire _06521_;
	wire _06522_;
	wire _06523_;
	wire _06524_;
	wire _06525_;
	wire _06526_;
	wire _06527_;
	wire _06528_;
	wire _06529_;
	wire _06530_;
	wire _06531_;
	wire _06532_;
	wire _06533_;
	wire _06534_;
	wire _06535_;
	wire _06536_;
	wire _06537_;
	wire _06538_;
	wire _06539_;
	wire _06540_;
	wire _06541_;
	wire _06542_;
	wire _06543_;
	wire _06544_;
	wire _06545_;
	wire _06546_;
	wire _06547_;
	wire _06548_;
	wire _06549_;
	wire _06550_;
	wire _06551_;
	wire _06552_;
	wire _06553_;
	wire _06554_;
	wire _06555_;
	wire _06556_;
	wire _06557_;
	wire _06558_;
	wire _06559_;
	wire _06560_;
	wire _06561_;
	wire _06562_;
	wire _06563_;
	wire _06564_;
	wire _06565_;
	wire _06566_;
	wire _06567_;
	wire _06568_;
	wire _06569_;
	wire _06570_;
	wire _06571_;
	wire _06572_;
	wire _06573_;
	wire _06574_;
	wire _06575_;
	wire _06576_;
	wire _06577_;
	wire _06578_;
	wire _06579_;
	wire _06580_;
	wire _06581_;
	wire _06582_;
	wire _06583_;
	wire _06584_;
	wire _06585_;
	wire _06586_;
	wire _06587_;
	wire _06588_;
	wire _06589_;
	wire _06590_;
	wire _06591_;
	wire _06592_;
	wire _06593_;
	wire _06594_;
	wire _06595_;
	wire _06596_;
	wire _06597_;
	wire _06598_;
	wire _06599_;
	wire _06600_;
	wire _06601_;
	wire _06602_;
	wire _06603_;
	wire _06604_;
	wire _06605_;
	wire _06606_;
	wire _06607_;
	wire _06608_;
	wire _06609_;
	wire _06610_;
	wire _06611_;
	wire _06612_;
	wire _06613_;
	wire _06614_;
	wire _06615_;
	wire _06616_;
	wire _06617_;
	wire _06618_;
	wire _06619_;
	wire _06620_;
	wire _06621_;
	wire _06622_;
	wire _06623_;
	wire _06624_;
	wire _06625_;
	wire _06626_;
	wire _06627_;
	wire _06628_;
	wire _06629_;
	wire _06630_;
	wire _06631_;
	wire _06632_;
	wire _06633_;
	wire _06634_;
	wire _06635_;
	wire _06636_;
	wire _06637_;
	wire _06638_;
	wire _06639_;
	wire _06640_;
	wire _06641_;
	wire _06642_;
	wire _06643_;
	wire _06644_;
	wire _06645_;
	wire _06646_;
	wire _06647_;
	wire _06648_;
	wire _06649_;
	wire _06650_;
	wire _06651_;
	wire _06652_;
	wire _06653_;
	wire _06654_;
	wire _06655_;
	wire _06656_;
	wire _06657_;
	wire _06658_;
	wire _06659_;
	wire _06660_;
	wire _06661_;
	wire _06662_;
	wire _06663_;
	wire _06664_;
	wire _06665_;
	wire _06666_;
	wire _06667_;
	wire _06668_;
	wire _06669_;
	wire _06670_;
	wire _06671_;
	wire _06672_;
	wire _06673_;
	wire _06674_;
	wire _06675_;
	wire _06676_;
	wire _06677_;
	wire _06678_;
	wire _06679_;
	wire _06680_;
	wire _06681_;
	wire _06682_;
	wire _06683_;
	wire _06684_;
	wire _06685_;
	wire _06686_;
	wire _06687_;
	wire _06688_;
	wire _06689_;
	wire _06690_;
	wire _06691_;
	wire _06692_;
	wire _06693_;
	wire _06694_;
	wire _06695_;
	wire _06696_;
	wire _06697_;
	wire _06698_;
	wire _06699_;
	wire _06700_;
	wire _06701_;
	wire _06702_;
	wire _06703_;
	wire _06704_;
	wire _06705_;
	wire _06706_;
	wire _06707_;
	wire _06708_;
	wire _06709_;
	wire _06710_;
	wire _06711_;
	wire _06712_;
	wire _06713_;
	wire _06714_;
	wire _06715_;
	wire _06716_;
	wire _06717_;
	wire _06718_;
	wire _06719_;
	wire _06720_;
	wire _06721_;
	wire _06722_;
	wire _06723_;
	wire _06724_;
	wire _06725_;
	wire _06726_;
	wire _06727_;
	wire _06728_;
	wire _06729_;
	wire _06730_;
	wire _06731_;
	wire _06732_;
	wire _06733_;
	wire _06734_;
	wire _06735_;
	wire _06736_;
	wire _06737_;
	wire _06738_;
	wire _06739_;
	wire _06740_;
	wire _06741_;
	wire _06742_;
	wire _06743_;
	wire _06744_;
	wire _06745_;
	wire _06746_;
	wire _06747_;
	wire _06748_;
	wire _06749_;
	wire _06750_;
	wire _06751_;
	wire _06752_;
	wire _06753_;
	wire _06754_;
	wire _06755_;
	wire _06756_;
	wire _06757_;
	wire _06758_;
	wire _06759_;
	wire _06760_;
	wire _06761_;
	wire _06762_;
	wire _06763_;
	wire _06764_;
	wire _06765_;
	wire _06766_;
	wire _06767_;
	wire _06768_;
	wire _06769_;
	wire _06770_;
	wire _06771_;
	wire _06772_;
	wire _06773_;
	wire _06774_;
	wire _06775_;
	wire _06776_;
	wire _06777_;
	wire _06778_;
	wire _06779_;
	wire _06780_;
	wire _06781_;
	wire _06782_;
	wire _06783_;
	wire _06784_;
	wire _06785_;
	wire _06786_;
	wire _06787_;
	wire _06788_;
	wire _06789_;
	wire _06790_;
	wire _06791_;
	wire _06792_;
	wire _06793_;
	wire _06794_;
	wire _06795_;
	wire _06796_;
	wire _06797_;
	wire _06798_;
	wire _06799_;
	wire _06800_;
	wire _06801_;
	wire _06802_;
	wire _06803_;
	wire _06804_;
	wire _06805_;
	wire _06806_;
	wire _06807_;
	wire _06808_;
	wire _06809_;
	wire _06810_;
	wire _06811_;
	wire _06812_;
	wire _06813_;
	wire _06814_;
	wire _06815_;
	wire _06816_;
	wire _06817_;
	wire _06818_;
	wire _06819_;
	wire _06820_;
	wire _06821_;
	wire _06822_;
	wire _06823_;
	wire _06824_;
	wire _06825_;
	wire _06826_;
	wire _06827_;
	wire _06828_;
	wire _06829_;
	wire _06830_;
	wire _06831_;
	wire _06832_;
	wire _06833_;
	wire _06834_;
	wire _06835_;
	wire _06836_;
	wire _06837_;
	wire _06838_;
	wire _06839_;
	wire _06840_;
	wire _06841_;
	wire _06842_;
	wire _06843_;
	wire _06844_;
	wire _06845_;
	wire _06846_;
	wire _06847_;
	wire _06848_;
	wire _06849_;
	wire _06850_;
	wire _06851_;
	wire _06852_;
	wire _06853_;
	wire _06854_;
	wire _06855_;
	wire _06856_;
	wire _06857_;
	wire _06858_;
	wire _06859_;
	wire _06860_;
	wire _06861_;
	wire _06862_;
	wire _06863_;
	wire _06864_;
	wire _06865_;
	wire _06866_;
	wire _06867_;
	wire _06868_;
	wire _06869_;
	wire _06870_;
	wire _06871_;
	wire _06872_;
	wire _06873_;
	wire _06874_;
	wire _06875_;
	wire _06876_;
	wire _06877_;
	wire _06878_;
	wire _06879_;
	wire _06880_;
	wire _06881_;
	wire _06882_;
	wire _06883_;
	wire _06884_;
	wire _06885_;
	wire _06886_;
	wire _06887_;
	wire _06888_;
	wire _06889_;
	wire _06890_;
	wire _06891_;
	wire _06892_;
	wire _06893_;
	wire _06894_;
	wire _06895_;
	wire _06896_;
	wire _06897_;
	wire _06898_;
	wire _06899_;
	wire _06900_;
	wire _06901_;
	wire _06902_;
	wire _06903_;
	wire _06904_;
	wire _06905_;
	wire _06906_;
	wire _06907_;
	wire _06908_;
	wire _06909_;
	wire _06910_;
	wire _06911_;
	wire _06912_;
	wire _06913_;
	wire _06914_;
	wire _06915_;
	wire _06916_;
	wire _06917_;
	wire _06918_;
	wire _06919_;
	wire _06920_;
	wire _06921_;
	wire _06922_;
	wire _06923_;
	wire _06924_;
	wire _06925_;
	wire _06926_;
	wire _06927_;
	wire _06928_;
	wire _06929_;
	wire _06930_;
	wire _06931_;
	wire _06932_;
	wire _06933_;
	wire _06934_;
	wire _06935_;
	wire _06936_;
	wire _06937_;
	wire _06938_;
	wire _06939_;
	wire _06940_;
	wire _06941_;
	wire _06942_;
	wire _06943_;
	wire _06944_;
	wire _06945_;
	wire _06946_;
	wire _06947_;
	wire _06948_;
	wire _06949_;
	wire _06950_;
	wire _06951_;
	wire _06952_;
	wire _06953_;
	wire _06954_;
	wire _06955_;
	wire _06956_;
	wire _06957_;
	wire _06958_;
	wire _06959_;
	wire _06960_;
	wire _06961_;
	wire _06962_;
	wire _06963_;
	wire _06964_;
	wire _06965_;
	wire _06966_;
	wire _06967_;
	wire _06968_;
	wire _06969_;
	wire _06970_;
	wire _06971_;
	wire _06972_;
	wire _06973_;
	wire _06974_;
	wire _06975_;
	wire _06976_;
	wire _06977_;
	wire _06978_;
	wire _06979_;
	wire _06980_;
	wire _06981_;
	wire _06982_;
	wire _06983_;
	wire _06984_;
	wire _06985_;
	wire _06986_;
	wire _06987_;
	wire _06988_;
	wire _06989_;
	wire _06990_;
	wire _06991_;
	wire _06992_;
	wire _06993_;
	wire _06994_;
	wire _06995_;
	wire _06996_;
	wire _06997_;
	wire _06998_;
	wire _06999_;
	wire _07000_;
	wire _07001_;
	wire _07002_;
	wire _07003_;
	wire _07004_;
	wire _07005_;
	wire _07006_;
	wire _07007_;
	wire _07008_;
	wire _07009_;
	wire _07010_;
	wire _07011_;
	wire _07012_;
	wire _07013_;
	wire _07014_;
	wire _07015_;
	wire _07016_;
	wire _07017_;
	wire _07018_;
	wire _07019_;
	wire _07020_;
	wire _07021_;
	wire _07022_;
	wire _07023_;
	wire _07024_;
	wire _07025_;
	wire _07026_;
	wire _07027_;
	wire _07028_;
	wire _07029_;
	wire _07030_;
	wire _07031_;
	wire _07032_;
	wire _07033_;
	wire _07034_;
	wire _07035_;
	wire _07036_;
	wire _07037_;
	wire _07038_;
	wire _07039_;
	wire _07040_;
	wire _07041_;
	wire _07042_;
	wire _07043_;
	wire _07044_;
	wire _07045_;
	wire _07046_;
	wire _07047_;
	wire _07048_;
	wire _07049_;
	wire _07050_;
	wire _07051_;
	wire _07052_;
	wire _07053_;
	wire _07054_;
	wire _07055_;
	wire _07056_;
	wire _07057_;
	wire _07058_;
	wire _07059_;
	wire _07060_;
	wire _07061_;
	wire _07062_;
	wire _07063_;
	wire _07064_;
	wire _07065_;
	wire _07066_;
	wire _07067_;
	wire _07068_;
	wire _07069_;
	wire _07070_;
	wire _07071_;
	wire _07072_;
	wire _07073_;
	wire _07074_;
	wire _07075_;
	wire _07076_;
	wire _07077_;
	wire _07078_;
	wire _07079_;
	wire _07080_;
	wire _07081_;
	wire _07082_;
	wire _07083_;
	wire _07084_;
	wire _07085_;
	wire _07086_;
	wire _07087_;
	wire _07088_;
	wire _07089_;
	wire _07090_;
	wire _07091_;
	wire _07092_;
	wire _07093_;
	wire _07094_;
	wire _07095_;
	wire _07096_;
	wire _07097_;
	wire _07098_;
	wire _07099_;
	wire _07100_;
	wire _07101_;
	wire _07102_;
	wire _07103_;
	wire _07104_;
	wire _07105_;
	wire _07106_;
	wire _07107_;
	wire _07108_;
	wire _07109_;
	wire _07110_;
	wire _07111_;
	wire _07112_;
	wire _07113_;
	wire _07114_;
	wire _07115_;
	wire _07116_;
	wire _07117_;
	wire _07118_;
	wire _07119_;
	wire _07120_;
	wire _07121_;
	wire _07122_;
	wire _07123_;
	wire _07124_;
	wire _07125_;
	wire _07126_;
	wire _07127_;
	wire _07128_;
	wire _07129_;
	wire _07130_;
	wire _07131_;
	wire _07132_;
	wire _07133_;
	wire _07134_;
	wire _07135_;
	wire _07136_;
	wire _07137_;
	wire _07138_;
	wire _07139_;
	wire _07140_;
	wire _07141_;
	wire _07142_;
	wire _07143_;
	wire _07144_;
	wire _07145_;
	wire _07146_;
	wire _07147_;
	wire _07148_;
	wire _07149_;
	wire _07150_;
	wire _07151_;
	wire _07152_;
	wire _07153_;
	wire _07154_;
	wire _07155_;
	wire _07156_;
	wire _07157_;
	wire _07158_;
	wire _07159_;
	wire _07160_;
	wire _07161_;
	wire _07162_;
	wire _07163_;
	wire _07164_;
	wire _07165_;
	wire _07166_;
	wire _07167_;
	wire _07168_;
	wire _07169_;
	wire _07170_;
	wire _07171_;
	wire _07172_;
	wire _07173_;
	wire _07174_;
	wire _07175_;
	wire _07176_;
	wire _07177_;
	wire _07178_;
	wire _07179_;
	wire _07180_;
	wire _07181_;
	wire _07182_;
	wire _07183_;
	wire _07184_;
	wire _07185_;
	wire _07186_;
	wire _07187_;
	wire _07188_;
	wire _07189_;
	wire _07190_;
	wire _07191_;
	wire _07192_;
	wire _07193_;
	wire _07194_;
	wire _07195_;
	wire _07196_;
	wire _07197_;
	wire _07198_;
	wire _07199_;
	wire _07200_;
	wire _07201_;
	wire _07202_;
	wire _07203_;
	wire _07204_;
	wire _07205_;
	wire _07206_;
	wire _07207_;
	wire _07208_;
	wire _07209_;
	wire _07210_;
	wire _07211_;
	wire _07212_;
	wire _07213_;
	wire _07214_;
	wire _07215_;
	wire _07216_;
	wire _07217_;
	wire _07218_;
	wire _07219_;
	wire _07220_;
	wire _07221_;
	wire _07222_;
	wire _07223_;
	wire _07224_;
	wire _07225_;
	wire _07226_;
	wire _07227_;
	wire _07228_;
	wire _07229_;
	wire _07230_;
	wire _07231_;
	wire _07232_;
	wire _07233_;
	wire _07234_;
	wire _07235_;
	wire _07236_;
	wire _07237_;
	wire _07238_;
	wire _07239_;
	wire _07240_;
	wire _07241_;
	wire _07242_;
	wire _07243_;
	wire _07244_;
	wire _07245_;
	wire _07246_;
	wire _07247_;
	wire _07248_;
	wire _07249_;
	wire _07250_;
	wire _07251_;
	wire _07252_;
	wire _07253_;
	wire _07254_;
	wire _07255_;
	wire _07256_;
	wire _07257_;
	wire _07258_;
	wire _07259_;
	wire _07260_;
	wire _07261_;
	wire _07262_;
	wire _07263_;
	wire _07264_;
	wire _07265_;
	wire _07266_;
	wire _07267_;
	wire _07268_;
	wire _07269_;
	wire _07270_;
	wire _07271_;
	wire _07272_;
	wire _07273_;
	wire _07274_;
	wire _07275_;
	wire _07276_;
	wire _07277_;
	wire _07278_;
	wire _07279_;
	wire _07280_;
	wire _07281_;
	wire _07282_;
	wire _07283_;
	wire _07284_;
	wire _07285_;
	wire _07286_;
	wire _07287_;
	wire _07288_;
	wire _07289_;
	wire _07290_;
	wire _07291_;
	wire _07292_;
	wire _07293_;
	wire _07294_;
	wire _07295_;
	wire _07296_;
	wire _07297_;
	wire _07298_;
	wire _07299_;
	wire _07300_;
	wire _07301_;
	wire _07302_;
	wire _07303_;
	wire _07304_;
	wire _07305_;
	wire _07306_;
	wire _07307_;
	wire _07308_;
	wire _07309_;
	wire _07310_;
	wire _07311_;
	wire _07312_;
	wire _07313_;
	wire _07314_;
	wire _07315_;
	wire _07316_;
	wire _07317_;
	wire _07318_;
	wire _07319_;
	wire _07320_;
	wire _07321_;
	wire _07322_;
	wire _07323_;
	wire _07324_;
	wire _07325_;
	wire _07326_;
	wire _07327_;
	wire _07328_;
	wire _07329_;
	wire _07330_;
	wire _07331_;
	wire _07332_;
	wire _07333_;
	wire _07334_;
	wire _07335_;
	wire _07336_;
	wire _07337_;
	wire _07338_;
	wire _07339_;
	wire _07340_;
	wire _07341_;
	wire _07342_;
	wire _07343_;
	wire _07344_;
	wire _07345_;
	wire _07346_;
	wire _07347_;
	wire _07348_;
	wire _07349_;
	wire _07350_;
	wire _07351_;
	wire _07352_;
	wire _07353_;
	wire _07354_;
	wire _07355_;
	wire _07356_;
	wire _07357_;
	wire _07358_;
	wire _07359_;
	wire _07360_;
	wire _07361_;
	wire _07362_;
	wire _07363_;
	wire _07364_;
	wire _07365_;
	wire _07366_;
	wire _07367_;
	wire _07368_;
	wire _07369_;
	wire _07370_;
	wire _07371_;
	wire _07372_;
	wire _07373_;
	wire _07374_;
	wire _07375_;
	wire _07376_;
	wire _07377_;
	wire _07378_;
	wire _07379_;
	wire _07380_;
	wire _07381_;
	wire _07382_;
	wire _07383_;
	wire _07384_;
	wire _07385_;
	wire _07386_;
	wire _07387_;
	wire _07388_;
	wire _07389_;
	wire _07390_;
	wire _07391_;
	wire _07392_;
	wire _07393_;
	wire _07394_;
	wire _07395_;
	wire _07396_;
	wire _07397_;
	wire _07398_;
	wire _07399_;
	wire _07400_;
	wire _07401_;
	wire _07402_;
	wire _07403_;
	wire _07404_;
	wire _07405_;
	wire _07406_;
	wire _07407_;
	wire _07408_;
	wire _07409_;
	wire _07410_;
	wire _07411_;
	wire _07412_;
	wire _07413_;
	wire _07414_;
	wire _07415_;
	wire _07416_;
	wire _07417_;
	wire _07418_;
	wire _07419_;
	wire _07420_;
	wire _07421_;
	wire _07422_;
	wire _07423_;
	wire _07424_;
	wire _07425_;
	wire _07426_;
	wire _07427_;
	wire _07428_;
	wire _07429_;
	wire _07430_;
	wire _07431_;
	wire _07432_;
	wire _07433_;
	wire _07434_;
	wire _07435_;
	wire _07436_;
	wire _07437_;
	wire _07438_;
	wire _07439_;
	wire _07440_;
	wire _07441_;
	wire _07442_;
	wire _07443_;
	wire _07444_;
	wire _07445_;
	wire _07446_;
	wire _07447_;
	wire _07448_;
	wire _07449_;
	wire _07450_;
	wire _07451_;
	wire _07452_;
	wire _07453_;
	wire _07454_;
	wire _07455_;
	wire _07456_;
	wire _07457_;
	wire _07458_;
	wire _07459_;
	wire _07460_;
	wire _07461_;
	wire _07462_;
	wire _07463_;
	wire _07464_;
	wire _07465_;
	wire _07466_;
	wire _07467_;
	wire _07468_;
	wire _07469_;
	wire _07470_;
	wire _07471_;
	wire _07472_;
	wire _07473_;
	wire _07474_;
	wire _07475_;
	wire _07476_;
	wire _07477_;
	wire _07478_;
	wire _07479_;
	wire _07480_;
	wire _07481_;
	wire _07482_;
	wire _07483_;
	wire _07484_;
	wire _07485_;
	wire _07486_;
	wire _07487_;
	wire _07488_;
	wire _07489_;
	wire _07490_;
	wire _07491_;
	wire _07492_;
	wire _07493_;
	wire _07494_;
	wire _07495_;
	wire _07496_;
	wire _07497_;
	wire _07498_;
	wire _07499_;
	wire _07500_;
	wire _07501_;
	wire _07502_;
	wire _07503_;
	wire _07504_;
	wire _07505_;
	wire _07506_;
	wire _07507_;
	wire _07508_;
	wire _07509_;
	wire _07510_;
	input wire [13:0] io_in;
	output wire [13:0] io_out;
	wire \mchip.clock ;
	wire [11:0] \mchip.io_in ;
	wire [11:0] \mchip.io_out ;
	wire \mchip.reset ;
	wire [7:0] \mchip.val ;
	assign _01208_ = ~io_in[8];
	assign _01319_ = ~io_in[3];
	assign _01430_ = ~(io_in[1] & io_in[2]);
	assign _01541_ = _01430_ | _01319_;
	assign _01652_ = _01541_ | io_in[6];
	assign _01763_ = _01652_ | io_in[7];
	assign _01874_ = _01208_ & ~_01763_;
	assign _01985_ = ~io_in[11];
	assign _02096_ = ~io_in[9];
	assign _02207_ = ~io_in[7];
	assign _02317_ = ~(io_in[1] & io_in[0]);
	assign _02428_ = _02317_ | io_in[2];
	assign _02539_ = _02428_ | io_in[4];
	assign _02650_ = _02539_ | _02207_;
	assign _02761_ = _02650_ | _01208_;
	assign _02872_ = _02761_ | _02096_;
	assign _02983_ = _01985_ & ~_02872_;
	assign _03094_ = ~io_in[5];
	assign _03205_ = io_in[3] | ~io_in[2];
	assign _03316_ = _03205_ | _03094_;
	assign _03427_ = _03316_ | io_in[8];
	assign _03537_ = _03427_ | io_in[9];
	assign _03648_ = io_in[10] & ~_03537_;
	assign _03759_ = ~io_in[6];
	assign _03870_ = io_in[1] | io_in[2];
	assign _03981_ = _03870_ | io_in[3];
	assign _04092_ = _03981_ | io_in[5];
	assign _04203_ = _04092_ | _03759_;
	assign _04314_ = _04203_ | io_in[9];
	assign _04425_ = _04314_ | io_in[10];
	assign _04536_ = io_in[11] & ~_04425_;
	assign _04647_ = io_in[1] | ~io_in[2];
	assign _04758_ = _04647_ | io_in[4];
	assign _04868_ = _04758_ | _03094_;
	assign _04979_ = _04868_ | io_in[7];
	assign _05090_ = io_in[11] & ~_04979_;
	assign _05201_ = _03870_ | io_in[5];
	assign _05312_ = _05201_ | io_in[6];
	assign _05423_ = _05312_ | io_in[8];
	assign _05534_ = _05423_ | _02096_;
	assign _05645_ = _05534_ | io_in[10];
	assign _05756_ = io_in[11] & ~_05645_;
	assign _05867_ = _04647_ | io_in[6];
	assign _05978_ = _05867_ | io_in[7];
	assign _06088_ = _05978_ | _02096_;
	assign _06199_ = _01985_ & ~_06088_;
	assign _06310_ = ~io_in[10];
	assign _06421_ = ~io_in[2];
	assign _06532_ = io_in[0] | ~io_in[1];
	assign _06643_ = _06532_ | _06421_;
	assign _06754_ = _06643_ | _01319_;
	assign _06865_ = _06754_ | io_in[4];
	assign _06976_ = _06865_ | _03759_;
	assign _07087_ = _06310_ & ~_06976_;
	assign _07198_ = io_in[1] | io_in[0];
	assign _07246_ = _07198_ | io_in[2];
	assign _07257_ = _07246_ | _01319_;
	assign _07268_ = _07257_ | io_in[8];
	assign _07279_ = _07268_ | io_in[9];
	assign _07290_ = _06310_ & ~_07279_;
	assign _07301_ = _04647_ | io_in[3];
	assign _07312_ = _07301_ | io_in[6];
	assign _07323_ = _07312_ | _02096_;
	assign _07334_ = _07323_ | io_in[10];
	assign _07345_ = _01985_ & ~_07334_;
	assign _07356_ = io_in[2] | ~io_in[0];
	assign _07367_ = _07356_ | _01319_;
	assign _07378_ = _07367_ | io_in[4];
	assign _07389_ = _07378_ | io_in[6];
	assign _07400_ = _07389_ | io_in[7];
	assign _07411_ = io_in[10] & ~_07400_;
	assign _07422_ = ~io_in[4];
	assign _07433_ = io_in[2] | ~io_in[1];
	assign _07444_ = _07433_ | _01319_;
	assign _07455_ = _07444_ | _07422_;
	assign _07466_ = _07455_ | _02207_;
	assign _07477_ = _07466_ | io_in[8];
	assign _07488_ = _06310_ & ~_07477_;
	assign _07499_ = _07198_ | _06421_;
	assign _07510_ = _07499_ | io_in[3];
	assign _00010_ = _07510_ | io_in[4];
	assign _00021_ = _00010_ | io_in[10];
	assign _00032_ = io_in[11] & ~_00021_;
	assign _00043_ = io_in[2] | io_in[0];
	assign _00054_ = _00043_ | io_in[4];
	assign _00065_ = _00054_ | io_in[5];
	assign _00076_ = _00065_ | _02207_;
	assign _00087_ = _00076_ | _01208_;
	assign _00098_ = _00087_ | _02096_;
	assign _00109_ = io_in[10] & ~_00098_;
	assign _00120_ = _07198_ | io_in[3];
	assign _00131_ = _00120_ | io_in[4];
	assign _00142_ = _00131_ | io_in[7];
	assign _00153_ = _00142_ | _06310_;
	assign _00163_ = _01985_ & ~_00153_;
	assign _00174_ = _01541_ | io_in[4];
	assign _00185_ = _00174_ | _02207_;
	assign _00196_ = _00185_ | _02096_;
	assign _00207_ = _06310_ & ~_00196_;
	assign _00218_ = _07246_ | io_in[5];
	assign _00229_ = _00218_ | io_in[7];
	assign _00240_ = _00229_ | _01208_;
	assign _00251_ = _00240_ | io_in[10];
	assign _00262_ = _01985_ & ~_00251_;
	assign _00273_ = _03981_ | _03094_;
	assign _00284_ = _00273_ | _03759_;
	assign _00295_ = _00284_ | io_in[7];
	assign _00306_ = io_in[9] & ~_00295_;
	assign _00317_ = ~(io_in[1] & io_in[3]);
	assign _00328_ = _00317_ | io_in[4];
	assign _00339_ = _00328_ | io_in[7];
	assign _00350_ = _00339_ | io_in[9];
	assign _00361_ = _00350_ | io_in[10];
	assign _00372_ = _01985_ & ~_00361_;
	assign _00383_ = _07356_ | io_in[3];
	assign _00394_ = _00383_ | _03759_;
	assign _00405_ = _00394_ | io_in[7];
	assign _00416_ = _00405_ | io_in[8];
	assign _00427_ = io_in[9] & ~_00416_;
	assign _00438_ = ~(io_in[3] & io_in[0]);
	assign _00449_ = _00438_ | _03094_;
	assign _00460_ = _00449_ | _02096_;
	assign _00471_ = _01985_ & ~_00460_;
	assign _00482_ = io_in[1] | ~io_in[0];
	assign _00493_ = _00482_ | _06421_;
	assign _00504_ = _00493_ | io_in[4];
	assign _00515_ = _00504_ | _02207_;
	assign _00526_ = _00515_ | _06310_;
	assign _00537_ = _01985_ & ~_00526_;
	assign _00548_ = ~(io_in[2] & io_in[0]);
	assign _00559_ = _00548_ | io_in[4];
	assign _00570_ = _00559_ | io_in[5];
	assign _00581_ = _00570_ | _02207_;
	assign _00592_ = _00581_ | _01208_;
	assign _00603_ = _02096_ & ~_00592_;
	assign _00614_ = _00559_ | io_in[6];
	assign _00625_ = _00614_ | _02207_;
	assign _00636_ = _00625_ | _02096_;
	assign _00647_ = io_in[11] & ~_00636_;
	assign _00658_ = io_in[3] | io_in[2];
	assign _00669_ = _00658_ | io_in[5];
	assign _00680_ = _00669_ | _02207_;
	assign _00691_ = _00680_ | _01208_;
	assign _00702_ = _00691_ | _02096_;
	assign _00713_ = _01985_ & ~_00702_;
	assign _00724_ = _07198_ | _03094_;
	assign _00735_ = _00724_ | io_in[8];
	assign _00746_ = io_in[9] & ~_00735_;
	assign _00757_ = _06532_ | io_in[3];
	assign _00768_ = _00757_ | _07422_;
	assign _00779_ = _00768_ | io_in[8];
	assign _00790_ = _00779_ | io_in[9];
	assign _00801_ = _01985_ & ~_00790_;
	assign _00812_ = _06532_ | _01319_;
	assign _00823_ = _00812_ | io_in[4];
	assign _00834_ = _00823_ | _02207_;
	assign _00845_ = _00834_ | _01208_;
	assign _00856_ = _00845_ | _02096_;
	assign _00867_ = _01985_ & ~_00856_;
	assign _00878_ = _07433_ | io_in[3];
	assign _00889_ = _00878_ | _07422_;
	assign _00900_ = _00889_ | io_in[6];
	assign _00911_ = _00900_ | io_in[9];
	assign _00922_ = _06310_ & ~_00911_;
	assign _00933_ = _02317_ | io_in[4];
	assign _00944_ = _00933_ | io_in[7];
	assign _00955_ = _00944_ | io_in[8];
	assign _00966_ = _00955_ | io_in[9];
	assign _00976_ = _06310_ & ~_00966_;
	assign _00987_ = _00493_ | _07422_;
	assign _00998_ = _00987_ | _03759_;
	assign _01009_ = _00998_ | io_in[9];
	assign _01020_ = _01985_ & ~_01009_;
	assign _01031_ = _00482_ | io_in[2];
	assign _01042_ = _01031_ | io_in[3];
	assign _01053_ = _01042_ | _03759_;
	assign _01064_ = _01053_ | _02207_;
	assign _01075_ = _01208_ & ~_01064_;
	assign _01086_ = io_in[0] | ~io_in[3];
	assign _01097_ = _01086_ | _07422_;
	assign _01108_ = _01097_ | _03759_;
	assign _01119_ = _01108_ | _02207_;
	assign _01130_ = _01119_ | io_in[9];
	assign _01141_ = _06310_ & ~_01130_;
	assign _01152_ = _00658_ | io_in[4];
	assign _01163_ = _01152_ | _03759_;
	assign _01174_ = _01163_ | io_in[7];
	assign _01185_ = _01174_ | _02096_;
	assign _01196_ = _01185_ | _06310_;
	assign _01207_ = _01985_ & ~_01196_;
	assign _01219_ = io_in[3] | ~io_in[1];
	assign _01230_ = _01219_ | io_in[5];
	assign _01241_ = _01230_ | io_in[6];
	assign _01252_ = _01241_ | _01208_;
	assign _01263_ = _01252_ | _02096_;
	assign _01274_ = _01263_ | _06310_;
	assign _01285_ = _01985_ & ~_01274_;
	assign _01296_ = _07198_ | _01319_;
	assign _01307_ = _01296_ | _07422_;
	assign _01318_ = _01307_ | _03759_;
	assign _01330_ = _01318_ | _06310_;
	assign _01341_ = _01985_ & ~_01330_;
	assign _01352_ = io_in[3] | io_in[0];
	assign _01363_ = _01352_ | io_in[4];
	assign _01374_ = _01363_ | io_in[6];
	assign _01385_ = _01374_ | _02207_;
	assign _01396_ = _01385_ | io_in[8];
	assign _01407_ = _01396_ | _02096_;
	assign _01418_ = _01985_ & ~_01407_;
	assign _01429_ = _01219_ | _07422_;
	assign _01441_ = _01429_ | _02207_;
	assign _01452_ = _01441_ | _01208_;
	assign _01463_ = _01452_ | _02096_;
	assign _01474_ = _01985_ & ~_01463_;
	assign _01485_ = _07301_ | io_in[4];
	assign _01496_ = _01485_ | io_in[5];
	assign _01507_ = _01496_ | _03759_;
	assign _01518_ = _01507_ | io_in[8];
	assign _01529_ = io_in[9] & ~_01518_;
	assign _01540_ = _07356_ | _03759_;
	assign _01552_ = _01540_ | _02207_;
	assign _01563_ = _01552_ | io_in[8];
	assign _01574_ = _01563_ | io_in[9];
	assign _01585_ = io_in[10] & ~_01574_;
	assign _01596_ = _00043_ | _01319_;
	assign _01607_ = _01596_ | io_in[4];
	assign _01618_ = _01607_ | _02207_;
	assign _01629_ = _01618_ | _01208_;
	assign _01640_ = io_in[9] & ~_01629_;
	assign _01651_ = _00724_ | io_in[6];
	assign _01663_ = _01651_ | io_in[8];
	assign _01674_ = io_in[10] & ~_01663_;
	assign _01685_ = _01352_ | _03094_;
	assign _01696_ = _01685_ | _03759_;
	assign _01707_ = _01696_ | _01208_;
	assign _01718_ = _01985_ & ~_01707_;
	assign _01729_ = _00493_ | _02207_;
	assign _01740_ = _01729_ | io_in[8];
	assign _01751_ = io_in[10] & ~_01740_;
	assign _01762_ = _00054_ | _02207_;
	assign _01774_ = _01762_ | _01208_;
	assign _01785_ = _01774_ | _06310_;
	assign _01796_ = _01985_ & ~_01785_;
	assign _01807_ = io_in[2] | ~io_in[3];
	assign _01818_ = _01807_ | _07422_;
	assign _01829_ = _01818_ | _03759_;
	assign _01840_ = _01829_ | _01208_;
	assign _01851_ = _01840_ | _02096_;
	assign _01862_ = _01985_ & ~_01851_;
	assign _01873_ = _04647_ | _02207_;
	assign _01885_ = _01873_ | io_in[9];
	assign _01896_ = io_in[10] & ~_01885_;
	assign _01907_ = io_in[2] | ~io_in[4];
	assign _01918_ = _01907_ | _03759_;
	assign _01929_ = _01918_ | _02207_;
	assign _01940_ = _01929_ | io_in[9];
	assign _01951_ = io_in[11] & ~_01940_;
	assign _01962_ = io_in[0] | ~io_in[2];
	assign _01973_ = _01962_ | _03759_;
	assign _01984_ = _01973_ | io_in[7];
	assign _01996_ = _01984_ | io_in[8];
	assign _02007_ = io_in[9] & ~_01996_;
	assign _02018_ = _00043_ | io_in[3];
	assign _02029_ = _02018_ | _07422_;
	assign _02040_ = _02029_ | io_in[6];
	assign _02051_ = _02040_ | io_in[9];
	assign _02062_ = _01985_ & ~_02051_;
	assign _02073_ = _00724_ | _03759_;
	assign _02084_ = _02073_ | io_in[7];
	assign _02095_ = io_in[9] & ~_02084_;
	assign _02107_ = _01086_ | io_in[5];
	assign _02118_ = _02107_ | io_in[6];
	assign _02129_ = _02118_ | io_in[8];
	assign _02140_ = _02129_ | _02096_;
	assign _02151_ = io_in[10] & ~_02140_;
	assign _02162_ = _07246_ | io_in[7];
	assign _02173_ = _02162_ | io_in[8];
	assign _02184_ = _02173_ | _06310_;
	assign _02195_ = _01985_ & ~_02184_;
	assign _02206_ = io_in[1] | io_in[3];
	assign _02218_ = _02206_ | io_in[4];
	assign _02229_ = _02218_ | _03094_;
	assign _02240_ = _02229_ | io_in[6];
	assign _02251_ = _02240_ | _02207_;
	assign _02262_ = io_in[10] & ~_02251_;
	assign _02272_ = _01042_ | _07422_;
	assign _02283_ = _02272_ | _02207_;
	assign _02294_ = _01208_ & ~_02283_;
	assign _02305_ = _04758_ | io_in[5];
	assign _02316_ = _02305_ | io_in[6];
	assign _02328_ = _02316_ | _02207_;
	assign _02339_ = _02096_ & ~_02328_;
	assign _02350_ = _02428_ | _03094_;
	assign _02361_ = _02350_ | _03759_;
	assign _02372_ = io_in[10] & ~_02361_;
	assign _02383_ = io_in[1] | ~io_in[5];
	assign _02394_ = _02383_ | io_in[7];
	assign _02405_ = _02394_ | io_in[9];
	assign _02416_ = io_in[11] & ~_02405_;
	assign _02427_ = _01097_ | io_in[6];
	assign _02439_ = _02427_ | _02207_;
	assign _02450_ = _02439_ | _01208_;
	assign _02461_ = io_in[11] & ~_02450_;
	assign _02472_ = _01541_ | _02207_;
	assign _02483_ = _02472_ | io_in[9];
	assign _02494_ = io_in[11] & ~_02483_;
	assign _02505_ = _01962_ | io_in[3];
	assign _02516_ = _02505_ | io_in[6];
	assign _02527_ = _02516_ | io_in[8];
	assign _02538_ = _02527_ | io_in[9];
	assign _02550_ = io_in[11] & ~_02538_;
	assign _02561_ = io_in[1] | io_in[4];
	assign _02572_ = _02561_ | io_in[5];
	assign _02583_ = _02572_ | io_in[6];
	assign _02594_ = _02583_ | _01208_;
	assign _02605_ = _02594_ | _02096_;
	assign _02616_ = _02605_ | _06310_;
	assign _02627_ = io_in[11] & ~_02616_;
	assign _02638_ = _01973_ | io_in[8];
	assign _02649_ = _02638_ | _02096_;
	assign _02661_ = io_in[11] & ~_02649_;
	assign _02672_ = _06532_ | io_in[2];
	assign _02683_ = _02672_ | io_in[5];
	assign _02694_ = _02683_ | io_in[6];
	assign _02705_ = _02694_ | _02207_;
	assign _02716_ = io_in[9] & ~_02705_;
	assign _02727_ = _01962_ | io_in[4];
	assign _02738_ = _02727_ | io_in[6];
	assign _02749_ = _02738_ | io_in[9];
	assign _02760_ = io_in[10] & ~_02749_;
	assign _02772_ = _02317_ | _03094_;
	assign _02783_ = _02772_ | _03759_;
	assign _02794_ = _02783_ | _01208_;
	assign _02805_ = io_in[11] & ~_02794_;
	assign _02816_ = _02505_ | io_in[5];
	assign _02827_ = _02816_ | io_in[7];
	assign _02838_ = _02827_ | io_in[10];
	assign _02849_ = io_in[11] & ~_02838_;
	assign _02860_ = _07444_ | io_in[4];
	assign _02871_ = _02860_ | io_in[6];
	assign _02883_ = _02871_ | _02207_;
	assign _02894_ = _02883_ | io_in[8];
	assign _02905_ = _02096_ & ~_02894_;
	assign _02916_ = _00438_ | _07422_;
	assign _02927_ = _02916_ | _02207_;
	assign _02938_ = _02927_ | _02096_;
	assign _02949_ = _02938_ | _06310_;
	assign _02960_ = _01985_ & ~_02949_;
	assign _02971_ = _02317_ | io_in[3];
	assign _02982_ = _02971_ | _07422_;
	assign _02994_ = _02982_ | io_in[5];
	assign _03005_ = _02994_ | io_in[6];
	assign _03016_ = _02207_ & ~_03005_;
	assign _03027_ = _07510_ | _03759_;
	assign _03038_ = _03027_ | io_in[8];
	assign _03049_ = io_in[9] & ~_03038_;
	assign _03060_ = _00482_ | io_in[5];
	assign _03071_ = _03060_ | _02207_;
	assign _03082_ = _03071_ | io_in[8];
	assign _03093_ = _03082_ | io_in[9];
	assign _03105_ = io_in[10] & ~_03093_;
	assign _03116_ = _07257_ | io_in[5];
	assign _03127_ = _03116_ | _03759_;
	assign _03138_ = _02096_ & ~_03127_;
	assign _03149_ = _00482_ | io_in[3];
	assign _03160_ = _03149_ | io_in[5];
	assign _03171_ = _03160_ | io_in[6];
	assign _03182_ = _03171_ | _02207_;
	assign _03193_ = io_in[11] & ~_03182_;
	assign _03204_ = _02672_ | io_in[4];
	assign _03216_ = _03204_ | _03759_;
	assign _03227_ = _03216_ | _02207_;
	assign _03238_ = io_in[8] & ~_03227_;
	assign _03249_ = _04647_ | _01319_;
	assign _03260_ = _03249_ | io_in[4];
	assign _03271_ = _03260_ | io_in[7];
	assign _03282_ = _03271_ | _02096_;
	assign _03293_ = _01985_ & ~_03282_;
	assign _03304_ = _00548_ | _01319_;
	assign _03315_ = _03304_ | _07422_;
	assign _03327_ = _03315_ | _02207_;
	assign _03338_ = _03327_ | _02096_;
	assign _03349_ = _01985_ & ~_03338_;
	assign _03360_ = _07499_ | _03759_;
	assign _03371_ = _03360_ | _02207_;
	assign _03382_ = _03371_ | _06310_;
	assign _03393_ = _01985_ & ~_03382_;
	assign _03404_ = _00482_ | io_in[4];
	assign _03415_ = _03404_ | io_in[5];
	assign _03426_ = _03415_ | _03759_;
	assign _03438_ = _03426_ | io_in[8];
	assign _03449_ = io_in[10] & ~_03438_;
	assign _03460_ = _01540_ | io_in[8];
	assign _03471_ = _03460_ | _02096_;
	assign _03482_ = io_in[11] & ~_03471_;
	assign _03493_ = _01152_ | io_in[5];
	assign _03504_ = _03493_ | _06310_;
	assign _03515_ = _01985_ & ~_03504_;
	assign _03526_ = io_in[3] | ~io_in[0];
	assign _03536_ = _03526_ | io_in[5];
	assign _03548_ = _03536_ | io_in[7];
	assign _03559_ = _03548_ | _01208_;
	assign _03570_ = _03559_ | io_in[10];
	assign _03581_ = io_in[11] & ~_03570_;
	assign _03592_ = _03526_ | io_in[4];
	assign _03603_ = _03592_ | io_in[5];
	assign _03614_ = _03603_ | io_in[6];
	assign _03625_ = _03614_ | _02207_;
	assign _03636_ = io_in[10] & ~_03625_;
	assign _03647_ = _02916_ | _03759_;
	assign _03659_ = _03647_ | _02096_;
	assign _03670_ = _06310_ & ~_03659_;
	assign _03681_ = _01296_ | io_in[5];
	assign _03692_ = _03681_ | _01208_;
	assign _03703_ = _03692_ | io_in[9];
	assign _03714_ = io_in[10] & ~_03703_;
	assign _03725_ = _01962_ | _01319_;
	assign _03736_ = _03725_ | _07422_;
	assign _03747_ = _03736_ | io_in[6];
	assign _03758_ = _03747_ | _01208_;
	assign _03770_ = _01985_ & ~_03758_;
	assign _03781_ = _07356_ | _07422_;
	assign _03792_ = _03781_ | io_in[8];
	assign _03803_ = _03792_ | _02096_;
	assign _03814_ = io_in[11] & ~_03803_;
	assign _03825_ = _07433_ | _03759_;
	assign _03836_ = _03825_ | _02207_;
	assign _03847_ = _03836_ | _02096_;
	assign _03858_ = _03847_ | io_in[10];
	assign _03869_ = _01985_ & ~_03858_;
	assign _03881_ = _07433_ | io_in[4];
	assign _03892_ = _03881_ | io_in[5];
	assign _03903_ = _03892_ | io_in[8];
	assign _03914_ = _03903_ | _02096_;
	assign _03925_ = io_in[10] & ~_03914_;
	assign _03936_ = _02505_ | _03094_;
	assign _03947_ = _03936_ | io_in[7];
	assign _03958_ = _03947_ | _02096_;
	assign _03969_ = io_in[11] & ~_03958_;
	assign _03980_ = io_in[1] | ~io_in[3];
	assign _03992_ = _03980_ | io_in[4];
	assign _04003_ = _03992_ | io_in[8];
	assign _04014_ = _04003_ | io_in[9];
	assign _04025_ = _04014_ | io_in[10];
	assign _04036_ = _01985_ & ~_04025_;
	assign _04047_ = _00493_ | io_in[3];
	assign _04058_ = _04047_ | _03759_;
	assign _04069_ = _04058_ | _01208_;
	assign _04080_ = _06310_ & ~_04069_;
	assign _04091_ = _01430_ | io_in[3];
	assign _04103_ = _04091_ | _07422_;
	assign _04114_ = _04103_ | io_in[7];
	assign _04125_ = io_in[11] & ~_04114_;
	assign _04136_ = _00548_ | _03759_;
	assign _04147_ = _04136_ | io_in[7];
	assign _04158_ = _04147_ | io_in[8];
	assign _04169_ = _04158_ | io_in[9];
	assign _04180_ = io_in[10] & ~_04169_;
	assign _04191_ = _01430_ | _03759_;
	assign _04202_ = _04191_ | _02207_;
	assign _04214_ = _04202_ | io_in[8];
	assign _04225_ = _04214_ | io_in[10];
	assign _04236_ = _01985_ & ~_04225_;
	assign _04247_ = ~(io_in[1] & io_in[5]);
	assign _04258_ = _04247_ | io_in[6];
	assign _04269_ = _04258_ | _02207_;
	assign _04280_ = _04269_ | io_in[9];
	assign _04291_ = io_in[11] & ~_04280_;
	assign _04302_ = _06643_ | _07422_;
	assign _04313_ = _04302_ | _03759_;
	assign _04325_ = _04313_ | io_in[7];
	assign _04336_ = _01985_ & ~_04325_;
	assign _04347_ = _02206_ | _03759_;
	assign _04358_ = _04347_ | io_in[7];
	assign _04369_ = _04358_ | _01208_;
	assign _04380_ = _04369_ | io_in[9];
	assign _04391_ = _06310_ & ~_04380_;
	assign _04402_ = ~(io_in[3] & io_in[2]);
	assign _04413_ = _04402_ | io_in[6];
	assign _04424_ = _04413_ | io_in[8];
	assign _04436_ = _04424_ | _02096_;
	assign _04447_ = io_in[10] & ~_04436_;
	assign _04458_ = _02317_ | _01319_;
	assign _04469_ = _04458_ | io_in[5];
	assign _04480_ = _04469_ | io_in[6];
	assign _04491_ = _04480_ | _02207_;
	assign _04502_ = io_in[11] & ~_04491_;
	assign _04513_ = _01086_ | io_in[4];
	assign _04524_ = _04513_ | io_in[5];
	assign _04535_ = _04524_ | _02207_;
	assign _04547_ = _04535_ | _02096_;
	assign _04558_ = _04547_ | io_in[10];
	assign _04569_ = _01985_ & ~_04558_;
	assign _04580_ = _07198_ | _07422_;
	assign _04591_ = io_in[5] & ~_04580_;
	assign _04602_ = _03060_ | _03759_;
	assign _04613_ = _04602_ | io_in[8];
	assign _04624_ = _04613_ | io_in[9];
	assign _04635_ = io_in[10] & ~_04624_;
	assign _04646_ = _04136_ | _02207_;
	assign _04658_ = _04646_ | io_in[8];
	assign _04669_ = _04658_ | _02096_;
	assign _04680_ = io_in[10] & ~_04669_;
	assign _04691_ = _04103_ | _02207_;
	assign _04702_ = _04691_ | io_in[10];
	assign _04713_ = _01985_ & ~_04702_;
	assign _04724_ = _07499_ | _01208_;
	assign _04735_ = _04724_ | io_in[9];
	assign _04746_ = io_in[10] & ~_04735_;
	assign _04757_ = _02040_ | _01208_;
	assign _04769_ = _01985_ & ~_04757_;
	assign _04780_ = io_in[4] | ~io_in[2];
	assign _04791_ = _04780_ | io_in[5];
	assign _04802_ = _04791_ | io_in[6];
	assign _04813_ = _04802_ | _02207_;
	assign _04823_ = _04813_ | _01208_;
	assign _04834_ = _02096_ & ~_04823_;
	assign _04845_ = _03980_ | _07422_;
	assign _04856_ = _04845_ | io_in[7];
	assign _04867_ = _04856_ | io_in[8];
	assign _04879_ = _04867_ | io_in[9];
	assign _04890_ = io_in[11] & ~_04879_;
	assign _04901_ = _03736_ | _03759_;
	assign _04912_ = _04901_ | io_in[7];
	assign _04923_ = io_in[10] & ~_04912_;
	assign _04934_ = _00757_ | _03759_;
	assign _04945_ = _04934_ | _02207_;
	assign _04956_ = _04945_ | io_in[8];
	assign _04967_ = _06310_ & ~_04956_;
	assign _04978_ = _04047_ | _07422_;
	assign _04990_ = _04978_ | io_in[5];
	assign _05001_ = _04990_ | io_in[7];
	assign _05012_ = io_in[8] & ~_05001_;
	assign _05023_ = _01807_ | io_in[4];
	assign _05034_ = _05023_ | _03759_;
	assign _05045_ = _05034_ | _02207_;
	assign _05056_ = io_in[8] & ~_05045_;
	assign _05067_ = io_in[2] | io_in[4];
	assign _05078_ = _05067_ | _03759_;
	assign _05089_ = _05078_ | io_in[7];
	assign _05101_ = _05089_ | _01208_;
	assign _05112_ = _05101_ | io_in[9];
	assign _05123_ = _01985_ & ~_05112_;
	assign _05134_ = _03249_ | io_in[6];
	assign _05145_ = _05134_ | _02207_;
	assign _05156_ = _05145_ | io_in[8];
	assign _05167_ = _01985_ & ~_05156_;
	assign _05178_ = _04845_ | _03759_;
	assign _05189_ = _05178_ | _02207_;
	assign _05200_ = _05189_ | _01208_;
	assign _05212_ = _01985_ & ~_05200_;
	assign _05223_ = _02206_ | io_in[7];
	assign _05234_ = _05223_ | _01208_;
	assign _05245_ = _05234_ | io_in[9];
	assign _05256_ = _05245_ | io_in[10];
	assign _05267_ = io_in[11] & ~_05256_;
	assign _05278_ = _06643_ | _03759_;
	assign _05289_ = _05278_ | io_in[7];
	assign _05300_ = _05289_ | io_in[10];
	assign _05311_ = _01985_ & ~_05300_;
	assign _05323_ = _02383_ | io_in[6];
	assign _05334_ = _05323_ | _02096_;
	assign _05345_ = _01985_ & ~_05334_;
	assign _05356_ = _00043_ | _03759_;
	assign _05367_ = _05356_ | _02207_;
	assign _05378_ = _05367_ | _01208_;
	assign _05389_ = _05378_ | _06310_;
	assign _05400_ = _01985_ & ~_05389_;
	assign _05411_ = _07499_ | io_in[4];
	assign _05422_ = _05411_ | _03759_;
	assign _05434_ = _05422_ | _02207_;
	assign _05445_ = io_in[10] & ~_05434_;
	assign _05456_ = _03204_ | io_in[5];
	assign _05467_ = _05456_ | io_in[7];
	assign _05478_ = _01208_ & ~_05467_;
	assign _05489_ = _06532_ | io_in[4];
	assign _05500_ = _05489_ | io_in[5];
	assign _05511_ = _05500_ | io_in[6];
	assign _05522_ = _05511_ | _02207_;
	assign _05533_ = _05522_ | _02096_;
	assign _05545_ = _01985_ & ~_05533_;
	assign _05556_ = _05201_ | _02207_;
	assign _05567_ = _05556_ | _01208_;
	assign _05578_ = _05567_ | io_in[9];
	assign _05589_ = _05578_ | io_in[10];
	assign _05600_ = io_in[11] & ~_05589_;
	assign _05611_ = _04092_ | _02207_;
	assign _05622_ = _05611_ | _02096_;
	assign _05633_ = _05622_ | _06310_;
	assign _05644_ = _01985_ & ~_05633_;
	assign _05656_ = _05867_ | _01208_;
	assign _05667_ = _05656_ | io_in[9];
	assign _05678_ = io_in[10] & ~_05667_;
	assign _05689_ = _00394_ | io_in[8];
	assign _05700_ = io_in[11] & ~_05689_;
	assign _05711_ = _01241_ | io_in[7];
	assign _05722_ = _05711_ | io_in[10];
	assign _05733_ = io_in[11] & ~_05722_;
	assign _05744_ = _03992_ | io_in[6];
	assign _05755_ = _05744_ | io_in[7];
	assign _05767_ = _05755_ | _01208_;
	assign _05778_ = io_in[9] & ~_05767_;
	assign _05789_ = _00757_ | io_in[6];
	assign _05800_ = _05789_ | io_in[7];
	assign _05811_ = _05800_ | _02096_;
	assign _05822_ = io_in[11] & ~_05811_;
	assign _05833_ = _04402_ | io_in[5];
	assign _05844_ = _05833_ | io_in[6];
	assign _05855_ = _05844_ | _02207_;
	assign _05866_ = _05855_ | io_in[9];
	assign _05878_ = io_in[10] & ~_05866_;
	assign _05889_ = _01430_ | _07422_;
	assign _05900_ = _05889_ | _03759_;
	assign _05911_ = _05900_ | io_in[7];
	assign _05922_ = _05911_ | _02096_;
	assign _05933_ = io_in[11] & ~_05922_;
	assign _05944_ = _00273_ | _02207_;
	assign _05955_ = _05944_ | io_in[8];
	assign _05966_ = _01985_ & ~_05955_;
	assign _05977_ = _02672_ | io_in[3];
	assign _05989_ = _05977_ | _07422_;
	assign _06000_ = _05989_ | _02207_;
	assign _06011_ = _01985_ & ~_06000_;
	assign _06022_ = _06643_ | io_in[6];
	assign _06032_ = _06022_ | _02207_;
	assign _06043_ = _06032_ | _06310_;
	assign _06054_ = _01985_ & ~_06043_;
	assign _06065_ = _01307_ | io_in[6];
	assign _06076_ = _06065_ | io_in[8];
	assign _06087_ = io_in[9] & ~_06076_;
	assign _06099_ = _01485_ | _02207_;
	assign _06110_ = _06099_ | _02096_;
	assign _06121_ = _06310_ & ~_06110_;
	assign _06132_ = _03149_ | _03759_;
	assign _06143_ = _06132_ | _02207_;
	assign _06154_ = _06143_ | io_in[9];
	assign _06165_ = io_in[11] & ~_06154_;
	assign _06176_ = _01962_ | io_in[5];
	assign _06187_ = _06176_ | _03759_;
	assign _06198_ = _06187_ | io_in[8];
	assign _06210_ = _06198_ | io_in[9];
	assign _06221_ = _06210_ | io_in[10];
	assign _06232_ = _01985_ & ~_06221_;
	assign _06243_ = _03981_ | _07422_;
	assign _06254_ = _06243_ | _03759_;
	assign _06265_ = _06254_ | io_in[9];
	assign _06276_ = _06310_ & ~_06265_;
	assign _06287_ = _05067_ | io_in[6];
	assign _06298_ = _06287_ | _02207_;
	assign _06309_ = _06298_ | io_in[8];
	assign _06321_ = _06309_ | io_in[9];
	assign _06332_ = _06321_ | io_in[10];
	assign _06343_ = io_in[11] & ~_06332_;
	assign _06354_ = _00669_ | io_in[6];
	assign _06365_ = _06354_ | _02207_;
	assign _06376_ = _06365_ | _02096_;
	assign _06387_ = _06376_ | _06310_;
	assign _06398_ = _01985_ & ~_06387_;
	assign _06409_ = _02860_ | _01208_;
	assign _06420_ = _06409_ | io_in[10];
	assign _06432_ = _01985_ & ~_06420_;
	assign _06443_ = io_in[4] | ~io_in[1];
	assign _06454_ = _06443_ | io_in[5];
	assign _06465_ = _06454_ | _03759_;
	assign _06476_ = _06465_ | io_in[8];
	assign _06487_ = _06476_ | io_in[9];
	assign _06498_ = io_in[11] & ~_06487_;
	assign _06509_ = _00548_ | io_in[3];
	assign _06520_ = _06509_ | _07422_;
	assign _06531_ = _06520_ | io_in[7];
	assign _06543_ = _06531_ | io_in[9];
	assign _06554_ = _01985_ & ~_06543_;
	assign _06565_ = _00548_ | io_in[6];
	assign _06576_ = _06565_ | io_in[7];
	assign _06587_ = _06576_ | _02096_;
	assign _06598_ = _01985_ & ~_06587_;
	assign _06609_ = _07444_ | _03094_;
	assign _06620_ = _06609_ | _03759_;
	assign _06631_ = io_in[10] & ~_06620_;
	assign _06642_ = _03205_ | io_in[4];
	assign _06654_ = _06642_ | io_in[5];
	assign _06665_ = _06654_ | io_in[6];
	assign _06676_ = _06665_ | io_in[7];
	assign _06687_ = _06676_ | _01208_;
	assign _06698_ = _06687_ | _02096_;
	assign _06709_ = _01985_ & ~_06698_;
	assign _06720_ = _07246_ | _07422_;
	assign _06731_ = _06720_ | io_in[7];
	assign _06742_ = _06731_ | io_in[9];
	assign _06753_ = _06310_ & ~_06742_;
	assign _06765_ = _02971_ | io_in[5];
	assign _06776_ = _06765_ | _03759_;
	assign _06787_ = _06776_ | _02207_;
	assign _06798_ = _06787_ | _01208_;
	assign _06809_ = _01985_ & ~_06798_;
	assign _06820_ = _05977_ | _01208_;
	assign _06831_ = _06820_ | _06310_;
	assign _06842_ = _01985_ & ~_06831_;
	assign _06853_ = _02317_ | _06421_;
	assign _06864_ = _06853_ | _01319_;
	assign _06876_ = _06864_ | io_in[8];
	assign _06887_ = io_in[11] & ~_06876_;
	assign _06898_ = _02394_ | _01208_;
	assign _06909_ = _06898_ | _02096_;
	assign _06920_ = _01985_ & ~_06909_;
	assign _06931_ = _02428_ | io_in[3];
	assign _06942_ = _06931_ | _03094_;
	assign _06953_ = _06942_ | _02207_;
	assign _06964_ = io_in[11] & ~_06953_;
	assign _06975_ = ~(io_in[1] & io_in[4]);
	assign _06987_ = _06975_ | io_in[7];
	assign _06998_ = _06987_ | io_in[8];
	assign _07009_ = _06998_ | io_in[9];
	assign _07020_ = io_in[10] & ~_07009_;
	assign _07031_ = _00548_ | _07422_;
	assign _07042_ = _07031_ | io_in[7];
	assign _07053_ = _07042_ | io_in[8];
	assign _07064_ = io_in[10] & ~_07053_;
	assign _07075_ = _03149_ | _07422_;
	assign _07086_ = _07075_ | _03759_;
	assign _07098_ = _07086_ | io_in[7];
	assign _07109_ = _01985_ & ~_07098_;
	assign _07120_ = _00768_ | _02207_;
	assign _07131_ = _06310_ & ~_07120_;
	assign _07142_ = _01596_ | _07422_;
	assign _07153_ = _07142_ | _03759_;
	assign _07164_ = _07153_ | io_in[9];
	assign _07175_ = io_in[11] & ~_07164_;
	assign _07186_ = _00317_ | _07422_;
	assign _07197_ = _07186_ | _01208_;
	assign _07209_ = _07197_ | io_in[10];
	assign _07220_ = io_in[11] & ~_07209_;
	assign _07231_ = _03149_ | io_in[6];
	assign _07239_ = _07231_ | io_in[7];
	assign _07240_ = _07239_ | _01208_;
	assign _07241_ = io_in[11] & ~_07240_;
	assign _07242_ = _06654_ | _03759_;
	assign _07243_ = _07242_ | _02207_;
	assign _07244_ = _07243_ | _06310_;
	assign _07245_ = io_in[11] & ~_07244_;
	assign _07247_ = _03892_ | io_in[6];
	assign _07248_ = _07247_ | io_in[7];
	assign _07249_ = io_in[11] & ~_07248_;
	assign _07250_ = _07367_ | _07422_;
	assign _07251_ = _07250_ | _03759_;
	assign _07252_ = _07251_ | io_in[7];
	assign _07253_ = _07252_ | _01208_;
	assign _07254_ = io_in[9] & ~_07253_;
	assign _07255_ = _06931_ | io_in[4];
	assign _07256_ = _07255_ | io_in[7];
	assign _07258_ = _01208_ & ~_07256_;
	assign _07259_ = _07356_ | io_in[4];
	assign _07260_ = _07259_ | io_in[6];
	assign _07261_ = _07260_ | io_in[7];
	assign _07262_ = _07261_ | _01208_;
	assign _07263_ = io_in[10] & ~_07262_;
	assign _07264_ = _01430_ | io_in[4];
	assign _07265_ = _07264_ | io_in[7];
	assign _07266_ = _07265_ | _01208_;
	assign _07267_ = _07266_ | io_in[9];
	assign _07269_ = io_in[10] & ~_07267_;
	assign _07270_ = _03149_ | io_in[4];
	assign _07271_ = _07270_ | io_in[5];
	assign _07272_ = _07271_ | _02207_;
	assign _07273_ = io_in[9] & ~_07272_;
	assign _07274_ = _03781_ | io_in[6];
	assign _07275_ = _07274_ | _02207_;
	assign _07276_ = _07275_ | _01208_;
	assign _07277_ = _02096_ & ~_07276_;
	assign _07278_ = _07259_ | _03759_;
	assign _07280_ = _07278_ | io_in[7];
	assign _07281_ = _07280_ | io_in[10];
	assign _07282_ = io_in[11] & ~_07281_;
	assign _07283_ = _04402_ | io_in[4];
	assign _07284_ = _07283_ | _03759_;
	assign _07285_ = _07284_ | io_in[7];
	assign _07286_ = _07285_ | _01208_;
	assign _07287_ = _07286_ | _06310_;
	assign _07288_ = _01985_ & ~_07287_;
	assign _07289_ = _01962_ | _07422_;
	assign _07291_ = _07289_ | io_in[5];
	assign _07292_ = _07291_ | io_in[6];
	assign _07293_ = _07292_ | _02207_;
	assign _07294_ = _07293_ | _01208_;
	assign _07295_ = io_in[9] & ~_07294_;
	assign _07296_ = _02428_ | _01208_;
	assign _07297_ = _07296_ | _02096_;
	assign _07298_ = _07297_ | _06310_;
	assign _07299_ = _01985_ & ~_07298_;
	assign _07300_ = _03870_ | _01319_;
	assign _07302_ = _07300_ | io_in[4];
	assign _07303_ = _07302_ | io_in[6];
	assign _07304_ = _07303_ | _02207_;
	assign _07305_ = _06310_ & ~_07304_;
	assign _07306_ = _02727_ | io_in[5];
	assign _07307_ = _07306_ | _03759_;
	assign _07308_ = _07307_ | _02207_;
	assign _07309_ = _07308_ | io_in[8];
	assign _07310_ = _02096_ & ~_07309_;
	assign _07311_ = _06520_ | io_in[6];
	assign _07313_ = _07311_ | io_in[7];
	assign _07314_ = _02096_ & ~_07313_;
	assign _07315_ = _03160_ | io_in[8];
	assign _07316_ = _07315_ | io_in[9];
	assign _07317_ = io_in[10] & ~_07316_;
	assign _07318_ = _07433_ | _07422_;
	assign _07319_ = _07318_ | _03759_;
	assign _07320_ = _07319_ | _02096_;
	assign _07321_ = _06310_ & ~_07320_;
	assign _07322_ = _02218_ | _02207_;
	assign _07324_ = _07322_ | io_in[8];
	assign _07325_ = _07324_ | _02096_;
	assign _07326_ = _06310_ & ~_07325_;
	assign _07327_ = _06642_ | _02207_;
	assign _07328_ = _07327_ | io_in[8];
	assign _07329_ = io_in[10] & ~_07328_;
	assign _07330_ = _00043_ | _03094_;
	assign _07331_ = _07330_ | _03759_;
	assign _07332_ = _07331_ | _01208_;
	assign _07333_ = _06310_ & ~_07332_;
	assign _07335_ = _00482_ | _01319_;
	assign _07336_ = _07335_ | _07422_;
	assign _07337_ = _07336_ | _01208_;
	assign _07338_ = _07337_ | _02096_;
	assign _07339_ = _01985_ & ~_07338_;
	assign _07340_ = _03404_ | _02207_;
	assign _07341_ = _07340_ | _01208_;
	assign _07342_ = _02096_ & ~_07341_;
	assign _07343_ = _03304_ | io_in[6];
	assign _07344_ = _07343_ | io_in[7];
	assign _07346_ = _07344_ | _01208_;
	assign _07347_ = _06310_ & ~_07346_;
	assign _07348_ = _07257_ | _02207_;
	assign _07349_ = _07348_ | io_in[8];
	assign _07350_ = _06310_ & ~_07349_;
	assign _07351_ = _06509_ | io_in[4];
	assign _07352_ = _07351_ | io_in[5];
	assign _07353_ = _07352_ | _03759_;
	assign _07354_ = _07353_ | _02096_;
	assign _07355_ = _07354_ | io_in[10];
	assign _07357_ = _01985_ & ~_07355_;
	assign _07358_ = _02672_ | _07422_;
	assign _07359_ = _07358_ | _02207_;
	assign _07360_ = _07359_ | io_in[8];
	assign _07361_ = _02096_ & ~_07360_;
	assign _07362_ = _02971_ | io_in[4];
	assign _07363_ = _07362_ | _02207_;
	assign _07364_ = _07363_ | io_in[8];
	assign _07365_ = _07364_ | io_in[9];
	assign _07366_ = _01985_ & ~_07365_;
	assign _07368_ = ~(io_in[2] & io_in[4]);
	assign _07369_ = _07368_ | _03759_;
	assign _07370_ = _07369_ | io_in[7];
	assign _07371_ = _07370_ | io_in[8];
	assign _07372_ = io_in[9] & ~_07371_;
	assign _07373_ = _07455_ | io_in[7];
	assign _07374_ = _07373_ | io_in[9];
	assign _07375_ = io_in[10] & ~_07374_;
	assign _07376_ = _00174_ | io_in[6];
	assign _07377_ = _07376_ | _02096_;
	assign _07379_ = io_in[11] & ~_07377_;
	assign _07380_ = _03404_ | io_in[6];
	assign _07381_ = _07380_ | _01208_;
	assign _07382_ = io_in[11] & ~_07381_;
	assign _07383_ = _04402_ | _07422_;
	assign _07384_ = _07383_ | io_in[8];
	assign _07385_ = _07384_ | _02096_;
	assign _07386_ = io_in[10] & ~_07385_;
	assign _07387_ = _01086_ | io_in[7];
	assign _07388_ = _07387_ | io_in[8];
	assign _07390_ = _07388_ | _02096_;
	assign _07391_ = io_in[10] & ~_07390_;
	assign _07392_ = _07300_ | _07422_;
	assign _07393_ = _07392_ | io_in[7];
	assign _07394_ = _07393_ | _06310_;
	assign _07395_ = io_in[11] & ~_07394_;
	assign _07396_ = _06565_ | _02207_;
	assign _07397_ = _07396_ | _06310_;
	assign _07398_ = io_in[11] & ~_07397_;
	assign _07399_ = _04114_ | io_in[9];
	assign _07401_ = _06310_ & ~_07399_;
	assign _07402_ = _03304_ | io_in[4];
	assign _07403_ = _07402_ | io_in[6];
	assign _07404_ = io_in[11] & ~_07403_;
	assign _07405_ = _05201_ | io_in[7];
	assign _07406_ = _07405_ | _01208_;
	assign _07407_ = _07406_ | io_in[9];
	assign _07408_ = _07407_ | io_in[10];
	assign _07409_ = _01985_ & ~_07408_;
	assign _07410_ = _02428_ | _01319_;
	assign _07412_ = _07410_ | _07422_;
	assign _07413_ = _07412_ | _03759_;
	assign _07414_ = _07413_ | io_in[8];
	assign _07415_ = _01985_ & ~_07414_;
	assign _07416_ = _05889_ | io_in[6];
	assign _07417_ = _07416_ | io_in[8];
	assign _07418_ = _02096_ & ~_07417_;
	assign _07419_ = _05977_ | io_in[4];
	assign _07420_ = _07419_ | io_in[7];
	assign _07421_ = _02096_ & ~_07420_;
	assign _07423_ = _04758_ | io_in[7];
	assign _07424_ = _07423_ | _01208_;
	assign _07425_ = _07424_ | io_in[9];
	assign _07426_ = io_in[11] & ~_07425_;
	assign _07427_ = _07358_ | io_in[5];
	assign _07428_ = _07427_ | io_in[6];
	assign _07429_ = _07428_ | _01208_;
	assign _07430_ = io_in[9] & ~_07429_;
	assign _07431_ = _03304_ | _02207_;
	assign _07432_ = _07431_ | io_in[8];
	assign _07434_ = io_in[11] & ~_07432_;
	assign _07435_ = _05977_ | io_in[5];
	assign _07436_ = _07435_ | io_in[6];
	assign _07437_ = io_in[8] & ~_07436_;
	assign _07438_ = _03249_ | _03759_;
	assign _07439_ = _07438_ | io_in[8];
	assign _07440_ = _02096_ & ~_07439_;
	assign _07441_ = io_in[5] & ~_02029_;
	assign _07442_ = _07441_ | _07440_;
	assign _07443_ = _07442_ | _07437_;
	assign _07445_ = _07443_ | _07434_;
	assign _07446_ = _07445_ | _07430_;
	assign _07447_ = _07446_ | _07426_;
	assign _07448_ = _07447_ | _07421_;
	assign _07449_ = _07448_ | _07418_;
	assign _07450_ = _07449_ | _07415_;
	assign _07451_ = _07450_ | _07409_;
	assign _07452_ = _07451_ | _07404_;
	assign _07453_ = _07452_ | _07401_;
	assign _07454_ = _07453_ | _07398_;
	assign _07456_ = _07454_ | _07395_;
	assign _07457_ = _07456_ | _07391_;
	assign _07458_ = _07457_ | _07386_;
	assign _07459_ = _07458_ | _07382_;
	assign _07460_ = _07459_ | _07379_;
	assign _07461_ = _07460_ | _07375_;
	assign _07462_ = _07461_ | _07372_;
	assign _07463_ = _07462_ | _07366_;
	assign _07464_ = _07463_ | _07361_;
	assign _07465_ = _07464_ | _07357_;
	assign _07467_ = _07465_ | _07350_;
	assign _07468_ = _07467_ | _07347_;
	assign _07469_ = _07468_ | _07342_;
	assign _07470_ = _07469_ | _07339_;
	assign _07471_ = _07470_ | _07333_;
	assign _07472_ = _07471_ | _07329_;
	assign _07473_ = _07472_ | _07326_;
	assign _07474_ = _07473_ | _07321_;
	assign _07475_ = _07474_ | _07317_;
	assign _07476_ = _07475_ | _07314_;
	assign _07478_ = _07476_ | _07310_;
	assign _07479_ = _07478_ | _07305_;
	assign _07480_ = _07479_ | _07299_;
	assign _07481_ = _07480_ | _07295_;
	assign _07482_ = _07481_ | _07288_;
	assign _07483_ = _07482_ | _07282_;
	assign _07484_ = _07483_ | _07277_;
	assign _07485_ = _07484_ | _07273_;
	assign _07486_ = _07485_ | _07269_;
	assign _07487_ = _07486_ | _07263_;
	assign _07489_ = _07487_ | _07258_;
	assign _07490_ = _07489_ | _07254_;
	assign _07491_ = _07490_ | _07249_;
	assign _07492_ = _07491_ | _07245_;
	assign _07493_ = _07492_ | _07241_;
	assign _07494_ = _07493_ | _07220_;
	assign _07495_ = _07494_ | _07175_;
	assign _07496_ = _07495_ | _07131_;
	assign _07497_ = _07496_ | _07109_;
	assign _07498_ = _07497_ | _07064_;
	assign _07500_ = _07498_ | _07020_;
	assign _07501_ = _07500_ | _06964_;
	assign _07502_ = _07501_ | _06920_;
	assign _07503_ = _07502_ | _06887_;
	assign _07504_ = _07503_ | _06842_;
	assign _07505_ = _07504_ | _06809_;
	assign _07506_ = _07505_ | _06753_;
	assign _07507_ = _07506_ | _06709_;
	assign _07508_ = _07507_ | _06631_;
	assign _07509_ = _07508_ | _06598_;
	assign _00000_ = _07509_ | _06554_;
	assign _00001_ = _00000_ | _06498_;
	assign _00002_ = _00001_ | _06432_;
	assign _00003_ = _00002_ | _06398_;
	assign _00004_ = _00003_ | _06343_;
	assign _00005_ = _00004_ | _06276_;
	assign _00006_ = _00005_ | _06232_;
	assign _00007_ = _00006_ | _06165_;
	assign _00008_ = _00007_ | _06121_;
	assign _00009_ = _00008_ | _06087_;
	assign _00011_ = _00009_ | _06054_;
	assign _00012_ = _00011_ | _06011_;
	assign _00013_ = _00012_ | _05966_;
	assign _00014_ = _00013_ | _05933_;
	assign _00015_ = _00014_ | _05878_;
	assign _00016_ = _00015_ | _05822_;
	assign _00017_ = _00016_ | _05778_;
	assign _00018_ = _00017_ | _05733_;
	assign _00019_ = _00018_ | _05700_;
	assign _00020_ = _00019_ | _05678_;
	assign _00022_ = _00020_ | _05644_;
	assign _00023_ = _00022_ | _05600_;
	assign _00024_ = _00023_ | _05545_;
	assign _00025_ = _00024_ | _05478_;
	assign _00026_ = _00025_ | _05445_;
	assign _00027_ = _00026_ | _05400_;
	assign _00028_ = _00027_ | _05345_;
	assign _00029_ = _00028_ | _05311_;
	assign _00030_ = _00029_ | _05267_;
	assign _00031_ = _00030_ | _05212_;
	assign _00033_ = _00031_ | _05167_;
	assign _00034_ = _00033_ | _05123_;
	assign _00035_ = _00034_ | _05056_;
	assign _00036_ = _00035_ | _05012_;
	assign _00037_ = _00036_ | _04967_;
	assign _00038_ = _00037_ | _04923_;
	assign _00039_ = _00038_ | _04890_;
	assign _00040_ = _00039_ | _04834_;
	assign _00041_ = _00040_ | _04769_;
	assign _00042_ = _00041_ | _04746_;
	assign _00044_ = _00042_ | _04713_;
	assign _00045_ = _00044_ | _04680_;
	assign _00046_ = _00045_ | _04635_;
	assign _00047_ = _00046_ | _04591_;
	assign _00048_ = _00047_ | _04569_;
	assign _00049_ = _00048_ | _04502_;
	assign _00050_ = _00049_ | _04447_;
	assign _00051_ = _00050_ | _04391_;
	assign _00052_ = _00051_ | _04336_;
	assign _00053_ = _00052_ | _04291_;
	assign _00055_ = _00053_ | _04236_;
	assign _00056_ = _00055_ | _04180_;
	assign _00057_ = _00056_ | _04125_;
	assign _00058_ = _00057_ | _04080_;
	assign _00059_ = _00058_ | _04036_;
	assign _00060_ = _00059_ | _03969_;
	assign _00061_ = _00060_ | _03925_;
	assign _00062_ = _00061_ | _03869_;
	assign _00063_ = _00062_ | _03814_;
	assign _00064_ = _00063_ | _03770_;
	assign _00066_ = _00064_ | _03714_;
	assign _00067_ = _00066_ | _03670_;
	assign _00068_ = _00067_ | _03636_;
	assign _00069_ = _00068_ | _03581_;
	assign _00070_ = _00069_ | _03515_;
	assign _00071_ = _00070_ | _03482_;
	assign _00072_ = _00071_ | _03449_;
	assign _00073_ = _00072_ | _03393_;
	assign _00074_ = _00073_ | _03349_;
	assign _00075_ = _00074_ | _03293_;
	assign _00077_ = _00075_ | _03238_;
	assign _00078_ = _00077_ | _03193_;
	assign _00079_ = _00078_ | _03138_;
	assign _00080_ = _00079_ | _03105_;
	assign _00081_ = _00080_ | _03049_;
	assign _00082_ = _00081_ | _03016_;
	assign _00083_ = _00082_ | _02960_;
	assign _00084_ = _00083_ | _02905_;
	assign _00085_ = _00084_ | _02849_;
	assign _00086_ = _00085_ | _02805_;
	assign _00088_ = _00086_ | _02760_;
	assign _00089_ = _00088_ | _02716_;
	assign _00090_ = _00089_ | _02661_;
	assign _00091_ = _00090_ | _02627_;
	assign _00092_ = _00091_ | _02550_;
	assign _00093_ = _00092_ | _02494_;
	assign _00094_ = _00093_ | _02461_;
	assign _00095_ = _00094_ | _02416_;
	assign _00096_ = _00095_ | _02372_;
	assign _00097_ = _00096_ | _02339_;
	assign _00099_ = _00097_ | _02294_;
	assign _00100_ = _00099_ | _02262_;
	assign _00101_ = _00100_ | _02195_;
	assign _00102_ = _00101_ | _02151_;
	assign _00103_ = _00102_ | _02095_;
	assign _00104_ = _00103_ | _02062_;
	assign _00105_ = _00104_ | _02007_;
	assign _00106_ = _00105_ | _01951_;
	assign _00107_ = _00106_ | _01896_;
	assign _00108_ = _00107_ | _01862_;
	assign _00110_ = _00108_ | _01796_;
	assign _00111_ = _00110_ | _01751_;
	assign _00112_ = _00111_ | _01718_;
	assign _00113_ = _00112_ | _01674_;
	assign _00114_ = _00113_ | _01640_;
	assign _00115_ = _00114_ | _01585_;
	assign _00116_ = _00115_ | _01529_;
	assign _00117_ = _00116_ | _01474_;
	assign _00118_ = _00117_ | _01418_;
	assign _00119_ = _00118_ | _01341_;
	assign _00121_ = _00119_ | _01285_;
	assign _00122_ = _00121_ | _01207_;
	assign _00123_ = _00122_ | _01141_;
	assign _00124_ = _00123_ | _01075_;
	assign _00125_ = _00124_ | _01020_;
	assign _00126_ = _00125_ | _00976_;
	assign _00127_ = _00126_ | _00922_;
	assign _00128_ = _00127_ | _00867_;
	assign _00129_ = _00128_ | _00801_;
	assign _00130_ = _00129_ | _00746_;
	assign _00132_ = _00130_ | _00713_;
	assign _00133_ = _00132_ | _00647_;
	assign _00134_ = _00133_ | _00603_;
	assign _00135_ = _05989_ | io_in[6];
	assign _00136_ = _00134_ | ~_00135_;
	assign _00137_ = _00136_ | _00537_;
	assign _00138_ = _00137_ | _00471_;
	assign _00139_ = _00138_ | _00427_;
	assign _00140_ = _00139_ | _00372_;
	assign _00141_ = _00140_ | _00306_;
	assign _00143_ = _00141_ | _00262_;
	assign _00144_ = _00143_ | _00207_;
	assign _00145_ = _00144_ | _00163_;
	assign _00146_ = _00145_ | _00109_;
	assign _00147_ = _00146_ | _00032_;
	assign _00148_ = _00147_ | _07488_;
	assign _00149_ = _00148_ | _07411_;
	assign _00150_ = _00149_ | _07345_;
	assign _00151_ = _00150_ | _07290_;
	assign _00152_ = _00151_ | _07087_;
	assign _00154_ = _00152_ | _06199_;
	assign _00155_ = _00154_ | _05756_;
	assign _00156_ = _00155_ | _05090_;
	assign _00157_ = _00156_ | _04536_;
	assign _00158_ = _00157_ | _03648_;
	assign _00159_ = _00158_ | _02983_;
	assign \mchip.val [6] = _00159_ | _01874_;
	assign _00160_ = io_in[6] | ~io_in[0];
	assign _00161_ = _00160_ | _02207_;
	assign _00162_ = _00161_ | io_in[8];
	assign _00164_ = _00162_ | _02096_;
	assign _00165_ = _01985_ & ~_00164_;
	assign _00166_ = _03249_ | _07422_;
	assign _00167_ = _00166_ | _02096_;
	assign _00168_ = io_in[11] & ~_00167_;
	assign _00169_ = _00166_ | io_in[6];
	assign _00170_ = _00169_ | _02207_;
	assign _00171_ = _00170_ | io_in[8];
	assign _00172_ = io_in[9] & ~_00171_;
	assign _00173_ = _03870_ | _07422_;
	assign _00175_ = _00173_ | io_in[6];
	assign _00176_ = _00175_ | io_in[10];
	assign _00177_ = _01985_ & ~_00176_;
	assign _00178_ = _03870_ | _03094_;
	assign _00179_ = _00178_ | _02096_;
	assign _00180_ = io_in[11] & ~_00179_;
	assign _00181_ = io_in[10] & ~_04114_;
	assign _00182_ = _07356_ | io_in[5];
	assign _00183_ = _00182_ | io_in[7];
	assign _00184_ = _00183_ | io_in[8];
	assign _00186_ = _02096_ & ~_00184_;
	assign _00187_ = io_in[6] | ~io_in[2];
	assign _00188_ = _00187_ | io_in[7];
	assign _00189_ = _00188_ | _01208_;
	assign _00190_ = _00189_ | io_in[9];
	assign _00191_ = io_in[10] & ~_00190_;
	assign _00192_ = _04091_ | io_in[5];
	assign _00193_ = _00192_ | io_in[6];
	assign _00194_ = _00193_ | _01208_;
	assign _00195_ = _02096_ & ~_00194_;
	assign _00197_ = io_in[10] & ~_05467_;
	assign _00198_ = _01296_ | io_in[4];
	assign _00199_ = _00198_ | _02207_;
	assign _00200_ = _00199_ | io_in[8];
	assign _00201_ = io_in[10] & ~_00200_;
	assign _00202_ = io_in[0] | ~io_in[4];
	assign _00203_ = _00202_ | io_in[6];
	assign _00204_ = _00203_ | _02207_;
	assign _00205_ = _00204_ | io_in[8];
	assign _00206_ = _00205_ | io_in[9];
	assign _00208_ = _06310_ & ~_00206_;
	assign _00209_ = _01430_ | io_in[5];
	assign _00210_ = _00209_ | io_in[6];
	assign _00211_ = _00210_ | io_in[7];
	assign _00212_ = _00211_ | _01208_;
	assign _00213_ = io_in[10] & ~_00212_;
	assign _00214_ = _07367_ | _03759_;
	assign _00215_ = _00214_ | _01208_;
	assign _00216_ = io_in[9] & ~_00215_;
	assign _00217_ = _00182_ | io_in[6];
	assign _00219_ = _00217_ | _02207_;
	assign _00220_ = io_in[9] & ~_00219_;
	assign _00221_ = io_in[5] | ~io_in[0];
	assign _00222_ = _00221_ | _03759_;
	assign _00223_ = _00222_ | _02207_;
	assign _00224_ = _00223_ | io_in[8];
	assign _00225_ = _00224_ | io_in[9];
	assign _00226_ = io_in[11] & ~_00225_;
	assign _00227_ = _07300_ | _03759_;
	assign _00228_ = _00227_ | io_in[8];
	assign _00230_ = _00228_ | io_in[10];
	assign _00231_ = _01985_ & ~_00230_;
	assign _00232_ = _00823_ | io_in[6];
	assign _00233_ = _00232_ | io_in[7];
	assign _00234_ = io_in[8] & ~_00233_;
	assign _00235_ = _00933_ | io_in[5];
	assign _00236_ = _00235_ | io_in[7];
	assign _00237_ = _00236_ | _02096_;
	assign _00238_ = io_in[11] & ~_00237_;
	assign _00239_ = _02206_ | _03094_;
	assign _00241_ = _00239_ | io_in[6];
	assign _00242_ = _00241_ | _02207_;
	assign _00243_ = _00242_ | _01208_;
	assign _00244_ = io_in[9] & ~_00243_;
	assign _00245_ = _07246_ | io_in[3];
	assign _00246_ = _00245_ | _07422_;
	assign _00247_ = _00246_ | io_in[7];
	assign _00248_ = io_in[10] & ~_00247_;
	assign _00249_ = _01985_ & ~_03537_;
	assign _00250_ = _02505_ | _07422_;
	assign _00252_ = _00250_ | _01208_;
	assign _00253_ = _06310_ & ~_00252_;
	assign _00254_ = _00878_ | io_in[5];
	assign _00255_ = _00254_ | _03759_;
	assign _00256_ = _00255_ | _02096_;
	assign _00257_ = _06310_ & ~_00256_;
	assign _00258_ = _04780_ | _03759_;
	assign _00259_ = _00258_ | io_in[7];
	assign _00260_ = _00259_ | _01208_;
	assign _00261_ = _00260_ | io_in[9];
	assign _00263_ = _06310_ & ~_00261_;
	assign _00264_ = _05977_ | io_in[6];
	assign _00265_ = _00264_ | _02207_;
	assign _00266_ = _01985_ & ~_00265_;
	assign _00267_ = _01352_ | _07422_;
	assign _00268_ = _00267_ | _01208_;
	assign _00269_ = _00268_ | io_in[9];
	assign _00270_ = _06310_ & ~_00269_;
	assign _00271_ = _00178_ | io_in[6];
	assign _00272_ = io_in[9] & ~_00271_;
	assign _00274_ = _04047_ | io_in[4];
	assign _00275_ = io_in[11] & ~_00274_;
	assign _00276_ = _00328_ | io_in[6];
	assign _00277_ = _00276_ | io_in[8];
	assign _00278_ = _06310_ & ~_00277_;
	assign _00279_ = _07231_ | _02096_;
	assign _00280_ = _06310_ & ~_00279_;
	assign _00281_ = _00812_ | _07422_;
	assign _00282_ = _00281_ | _01208_;
	assign _00283_ = _00282_ | _02096_;
	assign _00285_ = _01985_ & ~_00283_;
	assign _00286_ = _06864_ | io_in[5];
	assign _00287_ = _00286_ | io_in[6];
	assign _00288_ = _01985_ & ~_00287_;
	assign _00289_ = _00173_ | io_in[7];
	assign _00290_ = _00289_ | io_in[8];
	assign _00291_ = _01985_ & ~_00290_;
	assign _00292_ = _07367_ | io_in[5];
	assign _00293_ = _00292_ | io_in[8];
	assign _00294_ = _00293_ | io_in[9];
	assign _00296_ = _06310_ & ~_00294_;
	assign _00297_ = io_in[5] | io_in[2];
	assign _00298_ = _00297_ | _03759_;
	assign _00299_ = _00298_ | io_in[7];
	assign _00300_ = _00299_ | _01208_;
	assign _00301_ = _00300_ | _02096_;
	assign _00302_ = _00301_ | _06310_;
	assign _00303_ = io_in[11] & ~_00302_;
	assign _00304_ = _00198_ | _03759_;
	assign _00305_ = io_in[11] & ~_00304_;
	assign _00307_ = io_in[4] | ~io_in[0];
	assign _00308_ = _00307_ | io_in[6];
	assign _00309_ = _00308_ | _02207_;
	assign _00310_ = _00309_ | io_in[8];
	assign _00311_ = _00310_ | io_in[9];
	assign _00312_ = io_in[11] & ~_00311_;
	assign _00313_ = _06642_ | io_in[7];
	assign _00314_ = _00313_ | _06310_;
	assign _00315_ = io_in[11] & ~_00314_;
	assign _00316_ = _02107_ | _03759_;
	assign _00318_ = _00316_ | io_in[7];
	assign _00319_ = _00318_ | io_in[8];
	assign _00320_ = _06310_ & ~_00319_;
	assign _00321_ = ~(io_in[0] & io_in[4]);
	assign _00322_ = _00321_ | _02207_;
	assign _00323_ = _00322_ | _01208_;
	assign _00324_ = io_in[11] & ~_00323_;
	assign _00325_ = _01962_ | _03094_;
	assign _00326_ = _00325_ | _03759_;
	assign _00327_ = _02207_ & ~_00326_;
	assign _00329_ = _03892_ | _03759_;
	assign _00330_ = _00329_ | _02096_;
	assign _00331_ = _00330_ | _06310_;
	assign _00332_ = _01985_ & ~_00331_;
	assign _00333_ = _00383_ | io_in[6];
	assign _00334_ = _00333_ | io_in[7];
	assign _00335_ = io_in[11] & ~_00334_;
	assign _00336_ = _07433_ | io_in[5];
	assign _00337_ = _00336_ | io_in[7];
	assign _00338_ = _00337_ | _02096_;
	assign _00340_ = io_in[11] & ~_00338_;
	assign _00341_ = _07396_ | _01208_;
	assign _00342_ = _06310_ & ~_00341_;
	assign _00343_ = _00173_ | io_in[9];
	assign _00344_ = _01985_ & ~_00343_;
	assign _00345_ = _07270_ | io_in[6];
	assign _00346_ = _01208_ & ~_00345_;
	assign _00347_ = _00307_ | io_in[5];
	assign _00348_ = _00347_ | io_in[6];
	assign _00349_ = _00348_ | _02096_;
	assign _00351_ = _00349_ | io_in[10];
	assign _00352_ = _01985_ & ~_00351_;
	assign _00353_ = _00286_ | io_in[7];
	assign _00354_ = io_in[9] & ~_00353_;
	assign _00355_ = _07318_ | _02207_;
	assign _00356_ = _00355_ | io_in[10];
	assign _00357_ = io_in[11] & ~_00356_;
	assign _00358_ = _04524_ | _02096_;
	assign _00359_ = io_in[11] & ~_00358_;
	assign _00360_ = _06853_ | _07422_;
	assign _00362_ = _00360_ | _01208_;
	assign _00363_ = io_in[11] & ~_00362_;
	assign _00364_ = _00174_ | io_in[8];
	assign _00365_ = _06310_ & ~_00364_;
	assign _00366_ = _00173_ | _06310_;
	assign _00367_ = io_in[11] & ~_00366_;
	assign _00368_ = _02206_ | _07422_;
	assign _00369_ = _00368_ | io_in[8];
	assign _00370_ = _00369_ | _02096_;
	assign _00371_ = io_in[10] & ~_00370_;
	assign _00373_ = _00120_ | _03094_;
	assign _00374_ = _00373_ | _03759_;
	assign _00375_ = _00374_ | _02207_;
	assign _00376_ = _01985_ & ~_00375_;
	assign _00377_ = _00317_ | io_in[7];
	assign _00378_ = _00377_ | io_in[9];
	assign _00379_ = _00378_ | io_in[10];
	assign _00380_ = _01985_ & ~_00379_;
	assign _00381_ = _00515_ | io_in[8];
	assign _00382_ = _02096_ & ~_00381_;
	assign _00384_ = _00328_ | _02207_;
	assign _00385_ = _00384_ | _01208_;
	assign _00386_ = io_in[10] & ~_00385_;
	assign _00387_ = io_in[10] & ~_06198_;
	assign _00388_ = _03725_ | io_in[4];
	assign _00389_ = _00388_ | io_in[7];
	assign _00390_ = _06310_ & ~_00389_;
	assign _00391_ = _07301_ | _07422_;
	assign _00392_ = _00391_ | _02096_;
	assign _00393_ = _00392_ | _06310_;
	assign _00395_ = _01985_ & ~_00393_;
	assign _00396_ = _01918_ | _06310_;
	assign _00397_ = io_in[11] & ~_00396_;
	assign _00398_ = _00383_ | io_in[5];
	assign _00399_ = _00398_ | io_in[9];
	assign _00400_ = io_in[10] & ~_00399_;
	assign _00401_ = _01652_ | _02096_;
	assign _00402_ = io_in[10] & ~_00401_;
	assign _00403_ = _00254_ | io_in[6];
	assign _00404_ = _00403_ | _02207_;
	assign _00406_ = io_in[9] & ~_00404_;
	assign _00407_ = _00878_ | io_in[4];
	assign _00408_ = _00407_ | _03759_;
	assign _00409_ = _00408_ | io_in[9];
	assign _00410_ = io_in[11] & ~_00409_;
	assign _00411_ = _00482_ | _01208_;
	assign _00412_ = _00411_ | io_in[9];
	assign _00413_ = io_in[10] & ~_00412_;
	assign _00414_ = _07510_ | io_in[5];
	assign _00415_ = _00414_ | _03759_;
	assign _00417_ = io_in[9] & ~_00415_;
	assign _00418_ = _04580_ | io_in[5];
	assign _00419_ = _00418_ | io_in[6];
	assign _00420_ = _00419_ | io_in[7];
	assign _00421_ = io_in[8] & ~_00420_;
	assign _00422_ = _01485_ | io_in[7];
	assign _00423_ = _00422_ | _01208_;
	assign _00424_ = io_in[10] & ~_00423_;
	assign _00425_ = io_in[5] | ~io_in[2];
	assign _00426_ = _00425_ | _03759_;
	assign _00428_ = _00426_ | io_in[7];
	assign _00429_ = _00428_ | _02096_;
	assign _00430_ = _00429_ | _06310_;
	assign _00431_ = _01985_ & ~_00430_;
	assign _00432_ = _06864_ | _02207_;
	assign _00433_ = io_in[8] & ~_00432_;
	assign _00434_ = _00438_ | io_in[4];
	assign _00435_ = _00434_ | _03759_;
	assign _00436_ = _00435_ | _01208_;
	assign _00437_ = _01985_ & ~_00436_;
	assign _00439_ = _00383_ | io_in[4];
	assign _00440_ = _00439_ | _01208_;
	assign _00441_ = _00440_ | _06310_;
	assign _00442_ = _01985_ & ~_00441_;
	assign _00443_ = _05977_ | _03094_;
	assign _00444_ = _00443_ | io_in[7];
	assign _00445_ = io_in[8] & ~_00444_;
	assign _00446_ = io_in[4] | ~io_in[3];
	assign _00447_ = _00446_ | io_in[5];
	assign _00448_ = _00447_ | _03759_;
	assign _00450_ = _00448_ | _01208_;
	assign _00451_ = io_in[10] & ~_00450_;
	assign _00452_ = _02096_ & ~_00289_;
	assign _00453_ = _07303_ | io_in[7];
	assign _00454_ = io_in[9] & ~_00453_;
	assign _00455_ = _03980_ | io_in[7];
	assign _00456_ = _00455_ | _06310_;
	assign _00457_ = io_in[11] & ~_00456_;
	assign _00458_ = _05977_ | _02207_;
	assign _00459_ = _00458_ | io_in[8];
	assign _00461_ = _02096_ & ~_00459_;
	assign _00462_ = _00398_ | _02207_;
	assign _00463_ = _00462_ | _06310_;
	assign _00464_ = _01985_ & ~_00463_;
	assign _00465_ = _02572_ | _03759_;
	assign _00466_ = _00465_ | io_in[7];
	assign _00467_ = _00466_ | io_in[8];
	assign _00468_ = _00467_ | io_in[9];
	assign _00469_ = _00468_ | io_in[10];
	assign _00470_ = _01985_ & ~_00469_;
	assign _00472_ = _02317_ | _07422_;
	assign _00473_ = _00472_ | _02207_;
	assign _00474_ = _00473_ | _01208_;
	assign _00475_ = io_in[9] & ~_00474_;
	assign _00476_ = _03205_ | _07422_;
	assign _00477_ = _00476_ | _03759_;
	assign _00478_ = _00477_ | io_in[7];
	assign _00479_ = _00478_ | _02096_;
	assign _00480_ = _01985_ & ~_00479_;
	assign _00481_ = _07410_ | io_in[6];
	assign _00483_ = _01208_ & ~_00481_;
	assign _00484_ = _01031_ | _03759_;
	assign _00485_ = _00484_ | _01208_;
	assign _00486_ = _06310_ & ~_00485_;
	assign _00487_ = _01241_ | _02207_;
	assign _00488_ = _00487_ | _02096_;
	assign _00489_ = _00488_ | io_in[10];
	assign _00490_ = _01985_ & ~_00489_;
	assign _00491_ = _00878_ | _03759_;
	assign _00492_ = _00491_ | _02207_;
	assign _00494_ = _00492_ | io_in[9];
	assign _00495_ = _06310_ & ~_00494_;
	assign _00496_ = _05411_ | io_in[5];
	assign _00497_ = _00496_ | _02207_;
	assign _00498_ = _00497_ | _01208_;
	assign _00499_ = io_in[9] & ~_00498_;
	assign _00500_ = _01219_ | io_in[4];
	assign _00501_ = _00500_ | io_in[5];
	assign _00502_ = _00501_ | _03759_;
	assign _00503_ = _00502_ | io_in[8];
	assign _00505_ = io_in[9] & ~_00503_;
	assign _00506_ = _02982_ | io_in[8];
	assign _00507_ = _02096_ & ~_00506_;
	assign _00508_ = _00178_ | io_in[7];
	assign _00509_ = io_in[11] & ~_00508_;
	assign _00510_ = _00325_ | io_in[7];
	assign _00511_ = _01208_ & ~_00510_;
	assign _00512_ = _00333_ | _01208_;
	assign _00513_ = io_in[10] & ~_00512_;
	assign _00514_ = _02029_ | _03759_;
	assign _00516_ = _00514_ | io_in[7];
	assign _00517_ = _02096_ & ~_00516_;
	assign _00518_ = _04136_ | io_in[8];
	assign _00519_ = _00518_ | io_in[10];
	assign _00520_ = _01985_ & ~_00519_;
	assign _00521_ = _06643_ | io_in[3];
	assign _00522_ = _00521_ | io_in[8];
	assign _00523_ = io_in[10] & ~_00522_;
	assign _00524_ = _01762_ | io_in[8];
	assign _00525_ = _00524_ | io_in[9];
	assign _00527_ = _00525_ | io_in[10];
	assign _00528_ = _01985_ & ~_00527_;
	assign _00529_ = _03315_ | _02096_;
	assign _00530_ = io_in[10] & ~_00529_;
	assign _00531_ = _06643_ | io_in[5];
	assign _00532_ = _00531_ | io_in[6];
	assign _00533_ = _00532_ | io_in[7];
	assign _00534_ = io_in[8] & ~_00533_;
	assign _00535_ = io_in[10] & ~_07308_;
	assign _00536_ = _00472_ | io_in[6];
	assign _00538_ = _00536_ | io_in[7];
	assign _00539_ = io_in[10] & ~_00538_;
	assign _00540_ = _06931_ | io_in[6];
	assign _00541_ = io_in[11] & ~_00540_;
	assign _00542_ = io_in[0] | io_in[4];
	assign _00543_ = _00542_ | _03094_;
	assign _00544_ = _00543_ | io_in[6];
	assign _00545_ = _00544_ | _06310_;
	assign _00546_ = io_in[11] & ~_00545_;
	assign _00547_ = _00482_ | _07422_;
	assign _00549_ = _00547_ | io_in[5];
	assign _00550_ = _00549_ | _02207_;
	assign _00551_ = io_in[10] & ~_00550_;
	assign _00552_ = _02305_ | io_in[7];
	assign _00553_ = _00552_ | _01208_;
	assign _00554_ = io_in[11] & ~_00553_;
	assign _00555_ = _04845_ | _01208_;
	assign _00556_ = _00555_ | io_in[9];
	assign _00557_ = _01985_ & ~_00556_;
	assign _00558_ = _02305_ | io_in[8];
	assign _00560_ = io_in[10] & ~_00558_;
	assign _00561_ = _04524_ | _01208_;
	assign _00562_ = io_in[11] & ~_00561_;
	assign _00563_ = _01208_ & ~_00271_;
	assign _00564_ = _02029_ | _02207_;
	assign _00565_ = _06310_ & ~_00564_;
	assign _00566_ = _02229_ | _03759_;
	assign _00567_ = _00566_ | _02207_;
	assign _00568_ = _01985_ & ~_00567_;
	assign _00569_ = _00336_ | _02207_;
	assign _00571_ = _00569_ | _01208_;
	assign _00572_ = _00571_ | _02096_;
	assign _00573_ = _01985_ & ~_00572_;
	assign _00574_ = _01962_ | io_in[6];
	assign _00575_ = _00574_ | io_in[9];
	assign _00576_ = _00575_ | io_in[10];
	assign _00577_ = _01985_ & ~_00576_;
	assign _00578_ = _02206_ | io_in[6];
	assign _00579_ = _00578_ | io_in[7];
	assign _00580_ = _00579_ | io_in[8];
	assign _00582_ = _00580_ | io_in[9];
	assign _00583_ = _00582_ | io_in[10];
	assign _00584_ = io_in[11] & ~_00583_;
	assign _00585_ = _07301_ | io_in[5];
	assign _00586_ = _00585_ | io_in[7];
	assign _00587_ = _00586_ | io_in[10];
	assign _00588_ = io_in[11] & ~_00587_;
	assign _00589_ = _03360_ | io_in[7];
	assign _00590_ = io_in[9] & ~_00589_;
	assign _00591_ = _06176_ | _02207_;
	assign _00593_ = _00591_ | io_in[8];
	assign _00594_ = io_in[11] & ~_00593_;
	assign _00595_ = _01485_ | _03759_;
	assign _00596_ = _00595_ | _02207_;
	assign _00597_ = _01985_ & ~_00596_;
	assign _00598_ = _02505_ | io_in[4];
	assign _00599_ = _00598_ | _03759_;
	assign _00600_ = _00599_ | _02207_;
	assign _00601_ = _00600_ | _02096_;
	assign _00602_ = _01985_ & ~_00601_;
	assign _00604_ = _03881_ | _03759_;
	assign _00605_ = _00604_ | _01208_;
	assign _00606_ = _00605_ | io_in[9];
	assign _00607_ = _01985_ & ~_00606_;
	assign _00608_ = _03980_ | _03759_;
	assign _00609_ = _00608_ | io_in[7];
	assign _00610_ = _00609_ | io_in[8];
	assign _00611_ = _02096_ & ~_00610_;
	assign _00612_ = _00214_ | io_in[7];
	assign _00613_ = _01985_ & ~_00612_;
	assign _00615_ = _07444_ | _02207_;
	assign _00616_ = _00615_ | _01208_;
	assign _00617_ = _00616_ | _02096_;
	assign _00618_ = _01985_ & ~_00617_;
	assign _00619_ = _06642_ | io_in[6];
	assign _00620_ = _00619_ | io_in[7];
	assign _00621_ = _00620_ | io_in[9];
	assign _00622_ = _01985_ & ~_00621_;
	assign _00623_ = _00438_ | io_in[5];
	assign _00624_ = _00623_ | _06310_;
	assign _00626_ = io_in[11] & ~_00624_;
	assign _00627_ = _03980_ | io_in[5];
	assign _00628_ = _00627_ | _03759_;
	assign _00629_ = _00628_ | _02207_;
	assign _00630_ = _00629_ | _01208_;
	assign _00631_ = io_in[9] & ~_00630_;
	assign _00632_ = _07416_ | io_in[7];
	assign _00633_ = _02096_ & ~_00632_;
	assign _00634_ = _07270_ | _02207_;
	assign _00635_ = _00634_ | io_in[8];
	assign _00637_ = io_in[9] & ~_00635_;
	assign _00638_ = _07331_ | _02207_;
	assign _00639_ = _02096_ & ~_00638_;
	assign _00640_ = _01696_ | _02207_;
	assign _00641_ = _01208_ & ~_00640_;
	assign _00642_ = _07330_ | io_in[7];
	assign _00643_ = _00642_ | _01208_;
	assign _00644_ = _06310_ & ~_00643_;
	assign _00645_ = _00473_ | io_in[9];
	assign _00646_ = _06310_ & ~_00645_;
	assign _00648_ = _04580_ | io_in[6];
	assign _00649_ = _00648_ | io_in[7];
	assign _00650_ = _02096_ & ~_00649_;
	assign _00651_ = _06032_ | io_in[9];
	assign _00652_ = _01985_ & ~_00651_;
	assign _00653_ = _00628_ | io_in[9];
	assign _00654_ = io_in[10] & ~_00653_;
	assign _00655_ = _05178_ | io_in[9];
	assign _00656_ = _01985_ & ~_00655_;
	assign _00657_ = _07250_ | io_in[9];
	assign _00659_ = _06310_ & ~_00657_;
	assign _00660_ = _02317_ | io_in[5];
	assign _00661_ = _00660_ | _06310_;
	assign _00662_ = io_in[11] & ~_00661_;
	assign _00663_ = _00548_ | io_in[5];
	assign _00664_ = _00663_ | _03759_;
	assign _00665_ = _00664_ | _02207_;
	assign _00666_ = _00665_ | io_in[8];
	assign _00667_ = _02096_ & ~_00666_;
	assign _00668_ = _01552_ | _01208_;
	assign _00670_ = _06310_ & ~_00668_;
	assign _00671_ = _00663_ | io_in[6];
	assign _00672_ = _00671_ | _02207_;
	assign _00673_ = _00672_ | io_in[8];
	assign _00674_ = io_in[10] & ~_00673_;
	assign _00675_ = _03526_ | _03094_;
	assign _00676_ = _00675_ | io_in[6];
	assign _00677_ = _00676_ | io_in[7];
	assign _00678_ = io_in[10] & ~_00677_;
	assign _00679_ = _07246_ | _03094_;
	assign _00681_ = _00679_ | io_in[8];
	assign _00682_ = io_in[10] & ~_00681_;
	assign _00683_ = _02207_ & ~_00540_;
	assign _00684_ = _00120_ | _07422_;
	assign _00685_ = _00684_ | io_in[10];
	assign _00686_ = io_in[11] & ~_00685_;
	assign _00687_ = _04647_ | _07422_;
	assign _00688_ = _00687_ | _02207_;
	assign _00689_ = _00688_ | _01208_;
	assign _00690_ = _02096_ & ~_00689_;
	assign _00692_ = _00316_ | _02207_;
	assign _00693_ = io_in[10] & ~_00692_;
	assign _00694_ = _01031_ | _01319_;
	assign _00695_ = _00694_ | _02207_;
	assign _00696_ = _06310_ & ~_00695_;
	assign _00697_ = _00694_ | io_in[10];
	assign _00698_ = _01985_ & ~_00697_;
	assign _00699_ = _00271_ | _02207_;
	assign _00700_ = io_in[10] & ~_00699_;
	assign _00701_ = io_in[10] & ~_07438_;
	assign _00703_ = _00178_ | io_in[8];
	assign _00704_ = io_in[9] & ~_00703_;
	assign _00705_ = _04791_ | _03759_;
	assign _00706_ = _00705_ | _02096_;
	assign _00707_ = io_in[11] & ~_00706_;
	assign _00708_ = _06643_ | io_in[4];
	assign _00709_ = _00708_ | io_in[5];
	assign _00710_ = _00709_ | _01208_;
	assign _00711_ = io_in[11] & ~_00710_;
	assign _00712_ = _04302_ | io_in[9];
	assign _00714_ = _01985_ & ~_00712_;
	assign _00715_ = _03316_ | _03759_;
	assign _00716_ = _00715_ | _02207_;
	assign _00717_ = _01985_ & ~_00716_;
	assign _00718_ = _00428_ | io_in[8];
	assign _00719_ = io_in[9] & ~_00718_;
	assign _00720_ = _00439_ | io_in[5];
	assign _00721_ = _00720_ | _02096_;
	assign _00722_ = _01985_ & ~_00721_;
	assign _00723_ = _04934_ | io_in[8];
	assign _00725_ = io_in[10] & ~_00723_;
	assign _00726_ = _07301_ | io_in[8];
	assign _00727_ = _00726_ | io_in[9];
	assign _00728_ = io_in[11] & ~_00727_;
	assign _00729_ = _00570_ | _03759_;
	assign _00730_ = _00729_ | io_in[7];
	assign _00731_ = io_in[11] & ~_00730_;
	assign _00732_ = _01429_ | io_in[5];
	assign _00733_ = _00732_ | _02207_;
	assign _00734_ = io_in[11] & ~_00733_;
	assign _00736_ = io_in[5] | io_in[0];
	assign _00737_ = _00736_ | _03759_;
	assign _00738_ = _00737_ | io_in[7];
	assign _00739_ = _00738_ | io_in[8];
	assign _00740_ = _00739_ | _02096_;
	assign _00741_ = _00740_ | io_in[10];
	assign _00742_ = io_in[11] & ~_00741_;
	assign _00743_ = _07300_ | io_in[5];
	assign _00744_ = _00743_ | _01208_;
	assign _00745_ = _00744_ | io_in[9];
	assign _00747_ = io_in[10] & ~_00745_;
	assign _00748_ = _00347_ | _03759_;
	assign _00749_ = _00748_ | io_in[7];
	assign _00750_ = _00749_ | _01208_;
	assign _00751_ = io_in[10] & ~_00750_;
	assign _00752_ = _02096_ & ~_00595_;
	assign _00753_ = io_in[11] & ~_05467_;
	assign _00754_ = _00336_ | io_in[6];
	assign _00755_ = _00754_ | io_in[7];
	assign _00756_ = _00755_ | _01208_;
	assign _00758_ = io_in[11] & ~_00756_;
	assign _00759_ = _00010_ | io_in[5];
	assign _00760_ = io_in[10] & ~_00759_;
	assign _00761_ = _06975_ | io_in[8];
	assign _00762_ = _00761_ | io_in[9];
	assign _00763_ = io_in[10] & ~_00762_;
	assign _00764_ = _02539_ | io_in[7];
	assign _00765_ = _01208_ & ~_00764_;
	assign _00766_ = _06532_ | _07422_;
	assign _00767_ = _00766_ | _02207_;
	assign _00769_ = _00767_ | io_in[8];
	assign _00770_ = io_in[10] & ~_00769_;
	assign _00771_ = _06620_ | _02207_;
	assign _00772_ = io_in[10] & ~_00771_;
	assign _00773_ = _01596_ | io_in[5];
	assign _00774_ = _00773_ | _02207_;
	assign _00775_ = _00774_ | io_in[9];
	assign _00776_ = io_in[10] & ~_00775_;
	assign _00777_ = _00776_ | _00772_;
	assign _00778_ = _00777_ | _00770_;
	assign _00780_ = _00778_ | _00765_;
	assign _00781_ = _00780_ | _00763_;
	assign _00782_ = _00781_ | _00760_;
	assign _00783_ = _00782_ | _00758_;
	assign _00784_ = _00783_ | _00753_;
	assign _00785_ = _00784_ | _00752_;
	assign _00786_ = _00785_ | _00751_;
	assign _00787_ = _00786_ | _00747_;
	assign _00788_ = _00787_ | _00742_;
	assign _00789_ = _00788_ | _00734_;
	assign _00791_ = _00789_ | _00731_;
	assign _00792_ = _00791_ | _00728_;
	assign _00793_ = _00792_ | _00725_;
	assign _00794_ = _00793_ | _00722_;
	assign _00795_ = _00794_ | _00719_;
	assign _00796_ = _00795_ | _00717_;
	assign _00797_ = _00796_ | _00714_;
	assign _00798_ = _00797_ | _00711_;
	assign _00799_ = _00798_ | _00707_;
	assign _00800_ = _00799_ | _00704_;
	assign _00802_ = _00800_ | _00701_;
	assign _00803_ = _00802_ | _00700_;
	assign _00804_ = _00803_ | _00698_;
	assign _00805_ = _00804_ | _07321_;
	assign _00806_ = _00805_ | _00696_;
	assign _00807_ = _00806_ | _00693_;
	assign _00808_ = _00807_ | _00690_;
	assign _00809_ = _00808_ | _00686_;
	assign _00810_ = _00809_ | _00683_;
	assign _00811_ = _00810_ | _00682_;
	assign _00813_ = _00811_ | _00678_;
	assign _00814_ = _00813_ | _00674_;
	assign _00815_ = _00814_ | _00670_;
	assign _00816_ = _00815_ | _00667_;
	assign _00817_ = _00816_ | _00662_;
	assign _00818_ = _00817_ | _00659_;
	assign _00819_ = _00818_ | _00656_;
	assign _00820_ = _00819_ | _00654_;
	assign _00821_ = _00820_ | _00652_;
	assign _00822_ = _00821_ | _00650_;
	assign _00824_ = _00822_ | _00646_;
	assign _00825_ = _00824_ | _00644_;
	assign _00826_ = _00825_ | _00641_;
	assign _00827_ = _00826_ | _00639_;
	assign _00828_ = _00827_ | _00637_;
	assign _00829_ = _00828_ | _00633_;
	assign _00830_ = _00829_ | _00631_;
	assign _00831_ = _00830_ | _00626_;
	assign _00832_ = _00831_ | _00622_;
	assign _00833_ = _00832_ | _00618_;
	assign _00835_ = _00833_ | _00613_;
	assign _00836_ = _00835_ | _00611_;
	assign _00837_ = _00836_ | _00607_;
	assign _00838_ = _00837_ | _00602_;
	assign _00839_ = _00838_ | _00597_;
	assign _00840_ = _00839_ | _00594_;
	assign _00841_ = _00840_ | _00590_;
	assign _00842_ = _00841_ | _00588_;
	assign _00843_ = _00842_ | _00584_;
	assign _00844_ = _00843_ | _00577_;
	assign _00846_ = _00844_ | _00573_;
	assign _00847_ = _00846_ | _00568_;
	assign _00848_ = _00847_ | _00565_;
	assign _00849_ = _00848_ | _00563_;
	assign _00850_ = _00849_ | _00562_;
	assign _00851_ = _00850_ | _00560_;
	assign _00852_ = _00851_ | _00557_;
	assign _00853_ = _00852_ | _00554_;
	assign _00854_ = _00853_ | _00551_;
	assign _00855_ = _00854_ | _00546_;
	assign _00857_ = _00855_ | _00541_;
	assign _00858_ = _00857_ | _00539_;
	assign _00859_ = _00858_ | _00535_;
	assign _00860_ = _00859_ | _00534_;
	assign _00861_ = _00860_ | _00530_;
	assign _00862_ = _00861_ | _00528_;
	assign _00863_ = _00862_ | _00523_;
	assign _00864_ = _00863_ | _00520_;
	assign _00865_ = _00864_ | _00517_;
	assign _00866_ = _00865_ | _00513_;
	assign _00868_ = _00866_ | _00511_;
	assign _00869_ = _00868_ | _00509_;
	assign _00870_ = _00869_ | _00507_;
	assign _00871_ = _00870_ | _00505_;
	assign _00872_ = _00871_ | _00499_;
	assign _00873_ = _00872_ | _00495_;
	assign _00874_ = _00873_ | _00490_;
	assign _00875_ = _00874_ | _00486_;
	assign _00876_ = _00875_ | _00483_;
	assign _00877_ = _00876_ | _00480_;
	assign _00879_ = _00877_ | _00475_;
	assign _00880_ = _00879_ | _00470_;
	assign _00881_ = _00880_ | _00464_;
	assign _00882_ = _00881_ | _00461_;
	assign _00883_ = _00882_ | _00457_;
	assign _00884_ = _00883_ | _00454_;
	assign _00885_ = _00884_ | _00452_;
	assign _00886_ = _00885_ | _00451_;
	assign _00887_ = _00886_ | _00445_;
	assign _00888_ = _00887_ | _00442_;
	assign _00890_ = _00888_ | _00437_;
	assign _00891_ = _00890_ | _00433_;
	assign _00892_ = _00891_ | _00431_;
	assign _00893_ = _00892_ | _00424_;
	assign _00894_ = _00893_ | _00421_;
	assign _00895_ = _00894_ | _00417_;
	assign _00896_ = _00895_ | _00413_;
	assign _00897_ = _00896_ | _00410_;
	assign _00898_ = _00897_ | _00406_;
	assign _00899_ = _00898_ | _00402_;
	assign _00901_ = _00899_ | _00400_;
	assign _00902_ = _00901_ | _00397_;
	assign _00903_ = _00902_ | _00395_;
	assign _00904_ = _00903_ | _00390_;
	assign _00905_ = _00904_ | _00387_;
	assign _00906_ = _00905_ | _00386_;
	assign _00907_ = _00906_ | _00382_;
	assign _00908_ = _00907_ | _00380_;
	assign _00909_ = _00908_ | _00376_;
	assign _00910_ = _00909_ | _00371_;
	assign _00912_ = _00910_ | _00367_;
	assign _00913_ = _00912_ | _00365_;
	assign _00914_ = _00913_ | _00363_;
	assign _00915_ = _00914_ | _00359_;
	assign _00916_ = _00915_ | _00357_;
	assign _00917_ = _00916_ | _00354_;
	assign _00918_ = _00917_ | _00352_;
	assign _00919_ = _00918_ | _00346_;
	assign _00920_ = _00919_ | _00344_;
	assign _00921_ = _00920_ | _00342_;
	assign _00923_ = _00921_ | _00340_;
	assign _00924_ = _00923_ | _00335_;
	assign _00925_ = _00924_ | _00332_;
	assign _00926_ = _00925_ | _00327_;
	assign _00927_ = _00926_ | _00324_;
	assign _00928_ = _00927_ | _00320_;
	assign _00929_ = _00928_ | _00315_;
	assign _00930_ = _00929_ | _00312_;
	assign _00931_ = _00930_ | _00305_;
	assign _00932_ = _00931_ | _00303_;
	assign _00934_ = _00932_ | _00296_;
	assign _00935_ = _00934_ | _00291_;
	assign _00936_ = _00935_ | _00288_;
	assign _00937_ = _00936_ | _00285_;
	assign _00938_ = _00937_ | _00280_;
	assign _00939_ = _00938_ | _00278_;
	assign _00940_ = _00939_ | _00275_;
	assign _00941_ = _00940_ | _00272_;
	assign _00942_ = _00941_ | _00270_;
	assign _00943_ = _00942_ | _00266_;
	assign _00945_ = _00943_ | _00263_;
	assign _00946_ = _00945_ | _00257_;
	assign _00947_ = _00946_ | _00253_;
	assign _00948_ = _00947_ | _00249_;
	assign _00949_ = _00948_ | _00248_;
	assign _00950_ = _00949_ | _00244_;
	assign _00951_ = _00950_ | _00238_;
	assign _00952_ = _00951_ | _00234_;
	assign _00953_ = _00952_ | _00231_;
	assign _00954_ = _00953_ | _00226_;
	assign _00956_ = _00954_ | _00220_;
	assign _00957_ = _00956_ | _00216_;
	assign _00958_ = _00957_ | _00213_;
	assign _00959_ = _00958_ | _00208_;
	assign _00960_ = _00959_ | _00201_;
	assign _00961_ = _00960_ | _00197_;
	assign _00962_ = _00961_ | _00195_;
	assign _00963_ = _00962_ | _00191_;
	assign _00964_ = _00963_ | _00186_;
	assign _00965_ = _00964_ | _00181_;
	assign _00967_ = _00965_ | _00180_;
	assign _00968_ = _00967_ | _00177_;
	assign _00969_ = _00968_ | _00172_;
	assign _00970_ = _00969_ | _00168_;
	assign \mchip.val [5] = _00970_ | _00165_;
	assign _00971_ = _06853_ | io_in[4];
	assign _00972_ = _00971_ | io_in[5];
	assign _00973_ = _00972_ | _03759_;
	assign _00974_ = _00973_ | _02207_;
	assign _00975_ = _00974_ | _01208_;
	assign _00977_ = _00975_ | _02096_;
	assign _00978_ = _06310_ & ~_00977_;
	assign _00979_ = _01042_ | io_in[5];
	assign _00980_ = _00979_ | _03759_;
	assign _00981_ = _00980_ | io_in[7];
	assign _00982_ = _00981_ | io_in[8];
	assign _00983_ = _00982_ | _02096_;
	assign _00984_ = io_in[10] & ~_00983_;
	assign _00985_ = _07499_ | _01319_;
	assign _00986_ = _00985_ | io_in[4];
	assign _00988_ = _00986_ | io_in[6];
	assign _00989_ = _00988_ | _02207_;
	assign _00990_ = _00989_ | _01208_;
	assign _00991_ = _00990_ | _02096_;
	assign _00992_ = _06310_ & ~_00991_;
	assign _00993_ = _00812_ | _03759_;
	assign _00994_ = _00993_ | _02207_;
	assign _00995_ = _00994_ | _06310_;
	assign _00996_ = io_in[11] & ~_00995_;
	assign _00997_ = _07098_ | _01208_;
	assign _00999_ = _00997_ | io_in[10];
	assign _01000_ = io_in[11] & ~_00999_;
	assign _01001_ = _07257_ | _07422_;
	assign _01002_ = _01001_ | io_in[6];
	assign _01003_ = _01002_ | _02207_;
	assign _01004_ = _01003_ | io_in[8];
	assign _01005_ = io_in[11] & ~_01004_;
	assign _01006_ = _00493_ | _01319_;
	assign _01007_ = _01006_ | io_in[4];
	assign _01008_ = _01007_ | io_in[8];
	assign _01010_ = _01008_ | io_in[9];
	assign _01011_ = _01010_ | io_in[10];
	assign _01012_ = _01985_ & ~_01011_;
	assign _01013_ = _07257_ | io_in[4];
	assign _01014_ = _01013_ | _02207_;
	assign _01015_ = _01014_ | _06310_;
	assign _01016_ = io_in[11] & ~_01015_;
	assign _01017_ = _00521_ | _07422_;
	assign _01018_ = _01017_ | io_in[6];
	assign _01019_ = _01018_ | _02207_;
	assign _01021_ = _01019_ | _02096_;
	assign _01022_ = _01021_ | _06310_;
	assign _01023_ = _01985_ & ~_01022_;
	assign _01024_ = _01006_ | _07422_;
	assign _01025_ = _01024_ | _03759_;
	assign _01026_ = _01025_ | _02207_;
	assign _01027_ = _01026_ | _01208_;
	assign _01028_ = io_in[9] & ~_01027_;
	assign _01029_ = _01001_ | _03759_;
	assign _01030_ = _01029_ | _02207_;
	assign _01032_ = _01030_ | io_in[8];
	assign _01033_ = _01032_ | _02096_;
	assign _01034_ = io_in[10] & ~_01033_;
	assign _01035_ = _01029_ | io_in[9];
	assign _01036_ = _01035_ | io_in[10];
	assign _01037_ = _01985_ & ~_01036_;
	assign _01038_ = _00274_ | io_in[5];
	assign _01039_ = _01038_ | _03759_;
	assign _01040_ = _01039_ | _02207_;
	assign _01041_ = _01040_ | _01208_;
	assign _01043_ = _01041_ | _02096_;
	assign _01044_ = _01043_ | _06310_;
	assign _01045_ = _01985_ & ~_01044_;
	assign _01046_ = _03260_ | io_in[6];
	assign _01047_ = _01046_ | io_in[7];
	assign _01048_ = _01047_ | _02096_;
	assign _01049_ = _01048_ | _06310_;
	assign _01050_ = _01985_ & ~_01049_;
	assign _01051_ = _00246_ | _03759_;
	assign _01052_ = _01051_ | io_in[7];
	assign _01054_ = _01052_ | io_in[8];
	assign _01055_ = _01054_ | io_in[9];
	assign _01056_ = io_in[11] & ~_01055_;
	assign _01057_ = _02018_ | io_in[4];
	assign _01058_ = _01057_ | io_in[5];
	assign _01059_ = _01058_ | _03759_;
	assign _01060_ = _01059_ | io_in[7];
	assign _01061_ = _01060_ | io_in[8];
	assign _01062_ = _01061_ | io_in[9];
	assign _01063_ = _01062_ | _06310_;
	assign _01065_ = _01985_ & ~_01063_;
	assign _01066_ = _00131_ | io_in[6];
	assign _01067_ = _01066_ | io_in[7];
	assign _01068_ = _01067_ | io_in[8];
	assign _01069_ = _01068_ | io_in[9];
	assign _01070_ = _01069_ | io_in[10];
	assign _01071_ = io_in[11] & ~_01070_;
	assign _01072_ = _07335_ | io_in[4];
	assign _01073_ = _01072_ | _03759_;
	assign _01074_ = _01073_ | _02207_;
	assign _01076_ = _01074_ | _01208_;
	assign _01077_ = _01076_ | io_in[10];
	assign _01078_ = io_in[11] & ~_01077_;
	assign _01079_ = _00250_ | _03759_;
	assign _01080_ = _01079_ | _02207_;
	assign _01081_ = _01080_ | _01208_;
	assign _01082_ = _01081_ | _02096_;
	assign _01083_ = io_in[10] & ~_01082_;
	assign _01084_ = _00724_ | _02207_;
	assign _01085_ = _01084_ | _02096_;
	assign _01087_ = _01085_ | io_in[10];
	assign _01088_ = io_in[11] & ~_01087_;
	assign _01089_ = _03249_ | _03094_;
	assign _01090_ = _01089_ | _03759_;
	assign _01091_ = _02096_ & ~_01090_;
	assign _01092_ = _00759_ | io_in[6];
	assign _01093_ = _01092_ | _02207_;
	assign _01094_ = _01093_ | _02096_;
	assign _01095_ = io_in[11] & ~_01094_;
	assign _01096_ = _03603_ | _03759_;
	assign _01098_ = _01096_ | io_in[7];
	assign _01099_ = _01098_ | _06310_;
	assign _01100_ = io_in[11] & ~_01099_;
	assign _01101_ = _01013_ | io_in[6];
	assign _01102_ = _01101_ | io_in[7];
	assign _01103_ = _01102_ | io_in[10];
	assign _01104_ = _01985_ & ~_01103_;
	assign _01105_ = _00709_ | _03759_;
	assign _01106_ = _01105_ | _02207_;
	assign _01107_ = _01106_ | io_in[8];
	assign _01109_ = _01107_ | io_in[9];
	assign _01110_ = io_in[10] & ~_01109_;
	assign _01111_ = _00246_ | io_in[6];
	assign _01112_ = _01111_ | io_in[7];
	assign _01113_ = _01112_ | _02096_;
	assign _01114_ = _06310_ & ~_01113_;
	assign _01115_ = _06931_ | _07422_;
	assign _01116_ = _01115_ | io_in[5];
	assign _01117_ = _01116_ | _03759_;
	assign _01118_ = _01117_ | _01208_;
	assign _01120_ = io_in[11] & ~_01118_;
	assign _01121_ = _07336_ | io_in[7];
	assign _01122_ = _01121_ | io_in[8];
	assign _01123_ = _01122_ | io_in[9];
	assign _01124_ = io_in[11] & ~_01123_;
	assign _01125_ = _07246_ | io_in[4];
	assign _01126_ = _01125_ | io_in[6];
	assign _01127_ = _01126_ | _02207_;
	assign _01128_ = _01127_ | io_in[8];
	assign _01129_ = _01128_ | _02096_;
	assign _01131_ = _01129_ | io_in[10];
	assign _01132_ = _01985_ & ~_01131_;
	assign _01133_ = _01072_ | io_in[6];
	assign _01134_ = _01133_ | io_in[7];
	assign _01135_ = _01134_ | _01208_;
	assign _01136_ = _01135_ | io_in[10];
	assign _01137_ = io_in[11] & ~_01136_;
	assign _01138_ = _07301_ | _03094_;
	assign _01139_ = _01138_ | _03759_;
	assign _01140_ = _01139_ | _02096_;
	assign _01142_ = _06310_ & ~_01140_;
	assign _01143_ = _06520_ | _03759_;
	assign _01144_ = _01143_ | _02207_;
	assign _01145_ = _01144_ | io_in[8];
	assign _01146_ = _01145_ | _02096_;
	assign _01147_ = io_in[10] & ~_01146_;
	assign _01148_ = _01541_ | _07422_;
	assign _01149_ = _01148_ | io_in[7];
	assign _01150_ = _01149_ | _01208_;
	assign _01151_ = _01150_ | _02096_;
	assign _01153_ = _06310_ & ~_01151_;
	assign _01154_ = _04325_ | _01208_;
	assign _01155_ = _01154_ | io_in[9];
	assign _01156_ = io_in[10] & ~_01155_;
	assign _01157_ = _01296_ | _03094_;
	assign _01158_ = _01157_ | io_in[6];
	assign _01159_ = _01158_ | _02207_;
	assign _01160_ = _01159_ | io_in[9];
	assign _01161_ = io_in[10] & ~_01160_;
	assign _01162_ = _00684_ | io_in[6];
	assign _01164_ = _01162_ | io_in[7];
	assign _01165_ = _01164_ | _01208_;
	assign _01166_ = _01165_ | io_in[9];
	assign _01167_ = io_in[11] & ~_01166_;
	assign _01168_ = _00759_ | _03759_;
	assign _01169_ = _01168_ | _02207_;
	assign _01170_ = _01169_ | io_in[8];
	assign _01171_ = io_in[10] & ~_01170_;
	assign _01172_ = _03981_ | io_in[4];
	assign _01173_ = _01172_ | io_in[5];
	assign _01175_ = _01173_ | _03759_;
	assign _01176_ = _01175_ | _01208_;
	assign _01177_ = _01176_ | _02096_;
	assign _01178_ = _01177_ | io_in[10];
	assign _01179_ = _01985_ & ~_01178_;
	assign _01180_ = _01115_ | _02207_;
	assign _01181_ = _01180_ | _01208_;
	assign _01182_ = _01181_ | io_in[10];
	assign _01183_ = io_in[11] & ~_01182_;
	assign _01184_ = _01115_ | io_in[6];
	assign _01186_ = _01184_ | io_in[7];
	assign _01187_ = _01186_ | _01208_;
	assign _01188_ = _01187_ | _02096_;
	assign _01189_ = _06310_ & ~_01188_;
	assign _01190_ = _06864_ | io_in[4];
	assign _01191_ = _01190_ | _03759_;
	assign _01192_ = _01191_ | io_in[7];
	assign _01193_ = _01192_ | io_in[8];
	assign _01194_ = io_in[11] & ~_01193_;
	assign _01195_ = _04978_ | io_in[6];
	assign _01197_ = _01195_ | io_in[8];
	assign _01198_ = _01197_ | io_in[9];
	assign _01199_ = io_in[11] & ~_01198_;
	assign _01200_ = _06853_ | io_in[3];
	assign _01201_ = _01200_ | _07422_;
	assign _01202_ = _01201_ | _03759_;
	assign _01203_ = _01202_ | io_in[7];
	assign _01204_ = _02096_ & ~_01203_;
	assign _01205_ = _01204_ & ~_06310_;
	assign _01206_ = _04458_ | _03759_;
	assign _01209_ = _01206_ | io_in[8];
	assign _01210_ = _01209_ | _02096_;
	assign _01211_ = _01210_ | io_in[10];
	assign _01212_ = _01985_ & ~_01211_;
	assign _01213_ = _01042_ | io_in[4];
	assign _01214_ = _01213_ | io_in[5];
	assign _01215_ = _01214_ | _03759_;
	assign _01216_ = _01215_ | _02096_;
	assign _01217_ = _01216_ | io_in[10];
	assign _01218_ = _01985_ & ~_01217_;
	assign _01220_ = _04647_ | _03094_;
	assign _01221_ = _01220_ | io_in[6];
	assign _01222_ = _01221_ | io_in[8];
	assign _01223_ = _01222_ | _02096_;
	assign _01224_ = io_in[10] & ~_01223_;
	assign _01225_ = _01200_ | io_in[4];
	assign _01226_ = _01225_ | io_in[6];
	assign _01227_ = _01226_ | _02207_;
	assign _01228_ = _01227_ | _02096_;
	assign _01229_ = _01228_ | io_in[10];
	assign _01231_ = io_in[11] & ~_01229_;
	assign _01232_ = _00353_ | _06310_;
	assign _01233_ = io_in[11] & ~_01232_;
	assign _01234_ = _00245_ | io_in[4];
	assign _01235_ = _01234_ | io_in[5];
	assign _01236_ = _01235_ | _03759_;
	assign _01237_ = _01236_ | io_in[7];
	assign _01238_ = _01237_ | io_in[9];
	assign _01239_ = _01238_ | io_in[10];
	assign _01240_ = _01985_ & ~_01239_;
	assign _01242_ = _00274_ | _01208_;
	assign _01243_ = _01242_ | io_in[9];
	assign _01244_ = _01243_ | io_in[10];
	assign _01245_ = _01985_ & ~_01244_;
	assign _01246_ = _07142_ | io_in[6];
	assign _01247_ = _01246_ | io_in[7];
	assign _01248_ = _01247_ | _01208_;
	assign _01249_ = _01248_ | io_in[9];
	assign _01250_ = io_in[10] & ~_01249_;
	assign _01251_ = _06864_ | _07422_;
	assign _01253_ = _01251_ | io_in[7];
	assign _01254_ = _01253_ | io_in[8];
	assign _01255_ = _01254_ | _02096_;
	assign _01256_ = io_in[10] & ~_01255_;
	assign _01257_ = _06000_ | _01208_;
	assign _01258_ = _01257_ | io_in[9];
	assign _01259_ = io_in[10] & ~_01258_;
	assign _01260_ = _07419_ | io_in[5];
	assign _01261_ = _01260_ | _02207_;
	assign _01262_ = _01261_ | io_in[8];
	assign _01264_ = _01262_ | _02096_;
	assign _01265_ = io_in[11] & ~_01264_;
	assign _01266_ = _07255_ | _03759_;
	assign _01267_ = _01266_ | io_in[8];
	assign _01268_ = _01267_ | io_in[9];
	assign _01269_ = io_in[10] & ~_01268_;
	assign _01270_ = _07413_ | _02096_;
	assign _01271_ = io_in[11] & ~_01270_;
	assign _01272_ = _00979_ | io_in[6];
	assign _01273_ = _01272_ | _02207_;
	assign _01275_ = _01273_ | _01208_;
	assign _01276_ = _06310_ & ~_01275_;
	assign _01277_ = _07255_ | io_in[5];
	assign _01278_ = _01277_ | io_in[6];
	assign _01279_ = _01278_ | _01208_;
	assign _01280_ = _01279_ | _06310_;
	assign _01281_ = _01985_ & ~_01280_;
	assign _01282_ = _00245_ | _03094_;
	assign _01283_ = _01282_ | _03759_;
	assign _01284_ = _01283_ | _01208_;
	assign _01286_ = _01284_ | _06310_;
	assign _01287_ = _01985_ & ~_01286_;
	assign _01288_ = _01214_ | _01208_;
	assign _01289_ = _01288_ | _02096_;
	assign _01290_ = _06310_ & ~_01289_;
	assign _01291_ = _01092_ | io_in[7];
	assign _01292_ = _01291_ | io_in[8];
	assign _01293_ = _02096_ & ~_01292_;
	assign _01294_ = _03116_ | io_in[6];
	assign _01295_ = _01294_ | io_in[7];
	assign _01297_ = _01295_ | io_in[8];
	assign _01298_ = io_in[10] & ~_01297_;
	assign _01299_ = _03647_ | _02207_;
	assign _01300_ = _01299_ | _06310_;
	assign _01301_ = io_in[11] & ~_01300_;
	assign _01302_ = _00660_ | _03759_;
	assign _01303_ = _01302_ | io_in[7];
	assign _01304_ = _01303_ | _06310_;
	assign _01305_ = io_in[11] & ~_01304_;
	assign _01306_ = _01007_ | io_in[5];
	assign _01308_ = _01306_ | io_in[6];
	assign _01309_ = _01308_ | _02207_;
	assign _01310_ = _01309_ | _02096_;
	assign _01311_ = io_in[11] & ~_01310_;
	assign _01312_ = _01168_ | io_in[7];
	assign _01313_ = io_in[11] & ~_01312_;
	assign _01314_ = _07433_ | _03094_;
	assign _01315_ = _01314_ | _03759_;
	assign _01316_ = _01315_ | _02207_;
	assign _01317_ = _01316_ | _02096_;
	assign _01320_ = io_in[11] & ~_01317_;
	assign _01321_ = _02428_ | _07422_;
	assign _01322_ = _01321_ | _03759_;
	assign _01323_ = _01322_ | _02207_;
	assign _01324_ = _01323_ | _02096_;
	assign _01325_ = _01324_ | io_in[10];
	assign _01326_ = _01985_ & ~_01325_;
	assign _01327_ = _01051_ | _02207_;
	assign _01328_ = _01327_ | _01208_;
	assign _01329_ = io_in[10] & ~_01328_;
	assign _01331_ = _05900_ | _02207_;
	assign _01332_ = _01331_ | _06310_;
	assign _01333_ = io_in[11] & ~_01332_;
	assign _01334_ = _07410_ | io_in[4];
	assign _01335_ = _01334_ | io_in[6];
	assign _01336_ = _01335_ | io_in[7];
	assign _01337_ = _01336_ | _01208_;
	assign _01338_ = _01337_ | _02096_;
	assign _01339_ = _06310_ & ~_01338_;
	assign _01340_ = _00245_ | io_in[5];
	assign _01342_ = _01340_ | io_in[6];
	assign _01343_ = _01342_ | io_in[7];
	assign _01344_ = _01343_ | _01208_;
	assign _01345_ = _01344_ | io_in[9];
	assign _01346_ = _01345_ | _06310_;
	assign _01347_ = _01985_ & ~_01346_;
	assign _01348_ = _01007_ | io_in[6];
	assign _01349_ = _01348_ | io_in[7];
	assign _01350_ = _01349_ | _01208_;
	assign _01351_ = _01350_ | _06310_;
	assign _01353_ = _01985_ & ~_01351_;
	assign _01354_ = _01172_ | _03759_;
	assign _01355_ = _01354_ | _02207_;
	assign _01356_ = _01355_ | _01208_;
	assign _01357_ = _01356_ | io_in[9];
	assign _01358_ = _01357_ | _06310_;
	assign _01359_ = _01985_ & ~_01358_;
	assign _01360_ = _00985_ | _07422_;
	assign _01361_ = _01360_ | io_in[6];
	assign _01362_ = _01361_ | io_in[7];
	assign _01364_ = _01362_ | _02096_;
	assign _01365_ = io_in[11] & ~_01364_;
	assign _01366_ = _01013_ | io_in[5];
	assign _01367_ = _01366_ | io_in[6];
	assign _01368_ = _01367_ | io_in[8];
	assign _01369_ = _01368_ | io_in[9];
	assign _01370_ = io_in[11] & ~_01369_;
	assign _01371_ = _06032_ | _01208_;
	assign _01372_ = _01371_ | _02096_;
	assign _01373_ = _01372_ | _06310_;
	assign _01375_ = _01985_ & ~_01373_;
	assign _01376_ = _01072_ | _02207_;
	assign _01377_ = _01376_ | io_in[8];
	assign _01378_ = _01377_ | _02096_;
	assign _01379_ = io_in[11] & ~_01378_;
	assign _01380_ = _04302_ | io_in[6];
	assign _01381_ = _01380_ | _01208_;
	assign _01382_ = _01381_ | _02096_;
	assign _01383_ = _01382_ | _06310_;
	assign _01384_ = _01985_ & ~_01383_;
	assign _01386_ = _06754_ | _07422_;
	assign _01387_ = _01386_ | _02207_;
	assign _01388_ = _01387_ | io_in[9];
	assign _01389_ = _01388_ | io_in[10];
	assign _01390_ = _01985_ & ~_01389_;
	assign _01391_ = _00493_ | _03094_;
	assign _01392_ = _01391_ | io_in[7];
	assign _01393_ = _01392_ | io_in[9];
	assign _01394_ = io_in[10] & ~_01393_;
	assign _01395_ = _04978_ | io_in[7];
	assign _01397_ = _01395_ | io_in[8];
	assign _01398_ = _01397_ | _02096_;
	assign _01399_ = io_in[10] & ~_01398_;
	assign _01400_ = _01541_ | _03759_;
	assign _01401_ = _01400_ | _02207_;
	assign _01402_ = _01401_ | _06310_;
	assign _01403_ = io_in[11] & ~_01402_;
	assign _01404_ = _02672_ | _01319_;
	assign _01405_ = _01404_ | _07422_;
	assign _01406_ = _01405_ | _03759_;
	assign _01408_ = _01406_ | _02207_;
	assign _01409_ = _01408_ | io_in[8];
	assign _01410_ = io_in[11] & ~_01409_;
	assign _01411_ = _02672_ | _03094_;
	assign _01412_ = _01411_ | io_in[6];
	assign _01413_ = _01412_ | io_in[7];
	assign _01414_ = _01413_ | io_in[8];
	assign _01415_ = io_in[11] & ~_01414_;
	assign _01416_ = _01201_ | io_in[6];
	assign _01417_ = _01416_ | _02207_;
	assign _01419_ = _01417_ | _01208_;
	assign _01420_ = io_in[9] & ~_01419_;
	assign _01421_ = _02860_ | io_in[5];
	assign _01422_ = _01421_ | io_in[6];
	assign _01423_ = _01422_ | _02207_;
	assign _01424_ = _01423_ | io_in[8];
	assign _01425_ = _01424_ | io_in[9];
	assign _01426_ = io_in[11] & ~_01425_;
	assign _01427_ = _06243_ | io_in[6];
	assign _01428_ = _01427_ | io_in[7];
	assign _01431_ = _01428_ | io_in[8];
	assign _01432_ = _01431_ | _02096_;
	assign _01433_ = io_in[11] & ~_01432_;
	assign _01434_ = _01405_ | io_in[6];
	assign _01435_ = _01434_ | _02207_;
	assign _01436_ = _01435_ | _01208_;
	assign _01437_ = io_in[11] & ~_01436_;
	assign _01438_ = _04458_ | io_in[4];
	assign _01439_ = _01438_ | _03759_;
	assign _01440_ = _01439_ | io_in[7];
	assign _01442_ = _01440_ | io_in[8];
	assign _01443_ = _01442_ | io_in[9];
	assign _01444_ = io_in[11] & ~_01443_;
	assign _01445_ = _03127_ | io_in[7];
	assign _01446_ = _01445_ | _06310_;
	assign _01447_ = io_in[11] & ~_01446_;
	assign _01448_ = _01039_ | io_in[8];
	assign _01449_ = _01448_ | io_in[9];
	assign _01450_ = io_in[10] & ~_01449_;
	assign _01451_ = _01235_ | io_in[6];
	assign _01453_ = _01451_ | _02207_;
	assign _01454_ = _01453_ | _02096_;
	assign _01455_ = _01985_ & ~_01454_;
	assign _01456_ = _00548_ | _03094_;
	assign _01457_ = _01456_ | _03759_;
	assign _01458_ = _01457_ | _01208_;
	assign _01459_ = _02096_ & ~_01458_;
	assign _01460_ = _00391_ | io_in[6];
	assign _01461_ = _01460_ | _02207_;
	assign _01462_ = _01461_ | io_in[8];
	assign _01464_ = _01462_ | io_in[9];
	assign _01465_ = io_in[11] & ~_01464_;
	assign _01466_ = _01192_ | _01208_;
	assign _01467_ = _01466_ | io_in[9];
	assign _01468_ = io_in[10] & ~_01467_;
	assign _01469_ = _00407_ | io_in[5];
	assign _01470_ = _01469_ | io_in[6];
	assign _01471_ = _01470_ | _02207_;
	assign _01472_ = _01471_ | _06310_;
	assign _01473_ = io_in[11] & ~_01472_;
	assign _01475_ = _02018_ | _03094_;
	assign _01476_ = _01475_ | io_in[6];
	assign _01477_ = _01476_ | io_in[8];
	assign _01478_ = _01477_ | io_in[9];
	assign _01479_ = io_in[11] & ~_01478_;
	assign _01480_ = _00481_ | io_in[7];
	assign _01481_ = _01480_ | io_in[8];
	assign _01482_ = _02096_ & ~_01481_;
	assign _01483_ = _00694_ | io_in[4];
	assign _01484_ = _01483_ | _03759_;
	assign _01486_ = _01484_ | _02207_;
	assign _01487_ = _01486_ | io_in[8];
	assign _01488_ = _01487_ | _02096_;
	assign _01489_ = io_in[10] & ~_01488_;
	assign _01490_ = _05977_ | _03759_;
	assign _01491_ = _01490_ | _01208_;
	assign _01492_ = _01491_ | io_in[9];
	assign _01493_ = io_in[10] & ~_01492_;
	assign _01494_ = _01112_ | _01208_;
	assign _01495_ = _01494_ | _06310_;
	assign _01497_ = _01985_ & ~_01495_;
	assign _01498_ = _01026_ | io_in[9];
	assign _01499_ = _01985_ & ~_01498_;
	assign _01500_ = _07351_ | io_in[6];
	assign _01501_ = _01500_ | io_in[7];
	assign _01502_ = _01501_ | io_in[8];
	assign _01503_ = _01502_ | _02096_;
	assign _01504_ = io_in[10] & ~_01503_;
	assign _01505_ = _02272_ | _03759_;
	assign _01506_ = _01505_ | _02207_;
	assign _01508_ = _01506_ | io_in[8];
	assign _01509_ = io_in[11] & ~_01508_;
	assign _01510_ = _01072_ | io_in[5];
	assign _01511_ = _01510_ | _02207_;
	assign _01512_ = _01511_ | io_in[9];
	assign _01513_ = _01512_ | io_in[10];
	assign _01514_ = _01985_ & ~_01513_;
	assign _01515_ = _02916_ | io_in[6];
	assign _01516_ = _01515_ | _02207_;
	assign _01517_ = _01516_ | _01208_;
	assign _01519_ = _01517_ | io_in[9];
	assign _01520_ = io_in[10] & ~_01519_;
	assign _01521_ = _07410_ | io_in[5];
	assign _01522_ = _01521_ | io_in[6];
	assign _01523_ = _01522_ | io_in[8];
	assign _01524_ = _01523_ | io_in[9];
	assign _01525_ = _06310_ & ~_01524_;
	assign _01526_ = _02040_ | io_in[7];
	assign _01527_ = _01526_ | _01208_;
	assign _01528_ = _01527_ | io_in[10];
	assign _01530_ = io_in[11] & ~_01528_;
	assign _01531_ = _01361_ | _01208_;
	assign _01532_ = _01531_ | io_in[9];
	assign _01533_ = io_in[10] & ~_01532_;
	assign _01534_ = _01017_ | _02207_;
	assign _01535_ = _01534_ | io_in[10];
	assign _01536_ = io_in[11] & ~_01535_;
	assign _01537_ = _04458_ | _07422_;
	assign _01538_ = _01537_ | io_in[6];
	assign _01539_ = _01538_ | io_in[7];
	assign _01542_ = _01539_ | io_in[9];
	assign _01543_ = io_in[11] & ~_01542_;
	assign _01544_ = _06976_ | io_in[7];
	assign _01545_ = _01544_ | io_in[9];
	assign _01546_ = io_in[11] & ~_01545_;
	assign _01547_ = _01321_ | io_in[6];
	assign _01548_ = _01547_ | _02207_;
	assign _01549_ = _01548_ | io_in[8];
	assign _01550_ = _01549_ | _02096_;
	assign _01551_ = io_in[11] & ~_01550_;
	assign _01553_ = _00598_ | io_in[6];
	assign _01554_ = _01553_ | io_in[7];
	assign _01555_ = _01554_ | io_in[10];
	assign _01556_ = _01985_ & ~_01555_;
	assign _01557_ = _01173_ | io_in[6];
	assign _01558_ = _01557_ | _02207_;
	assign _01559_ = _01558_ | _01208_;
	assign _01560_ = _01559_ | io_in[9];
	assign _01561_ = _01560_ | io_in[10];
	assign _01562_ = io_in[11] & ~_01561_;
	assign _01564_ = _03027_ | io_in[7];
	assign _01565_ = _01564_ | _01208_;
	assign _01566_ = _01565_ | io_in[9];
	assign _01567_ = io_in[10] & ~_01566_;
	assign _01568_ = _06931_ | _03759_;
	assign _01569_ = _01568_ | _02207_;
	assign _01570_ = _01569_ | io_in[8];
	assign _01571_ = _01570_ | io_in[9];
	assign _01572_ = io_in[10] & ~_01571_;
	assign _01573_ = _00135_ | io_in[7];
	assign _01575_ = _01573_ | io_in[8];
	assign _01576_ = _01575_ | _02096_;
	assign _01577_ = io_in[10] & ~_01576_;
	assign _01578_ = _01273_ | io_in[8];
	assign _01579_ = io_in[10] & ~_01578_;
	assign _01580_ = _01251_ | io_in[6];
	assign _01581_ = _01580_ | _02207_;
	assign _01582_ = _06310_ & ~_01581_;
	assign _01583_ = _06865_ | io_in[5];
	assign _01584_ = _01583_ | _02207_;
	assign _01586_ = _01584_ | io_in[8];
	assign _01587_ = _01586_ | io_in[9];
	assign _01588_ = io_in[10] & ~_01587_;
	assign _01589_ = _01485_ | _03094_;
	assign _01590_ = _01589_ | io_in[6];
	assign _01591_ = _01590_ | io_in[7];
	assign _01592_ = _01591_ | _06310_;
	assign _01593_ = io_in[11] & ~_01592_;
	assign _01594_ = _07402_ | io_in[5];
	assign _01595_ = _01594_ | _03759_;
	assign _01597_ = _01595_ | _02207_;
	assign _01598_ = _01597_ | io_in[8];
	assign _01599_ = _01598_ | _02096_;
	assign _01600_ = io_in[10] & ~_01599_;
	assign _01601_ = _00383_ | _03094_;
	assign _01602_ = _01601_ | _03759_;
	assign _01603_ = _01602_ | _02207_;
	assign _01604_ = _01603_ | io_in[9];
	assign _01605_ = io_in[10] & ~_01604_;
	assign _01606_ = _00504_ | _03094_;
	assign _01608_ = _01606_ | io_in[7];
	assign _01609_ = _01608_ | _02096_;
	assign _01610_ = io_in[11] & ~_01609_;
	assign _01611_ = _07380_ | _02207_;
	assign _01612_ = _01611_ | io_in[9];
	assign _01613_ = _01612_ | io_in[10];
	assign _01614_ = _01985_ & ~_01613_;
	assign _01615_ = _01283_ | _02207_;
	assign _01616_ = io_in[8] & ~_01615_;
	assign _01617_ = _01386_ | io_in[6];
	assign _01619_ = _01617_ | io_in[7];
	assign _01620_ = _01619_ | _02096_;
	assign _01621_ = io_in[10] & ~_01620_;
	assign _01622_ = _01234_ | io_in[6];
	assign _01623_ = _01622_ | _02207_;
	assign _01624_ = _01623_ | io_in[8];
	assign _01625_ = _01624_ | io_in[10];
	assign _01626_ = _01985_ & ~_01625_;
	assign _01627_ = _01072_ | _03094_;
	assign _01628_ = _01627_ | io_in[6];
	assign _01630_ = _02207_ & ~_01628_;
	assign _01631_ = _00281_ | io_in[6];
	assign _01632_ = _01631_ | _02207_;
	assign _01633_ = _01632_ | _01208_;
	assign _01634_ = _01633_ | _02096_;
	assign _01635_ = _06310_ & ~_01634_;
	assign _01636_ = _02539_ | _03759_;
	assign _01637_ = _01636_ | _02207_;
	assign _01638_ = _01637_ | io_in[8];
	assign _01639_ = _01638_ | io_in[9];
	assign _01641_ = io_in[10] & ~_01639_;
	assign _01642_ = _07510_ | _07422_;
	assign _01643_ = _01642_ | io_in[8];
	assign _01644_ = _01643_ | _02096_;
	assign _01645_ = _01644_ | io_in[10];
	assign _01646_ = _01985_ & ~_01645_;
	assign _01647_ = _01260_ | io_in[6];
	assign _01648_ = _01647_ | _06310_;
	assign _01649_ = io_in[11] & ~_01648_;
	assign _01650_ = _01007_ | io_in[7];
	assign _01653_ = _01650_ | _01208_;
	assign _01654_ = _01653_ | _02096_;
	assign _01655_ = _01654_ | _06310_;
	assign _01656_ = _01985_ & ~_01655_;
	assign _01657_ = _01125_ | io_in[5];
	assign _01658_ = _01657_ | _03759_;
	assign _01659_ = _01658_ | _01208_;
	assign _01660_ = _01659_ | _02096_;
	assign _01661_ = _01660_ | _06310_;
	assign _01662_ = io_in[11] & ~_01661_;
	assign _01664_ = _00989_ | io_in[8];
	assign _01665_ = io_in[10] & ~_01664_;
	assign _01666_ = _07455_ | _03759_;
	assign _01667_ = _01666_ | _02207_;
	assign _01668_ = _01667_ | _01208_;
	assign _01669_ = _01668_ | _02096_;
	assign _01670_ = io_in[10] & ~_01669_;
	assign _01671_ = _07499_ | _03094_;
	assign _01672_ = _01671_ | _03759_;
	assign _01673_ = _01672_ | _02207_;
	assign _01675_ = _01673_ | io_in[8];
	assign _01676_ = io_in[11] & ~_01675_;
	assign _01677_ = _01017_ | io_in[8];
	assign _01678_ = _01677_ | io_in[9];
	assign _01679_ = io_in[11] & ~_01678_;
	assign _01680_ = _01484_ | _01208_;
	assign _01681_ = _01680_ | io_in[10];
	assign _01682_ = io_in[11] & ~_01681_;
	assign _01683_ = _01200_ | _03094_;
	assign _01684_ = _01683_ | io_in[6];
	assign _01686_ = _01684_ | _02207_;
	assign _01687_ = io_in[11] & ~_01686_;
	assign _01688_ = _00533_ | _06310_;
	assign _01689_ = io_in[11] & ~_01688_;
	assign _01690_ = _02994_ | io_in[7];
	assign _01691_ = _01690_ | _06310_;
	assign _01692_ = io_in[11] & ~_01691_;
	assign _01693_ = _01348_ | _01208_;
	assign _01694_ = _01693_ | _02096_;
	assign _01695_ = _01694_ | _06310_;
	assign _01697_ = _01985_ & ~_01695_;
	assign _01698_ = _00757_ | io_in[4];
	assign _01699_ = _01698_ | _01208_;
	assign _01700_ = _01699_ | io_in[9];
	assign _01701_ = _01700_ | io_in[10];
	assign _01702_ = _01985_ & ~_01701_;
	assign _01703_ = _07302_ | _03759_;
	assign _01704_ = _01703_ | io_in[7];
	assign _01705_ = _01704_ | _01208_;
	assign _01706_ = _01705_ | _02096_;
	assign _01708_ = _01706_ | _06310_;
	assign _01709_ = _01985_ & ~_01708_;
	assign _01710_ = _01038_ | io_in[6];
	assign _01711_ = _01710_ | _02207_;
	assign _01712_ = _01711_ | io_in[8];
	assign _01713_ = _02096_ & ~_01712_;
	assign _01714_ = _00521_ | io_in[5];
	assign _01715_ = _01714_ | _02207_;
	assign _01716_ = _01715_ | io_in[8];
	assign _01717_ = _01716_ | io_in[9];
	assign _01719_ = io_in[11] & ~_01717_;
	assign _01720_ = _00521_ | _03094_;
	assign _01721_ = _01720_ | _03759_;
	assign _01722_ = _01721_ | io_in[7];
	assign _01723_ = _01722_ | _01208_;
	assign _01724_ = io_in[11] & ~_01723_;
	assign _01725_ = _01225_ | _03759_;
	assign _01726_ = _01725_ | _01208_;
	assign _01727_ = _01726_ | io_in[10];
	assign _01728_ = io_in[11] & ~_01727_;
	assign _01730_ = _00250_ | io_in[6];
	assign _01731_ = _01730_ | _02207_;
	assign _01732_ = _01731_ | _01208_;
	assign _01733_ = _01732_ | io_in[9];
	assign _01734_ = io_in[10] & ~_01733_;
	assign _01735_ = _00504_ | io_in[5];
	assign _01736_ = _01735_ | _03759_;
	assign _01737_ = _01736_ | _02207_;
	assign _01738_ = _01737_ | io_in[8];
	assign _01739_ = _01738_ | io_in[9];
	assign _01741_ = io_in[11] & ~_01739_;
	assign _01742_ = _01544_ | io_in[8];
	assign _01743_ = _01742_ | _02096_;
	assign _01744_ = io_in[10] & ~_01743_;
	assign _01745_ = _03315_ | io_in[6];
	assign _01746_ = _01745_ | _02207_;
	assign _01747_ = _01746_ | io_in[8];
	assign _01748_ = _01747_ | _02096_;
	assign _01749_ = io_in[10] & ~_01748_;
	assign _01750_ = _01583_ | io_in[6];
	assign _01752_ = _01750_ | io_in[7];
	assign _01753_ = _01752_ | _02096_;
	assign _01754_ = io_in[11] & ~_01753_;
	assign _01755_ = _01312_ | io_in[8];
	assign _01756_ = _06310_ & ~_01755_;
	assign _01757_ = _00694_ | _07422_;
	assign _01758_ = _01757_ | io_in[7];
	assign _01759_ = _01758_ | _01208_;
	assign _01760_ = _01759_ | _02096_;
	assign _01761_ = _01760_ | _06310_;
	assign _01764_ = _01985_ & ~_01761_;
	assign _01765_ = _07362_ | io_in[6];
	assign _01766_ = _01765_ | io_in[7];
	assign _01767_ = _01766_ | io_in[8];
	assign _01768_ = _01767_ | _02096_;
	assign _01769_ = io_in[10] & ~_01768_;
	assign _01770_ = _02539_ | io_in[6];
	assign _01771_ = _01770_ | _02207_;
	assign _01772_ = _01771_ | _01208_;
	assign _01773_ = _01772_ | _02096_;
	assign _01775_ = _01773_ | _06310_;
	assign _01776_ = _01985_ & ~_01775_;
	assign _01777_ = _01642_ | _02207_;
	assign _01778_ = _01777_ | io_in[8];
	assign _01779_ = _01778_ | io_in[9];
	assign _01780_ = io_in[10] & ~_01779_;
	assign _01781_ = _01405_ | _02207_;
	assign _01782_ = _01781_ | io_in[8];
	assign _01783_ = _01782_ | io_in[9];
	assign _01784_ = io_in[10] & ~_01783_;
	assign _01786_ = _05989_ | _03759_;
	assign _01787_ = _01786_ | _02207_;
	assign _01788_ = _01787_ | io_in[8];
	assign _01789_ = io_in[10] & ~_01788_;
	assign _01790_ = _01190_ | _02207_;
	assign _01791_ = _01790_ | io_in[8];
	assign _01792_ = _01791_ | _02096_;
	assign _01793_ = io_in[10] & ~_01792_;
	assign _01794_ = _06865_ | io_in[6];
	assign _01795_ = _01794_ | io_in[7];
	assign _01797_ = _01795_ | _01208_;
	assign _01798_ = _01797_ | io_in[9];
	assign _01799_ = io_in[10] & ~_01798_;
	assign _01800_ = _04524_ | _03759_;
	assign _01801_ = _01800_ | io_in[7];
	assign _01802_ = _01801_ | _06310_;
	assign _01803_ = io_in[11] & ~_01802_;
	assign _01804_ = _07428_ | _02207_;
	assign _01805_ = _01804_ | _06310_;
	assign _01806_ = io_in[11] & ~_01805_;
	assign _01808_ = _00496_ | _03759_;
	assign _01809_ = _01808_ | _02207_;
	assign _01810_ = _01809_ | io_in[9];
	assign _01811_ = _01810_ | io_in[10];
	assign _01812_ = _01985_ & ~_01811_;
	assign _01813_ = _01017_ | _03759_;
	assign _01814_ = _01813_ | io_in[7];
	assign _01815_ = _01814_ | _02096_;
	assign _01816_ = _01985_ & ~_01815_;
	assign _01817_ = _07510_ | io_in[6];
	assign _01819_ = _01817_ | io_in[8];
	assign _01820_ = _01819_ | _02096_;
	assign _01821_ = _01820_ | io_in[10];
	assign _01822_ = _01985_ & ~_01821_;
	assign _01823_ = _07031_ | io_in[5];
	assign _01824_ = _01823_ | io_in[6];
	assign _01825_ = _01824_ | io_in[7];
	assign _01826_ = _01825_ | _06310_;
	assign _01827_ = io_in[11] & ~_01826_;
	assign _01828_ = _00135_ | _02207_;
	assign _01830_ = _01828_ | _02096_;
	assign _01831_ = _01830_ | io_in[10];
	assign _01832_ = _01985_ & ~_01831_;
	assign _01833_ = _00889_ | io_in[5];
	assign _01834_ = _01833_ | _03759_;
	assign _01835_ = _01834_ | io_in[7];
	assign _01836_ = _01835_ | _01208_;
	assign _01837_ = _01836_ | _02096_;
	assign _01838_ = io_in[10] & ~_01837_;
	assign _01839_ = _00986_ | _03759_;
	assign _01841_ = _01839_ | _02207_;
	assign _01842_ = _01841_ | io_in[8];
	assign _01843_ = _01842_ | io_in[10];
	assign _01844_ = _01985_ & ~_01843_;
	assign _01845_ = _07383_ | _03759_;
	assign _01846_ = _01845_ | _02207_;
	assign _01847_ = _01846_ | _06310_;
	assign _01848_ = io_in[11] & ~_01847_;
	assign _01849_ = _00521_ | io_in[4];
	assign _01850_ = _01849_ | _03759_;
	assign _01852_ = _01850_ | _02207_;
	assign _01853_ = _01852_ | io_in[8];
	assign _01854_ = _01853_ | _02096_;
	assign _01855_ = _06310_ & ~_01854_;
	assign _01856_ = _01386_ | _03759_;
	assign _01857_ = _01856_ | _02207_;
	assign _01858_ = _01857_ | io_in[8];
	assign _01859_ = io_in[9] & ~_01858_;
	assign _01860_ = _01266_ | io_in[7];
	assign _01861_ = _01860_ | _02096_;
	assign _01863_ = io_in[11] & ~_01861_;
	assign _01864_ = _01225_ | io_in[5];
	assign _01865_ = _01864_ | _03759_;
	assign _01866_ = _01865_ | io_in[7];
	assign _01867_ = _01866_ | _01208_;
	assign _01868_ = _01867_ | _02096_;
	assign _01869_ = io_in[10] & ~_01868_;
	assign _01870_ = _01404_ | io_in[5];
	assign _01871_ = _01870_ | io_in[6];
	assign _01872_ = _01871_ | _02207_;
	assign _01875_ = _01872_ | io_in[8];
	assign _01876_ = _01875_ | _02096_;
	assign _01877_ = io_in[10] & ~_01876_;
	assign _01878_ = _01031_ | _07422_;
	assign _01879_ = _01878_ | _03759_;
	assign _01880_ = _01879_ | io_in[7];
	assign _01881_ = _01880_ | io_in[8];
	assign _01882_ = _01881_ | io_in[9];
	assign _01883_ = io_in[10] & ~_01882_;
	assign _01884_ = _00443_ | io_in[6];
	assign _01886_ = _01884_ | _02207_;
	assign _01887_ = _01886_ | io_in[8];
	assign _01888_ = _01887_ | _02096_;
	assign _01889_ = io_in[10] & ~_01888_;
	assign _01890_ = _01115_ | _03759_;
	assign _01891_ = _01890_ | _02207_;
	assign _01892_ = _01891_ | io_in[9];
	assign _01893_ = io_in[11] & ~_01892_;
	assign _01894_ = _07413_ | io_in[7];
	assign _01895_ = _01894_ | io_in[9];
	assign _01897_ = io_in[10] & ~_01895_;
	assign _01898_ = _07255_ | _03094_;
	assign _01899_ = _01898_ | io_in[7];
	assign _01900_ = _01899_ | _06310_;
	assign _01901_ = io_in[11] & ~_01900_;
	assign _01902_ = _07336_ | _03759_;
	assign _01903_ = _01902_ | io_in[7];
	assign _01904_ = _01903_ | io_in[8];
	assign _01905_ = io_in[11] & ~_01904_;
	assign _01906_ = _06942_ | _03759_;
	assign _01908_ = _01906_ | _02207_;
	assign _01909_ = _01208_ & ~_01908_;
	assign _01910_ = _07251_ | _02207_;
	assign _01911_ = _01910_ | _01208_;
	assign _01912_ = _01911_ | _02096_;
	assign _01913_ = _06310_ & ~_01912_;
	assign _01914_ = _01864_ | io_in[7];
	assign _01915_ = _01914_ | io_in[8];
	assign _01916_ = _01915_ | io_in[9];
	assign _01917_ = io_in[11] & ~_01916_;
	assign _01919_ = _01200_ | io_in[5];
	assign _01920_ = _01919_ | io_in[6];
	assign _01921_ = _01920_ | _02207_;
	assign _01922_ = _01921_ | io_in[8];
	assign _01923_ = _01922_ | io_in[9];
	assign _01924_ = io_in[10] & ~_01923_;
	assign _01925_ = _01484_ | io_in[7];
	assign _01926_ = _01925_ | _01208_;
	assign _01927_ = _01926_ | _06310_;
	assign _01928_ = _01985_ & ~_01927_;
	assign _01930_ = _06864_ | io_in[6];
	assign _01931_ = _01930_ | _02207_;
	assign _01932_ = _01931_ | _01208_;
	assign _01933_ = _01932_ | io_in[9];
	assign _01934_ = io_in[11] & ~_01933_;
	assign _01935_ = _01770_ | io_in[7];
	assign _01936_ = _01935_ | _01208_;
	assign _01937_ = _01936_ | io_in[9];
	assign _01938_ = io_in[10] & ~_01937_;
	assign _01939_ = _00170_ | _02096_;
	assign _01941_ = _01939_ | _06310_;
	assign _01942_ = _01985_ & ~_01941_;
	assign _01943_ = _01721_ | _02207_;
	assign _01944_ = _01943_ | _02096_;
	assign _01945_ = _01985_ & ~_01944_;
	assign _01946_ = _06720_ | io_in[6];
	assign _01947_ = _01946_ | io_in[7];
	assign _01948_ = _01947_ | _01208_;
	assign _01949_ = _01948_ | io_in[10];
	assign _01950_ = io_in[11] & ~_01949_;
	assign _01952_ = _01505_ | _06310_;
	assign _01953_ = io_in[11] & ~_01952_;
	assign _01954_ = _01427_ | _02207_;
	assign _01955_ = _01954_ | io_in[8];
	assign _01956_ = _01955_ | _02096_;
	assign _01957_ = io_in[10] & ~_01956_;
	assign _01958_ = _07362_ | io_in[5];
	assign _01959_ = _01958_ | io_in[6];
	assign _01960_ = _01959_ | _02207_;
	assign _01961_ = _01960_ | io_in[9];
	assign _01963_ = io_in[10] & ~_01961_;
	assign _01964_ = _01406_ | io_in[7];
	assign _01965_ = _01964_ | io_in[8];
	assign _01966_ = io_in[9] & ~_01965_;
	assign _01967_ = _00759_ | _01208_;
	assign _01968_ = _01967_ | io_in[9];
	assign _01969_ = io_in[11] & ~_01968_;
	assign _01970_ = _00504_ | _03759_;
	assign _01971_ = _01970_ | io_in[7];
	assign _01972_ = _01971_ | io_in[8];
	assign _01974_ = _01972_ | io_in[9];
	assign _01975_ = io_in[10] & ~_01974_;
	assign _01976_ = _01260_ | _03759_;
	assign _01977_ = _01976_ | _02207_;
	assign _01978_ = _01977_ | _01208_;
	assign _01979_ = _02096_ & ~_01978_;
	assign _01980_ = _01906_ | io_in[8];
	assign _01981_ = _01985_ & ~_01980_;
	assign _01982_ = _01698_ | io_in[5];
	assign _01983_ = _01982_ | _03759_;
	assign _01986_ = _01983_ | io_in[7];
	assign _01987_ = _01986_ | _01208_;
	assign _01988_ = _01987_ | _02096_;
	assign _01989_ = _01985_ & ~_01988_;
	assign _01990_ = _01031_ | _03094_;
	assign _01991_ = _01990_ | io_in[7];
	assign _01992_ = _01991_ | _01208_;
	assign _01993_ = _01992_ | io_in[9];
	assign _01994_ = io_in[11] & ~_01993_;
	assign _01995_ = _03216_ | io_in[7];
	assign _01997_ = _01995_ | _01208_;
	assign _01998_ = _01997_ | io_in[9];
	assign _01999_ = io_in[10] & ~_01998_;
	assign _02000_ = _00720_ | _03759_;
	assign _02001_ = _02000_ | _01208_;
	assign _02002_ = _02001_ | _02096_;
	assign _02003_ = _06310_ & ~_02002_;
	assign _02004_ = _07402_ | _03759_;
	assign _02005_ = _02004_ | _02207_;
	assign _02006_ = _02005_ | io_in[8];
	assign _02008_ = _02006_ | io_in[9];
	assign _02009_ = io_in[11] & ~_02008_;
	assign _02010_ = _03870_ | io_in[4];
	assign _02011_ = _02010_ | io_in[5];
	assign _02012_ = _02011_ | io_in[6];
	assign _02013_ = _02012_ | io_in[7];
	assign _02014_ = _02013_ | _01208_;
	assign _02015_ = _02014_ | _02096_;
	assign _02016_ = _02015_ | _06310_;
	assign _02017_ = io_in[11] & ~_02016_;
	assign _02019_ = _00521_ | io_in[6];
	assign _02020_ = _02019_ | _02207_;
	assign _02021_ = _02020_ | _01208_;
	assign _02022_ = _02021_ | _06310_;
	assign _02023_ = _01985_ & ~_02022_;
	assign _02024_ = _01451_ | io_in[8];
	assign _02025_ = _02024_ | _02096_;
	assign _02026_ = io_in[10] & ~_02025_;
	assign _02027_ = _06310_ & ~_00601_;
	assign _02028_ = (io_in[11] ? _02027_ : _02026_);
	assign _02030_ = _02028_ | _02023_;
	assign _02031_ = _02030_ | _02017_;
	assign _02032_ = _02031_ | _02009_;
	assign _02033_ = _02032_ | _02003_;
	assign _02034_ = _02033_ | _01999_;
	assign _02035_ = _02034_ | _01994_;
	assign _02036_ = _02035_ | _01989_;
	assign _02037_ = _02036_ | _01981_;
	assign _02038_ = _02037_ | _01979_;
	assign _02039_ = _02038_ | _01975_;
	assign _02041_ = _02039_ | _01969_;
	assign _02042_ = _02041_ | _01966_;
	assign _02043_ = _02042_ | _01963_;
	assign _02044_ = _02043_ | _01957_;
	assign _02045_ = _02044_ | _01953_;
	assign _02046_ = _02045_ | _01950_;
	assign _02047_ = _02046_ | _01945_;
	assign _02048_ = _02047_ | _01942_;
	assign _02049_ = _02048_ | _01938_;
	assign _02050_ = _02049_ | _01934_;
	assign _02052_ = _02050_ | _01928_;
	assign _02053_ = _02052_ | _01924_;
	assign _02054_ = _02053_ | _01917_;
	assign _02055_ = _02054_ | _01913_;
	assign _02056_ = _02055_ | _01909_;
	assign _02057_ = _02056_ | _01905_;
	assign _02058_ = _02057_ | _01901_;
	assign _02059_ = _02058_ | _01897_;
	assign _02060_ = _02059_ | _01893_;
	assign _02061_ = _02060_ | _01889_;
	assign _02063_ = _02061_ | _01883_;
	assign _02064_ = _02063_ | _01877_;
	assign _02065_ = _02064_ | _01869_;
	assign _02066_ = _02065_ | _01863_;
	assign _02067_ = _02066_ | _01859_;
	assign _02068_ = _02067_ | _01855_;
	assign _02069_ = _02068_ | _01848_;
	assign _02070_ = _02069_ | _01844_;
	assign _02071_ = _02070_ | _01838_;
	assign _02072_ = _02071_ | _01832_;
	assign _02074_ = _02072_ | _01827_;
	assign _02075_ = _02074_ | _01822_;
	assign _02076_ = _02075_ | _01816_;
	assign _02077_ = _02076_ | _01812_;
	assign _02078_ = _02077_ | _01806_;
	assign _02079_ = _02078_ | _01803_;
	assign _02080_ = _02079_ | _01799_;
	assign _02081_ = _02080_ | _01793_;
	assign _02082_ = _02081_ | _01789_;
	assign _02083_ = _02082_ | _01784_;
	assign _02085_ = _02083_ | _01780_;
	assign _02086_ = _02085_ | _01776_;
	assign _02087_ = _02086_ | _01769_;
	assign _02088_ = _02087_ | _01764_;
	assign _02089_ = _02088_ | _01756_;
	assign _02090_ = _02089_ | _01754_;
	assign _02091_ = _02090_ | _01749_;
	assign _02092_ = _02091_ | _01744_;
	assign _02093_ = _02092_ | _01741_;
	assign _02094_ = _02093_ | _01734_;
	assign _02097_ = _02094_ | _01728_;
	assign _02098_ = _02097_ | _01724_;
	assign _02099_ = _02098_ | _01719_;
	assign _02100_ = _02099_ | _01713_;
	assign _02101_ = _02100_ | _01709_;
	assign _02102_ = _02101_ | _01702_;
	assign _02103_ = _02102_ | _01697_;
	assign _02104_ = _02103_ | _01692_;
	assign _02105_ = _02104_ | _01689_;
	assign _02106_ = _02105_ | _01687_;
	assign _02108_ = _02106_ | _01682_;
	assign _02109_ = _02108_ | _01679_;
	assign _02110_ = _02109_ | _01676_;
	assign _02111_ = _02110_ | _01670_;
	assign _02112_ = _02111_ | _01665_;
	assign _02113_ = _02112_ | _01662_;
	assign _02114_ = _02113_ | _01656_;
	assign _02115_ = _02114_ | _01649_;
	assign _02116_ = _02115_ | _01646_;
	assign _02117_ = _02116_ | _01641_;
	assign _02119_ = _02117_ | _01635_;
	assign _02120_ = _02119_ | _01630_;
	assign _02121_ = _02120_ | _01626_;
	assign _02122_ = _02121_ | _01621_;
	assign _02123_ = _02122_ | _01616_;
	assign _02124_ = _02123_ | _01614_;
	assign _02125_ = _02124_ | _01610_;
	assign _02126_ = _02125_ | _01605_;
	assign _02127_ = _02126_ | _01600_;
	assign _02128_ = _02127_ | _01593_;
	assign _02130_ = _02128_ | _01588_;
	assign _02131_ = _02130_ | _01582_;
	assign _02132_ = _02131_ | _01579_;
	assign _02133_ = _02132_ | _01577_;
	assign _02134_ = _02133_ | _01572_;
	assign _02135_ = _02134_ | _01567_;
	assign _02136_ = _02135_ | _01562_;
	assign _02137_ = _02136_ | _01556_;
	assign _02138_ = _02137_ | _01551_;
	assign _02139_ = _02138_ | _01546_;
	assign _02141_ = _02139_ | _01543_;
	assign _02142_ = _02141_ | _01536_;
	assign _02143_ = _02142_ | _01533_;
	assign _02144_ = _02143_ | _01530_;
	assign _02145_ = _02144_ | _01525_;
	assign _02146_ = _02145_ | _01520_;
	assign _02147_ = _02146_ | _01514_;
	assign _02148_ = _02147_ | _01509_;
	assign _02149_ = _02148_ | _01504_;
	assign _02150_ = _02149_ | _01499_;
	assign _02152_ = _02150_ | _01497_;
	assign _02153_ = _02152_ | _01493_;
	assign _02154_ = _02153_ | _01489_;
	assign _02155_ = _02154_ | _01482_;
	assign _02156_ = _02155_ | _01479_;
	assign _02157_ = _02156_ | _01473_;
	assign _02158_ = _02157_ | _01468_;
	assign _02159_ = _02158_ | _01465_;
	assign _02160_ = _02159_ | _01459_;
	assign _02161_ = _02160_ | _01455_;
	assign _02163_ = _02161_ | _01450_;
	assign _02164_ = _02163_ | _01447_;
	assign _02165_ = _02164_ | _01444_;
	assign _02166_ = _02165_ | _01437_;
	assign _02167_ = _02166_ | _01433_;
	assign _02168_ = _02167_ | _01426_;
	assign _02169_ = _02168_ | _01420_;
	assign _02170_ = _02169_ | _01415_;
	assign _02171_ = _02170_ | _01410_;
	assign _02172_ = _02171_ | _01403_;
	assign _02174_ = _02172_ | _01399_;
	assign _02175_ = _02174_ | _01394_;
	assign _02176_ = _02175_ | _01390_;
	assign _02177_ = _02176_ | _01384_;
	assign _02178_ = _02177_ | _01379_;
	assign _02179_ = _02178_ | _01375_;
	assign _02180_ = _02179_ | _01370_;
	assign _02181_ = _02180_ | _01365_;
	assign _02182_ = _02181_ | _01359_;
	assign _02183_ = _02182_ | _01353_;
	assign _02185_ = _02183_ | _01347_;
	assign _02186_ = _02185_ | _01339_;
	assign _02187_ = _02186_ | _01333_;
	assign _02188_ = _02187_ | _01329_;
	assign _02189_ = _02188_ | _01326_;
	assign _02190_ = _02189_ | _01320_;
	assign _02191_ = _02190_ | _01313_;
	assign _02192_ = _02191_ | _01311_;
	assign _02193_ = _02192_ | _01305_;
	assign _02194_ = _02193_ | _01301_;
	assign _02196_ = _02194_ | _01298_;
	assign _02197_ = _02196_ | _01293_;
	assign _02198_ = _02197_ | _01290_;
	assign _02199_ = _02198_ | _01287_;
	assign _02200_ = _02199_ | _01281_;
	assign _02201_ = _02200_ | _01276_;
	assign _02202_ = _02201_ | _01271_;
	assign _02203_ = _02202_ | _01269_;
	assign _02204_ = _02203_ | _01265_;
	assign _02205_ = _02204_ | _01259_;
	assign _02208_ = _02205_ | _01256_;
	assign _02209_ = _02208_ | _01250_;
	assign _02210_ = _02209_ | _01245_;
	assign _02211_ = _02210_ | _01240_;
	assign _02212_ = _02211_ | _01233_;
	assign _02213_ = _02212_ | _01231_;
	assign _02214_ = _02213_ | _01224_;
	assign _02215_ = _02214_ | _01218_;
	assign _02216_ = _02215_ | _01212_;
	assign _02217_ = _02216_ | _01205_;
	assign _02219_ = _02217_ | _01199_;
	assign _02220_ = _02219_ | _01194_;
	assign _02221_ = _02220_ | _01189_;
	assign _02222_ = _02221_ | _01183_;
	assign _02223_ = _02222_ | _01179_;
	assign _02224_ = _02223_ | _01171_;
	assign _02225_ = _02224_ | _01167_;
	assign _02226_ = _02225_ | _01161_;
	assign _02227_ = _02226_ | _01156_;
	assign _02228_ = _02227_ | _01153_;
	assign _02230_ = _02228_ | _01147_;
	assign _02231_ = _02230_ | _01142_;
	assign _02232_ = _02231_ | _01137_;
	assign _02233_ = _02232_ | _01132_;
	assign _02234_ = _02233_ | _01124_;
	assign _02235_ = _02234_ | _01120_;
	assign _02236_ = _02235_ | _01114_;
	assign _02237_ = _02236_ | _01110_;
	assign _02238_ = _02237_ | _01104_;
	assign _02239_ = _02238_ | _01100_;
	assign _02241_ = _02239_ | _01095_;
	assign _02242_ = _02241_ | _01091_;
	assign _02243_ = _02242_ | _01088_;
	assign _02244_ = _02243_ | _01083_;
	assign _02245_ = _02244_ | _01078_;
	assign _02246_ = _02245_ | _01071_;
	assign _02247_ = _02246_ | _01065_;
	assign _02248_ = _02247_ | _01056_;
	assign _02249_ = _02248_ | _01050_;
	assign _02250_ = _02249_ | _01045_;
	assign _02252_ = _02250_ | _01037_;
	assign _02253_ = _02252_ | _01034_;
	assign _02254_ = _02253_ | _01028_;
	assign _02255_ = _02254_ | _01023_;
	assign _02256_ = _02255_ | _01016_;
	assign _02257_ = _02256_ | _01012_;
	assign _02258_ = _02257_ | _01005_;
	assign _02259_ = _02258_ | _01000_;
	assign _02260_ = _02259_ | _00996_;
	assign _02261_ = _02260_ | _00992_;
	assign _02263_ = _02261_ | _00984_;
	assign \mchip.val [4] = _02263_ | _00978_;
	assign _02264_ = _01865_ | _02207_;
	assign _02265_ = _02264_ | io_in[9];
	assign _02266_ = _01985_ & ~_02265_;
	assign _02267_ = _01878_ | _03094_;
	assign _02268_ = _02267_ | io_in[6];
	assign _02269_ = _02207_ & ~_02268_;
	assign _02270_ = _01794_ | io_in[8];
	assign _02271_ = _02270_ | _02096_;
	assign _02273_ = _02271_ | io_in[10];
	assign _02274_ = _01985_ & ~_02273_;
	assign _02275_ = _01391_ | _01208_;
	assign _02276_ = _02275_ | _02096_;
	assign _02277_ = _02276_ | _06310_;
	assign _02278_ = _01985_ & ~_02277_;
	assign _02279_ = io_in[11] & ~_06000_;
	assign _02280_ = _01344_ | _02096_;
	assign _02281_ = _01985_ & ~_02280_;
	assign _02282_ = _01480_ | io_in[9];
	assign _02284_ = io_in[11] & ~_02282_;
	assign _02285_ = _01404_ | io_in[4];
	assign _02286_ = _02285_ | _03759_;
	assign _02287_ = _02286_ | io_in[7];
	assign _02288_ = _02287_ | _01208_;
	assign _02289_ = _02288_ | _02096_;
	assign _02290_ = _01985_ & ~_02289_;
	assign _02291_ = _02350_ | _01208_;
	assign _02292_ = _02291_ | _02096_;
	assign _02293_ = _02292_ | _06310_;
	assign _02295_ = _01985_ & ~_02293_;
	assign _02296_ = _00481_ | _02207_;
	assign _02297_ = _02296_ | _06310_;
	assign _02298_ = io_in[11] & ~_02297_;
	assign _02299_ = _01671_ | _01208_;
	assign _02300_ = _02096_ & ~_02299_;
	assign _02301_ = _00514_ | _02207_;
	assign _02302_ = _02301_ | _01208_;
	assign _02303_ = _02096_ & ~_02302_;
	assign _02304_ = _07412_ | _02207_;
	assign _02306_ = _02304_ | io_in[9];
	assign _02307_ = _06310_ & ~_02306_;
	assign _02308_ = _07412_ | io_in[6];
	assign _02309_ = _02308_ | _02207_;
	assign _02310_ = _02309_ | _01208_;
	assign _02311_ = io_in[10] & ~_02310_;
	assign _02312_ = _00439_ | io_in[6];
	assign _02313_ = _02312_ | io_in[8];
	assign _02314_ = _02313_ | _02096_;
	assign _02315_ = _02314_ | io_in[10];
	assign _02318_ = _01985_ & ~_02315_;
	assign _02319_ = _01714_ | io_in[6];
	assign _02320_ = _02319_ | io_in[8];
	assign _02321_ = _02320_ | io_in[9];
	assign _02322_ = io_in[10] & ~_02321_;
	assign _02323_ = _02539_ | io_in[5];
	assign _02324_ = _02323_ | _03759_;
	assign _02325_ = _02324_ | _02207_;
	assign _02326_ = _02325_ | io_in[8];
	assign _02327_ = io_in[11] & ~_02326_;
	assign _02329_ = _01175_ | io_in[7];
	assign _02330_ = _02329_ | _01208_;
	assign _02331_ = _02330_ | _06310_;
	assign _02332_ = _01985_ & ~_02331_;
	assign _02333_ = _01986_ | _02096_;
	assign _02334_ = io_in[11] & ~_02333_;
	assign _02335_ = _01401_ | io_in[8];
	assign _02336_ = _02335_ | _02096_;
	assign _02337_ = io_in[11] & ~_02336_;
	assign _02338_ = io_in[9] & ~_01292_;
	assign _02340_ = _01475_ | _03759_;
	assign _02341_ = _02340_ | io_in[7];
	assign _02342_ = _02341_ | io_in[9];
	assign _02343_ = io_in[11] & ~_02342_;
	assign _02344_ = _01421_ | _03759_;
	assign _02345_ = _02344_ | _02207_;
	assign _02346_ = _02345_ | io_in[8];
	assign _02347_ = _02346_ | _02096_;
	assign _02348_ = io_in[10] & ~_02347_;
	assign _02349_ = _00985_ | io_in[5];
	assign _02351_ = _02349_ | _03759_;
	assign _02352_ = _02351_ | _02207_;
	assign _02353_ = _02352_ | _01208_;
	assign _02354_ = _06310_ & ~_02353_;
	assign _02355_ = _02272_ | io_in[7];
	assign _02356_ = _02355_ | _01208_;
	assign _02357_ = _02356_ | io_in[9];
	assign _02358_ = _06310_ & ~_02357_;
	assign _02359_ = _01596_ | io_in[6];
	assign _02360_ = _02359_ | _02207_;
	assign _02362_ = _02360_ | io_in[9];
	assign _02363_ = _02362_ | io_in[10];
	assign _02364_ = _01985_ & ~_02363_;
	assign _02365_ = _01990_ | _03759_;
	assign _02366_ = _02365_ | _02207_;
	assign _02367_ = _02366_ | io_in[8];
	assign _02368_ = _02096_ & ~_02367_;
	assign _02369_ = _00360_ | io_in[7];
	assign _02370_ = _02369_ | io_in[8];
	assign _02371_ = io_in[11] & ~_02370_;
	assign _02373_ = _07419_ | _03094_;
	assign _02374_ = _02373_ | io_in[7];
	assign _02375_ = _02374_ | _01208_;
	assign _02376_ = io_in[11] & ~_02375_;
	assign _02377_ = io_in[11] & ~_01393_;
	assign _02378_ = _07304_ | _01208_;
	assign _02379_ = _02378_ | _02096_;
	assign _02380_ = _06310_ & ~_02379_;
	assign _02381_ = _06976_ | _02207_;
	assign _02382_ = _02381_ | _01208_;
	assign _02384_ = io_in[9] & ~_02382_;
	assign _02385_ = _02384_ & ~io_in[11];
	assign _02386_ = _01483_ | io_in[6];
	assign _02387_ = _02386_ | _02096_;
	assign _02388_ = _02387_ | io_in[10];
	assign _02389_ = _01985_ & ~_02388_;
	assign _02390_ = _06065_ | _02207_;
	assign _02391_ = _02390_ | _01208_;
	assign _02392_ = io_in[11] & ~_02391_;
	assign _02393_ = _01647_ | io_in[7];
	assign _02395_ = _01208_ & ~_02393_;
	assign _02396_ = _02395_ & ~_02096_;
	assign _02397_ = _02285_ | _02207_;
	assign _02398_ = _02397_ | _01208_;
	assign _02399_ = _02398_ | io_in[9];
	assign _02400_ = io_in[10] & ~_02399_;
	assign _02401_ = _00333_ | _02207_;
	assign _02402_ = _02401_ | _01208_;
	assign _02403_ = _02402_ | _02096_;
	assign _02404_ = _02403_ | _06310_;
	assign _02406_ = _01985_ & ~_02404_;
	assign _02407_ = _00388_ | io_in[6];
	assign _02408_ = _02407_ | _01208_;
	assign _02409_ = _02408_ | io_in[9];
	assign _02410_ = _02409_ | io_in[10];
	assign _02411_ = _01985_ & ~_02410_;
	assign _02412_ = _01366_ | _02207_;
	assign _02413_ = _02412_ | io_in[8];
	assign _02414_ = _02413_ | io_in[9];
	assign _02415_ = _01985_ & ~_02414_;
	assign _02417_ = _01234_ | _03094_;
	assign _02418_ = _02417_ | _02207_;
	assign _02419_ = _02418_ | _02096_;
	assign _02420_ = _01985_ & ~_02419_;
	assign _02421_ = _02304_ | _01208_;
	assign _02422_ = io_in[11] & ~_02421_;
	assign _02423_ = _01387_ | _01208_;
	assign _02424_ = io_in[11] & ~_02423_;
	assign _02425_ = _04302_ | _02207_;
	assign _02426_ = _02425_ | io_in[8];
	assign _02429_ = _02426_ | io_in[9];
	assign _02430_ = io_in[10] & ~_02429_;
	assign _02431_ = _01092_ | io_in[8];
	assign _02432_ = _02431_ | _02096_;
	assign _02433_ = io_in[10] & ~_02432_;
	assign _02434_ = _01024_ | io_in[7];
	assign _02435_ = _02434_ | io_in[9];
	assign _02436_ = io_in[11] & ~_02435_;
	assign _02437_ = _01864_ | io_in[6];
	assign _02438_ = _02437_ | _02207_;
	assign _02440_ = _02438_ | _01208_;
	assign _02441_ = io_in[11] & ~_02440_;
	assign _02442_ = _01282_ | io_in[6];
	assign _02443_ = _02442_ | _02207_;
	assign _02444_ = _02443_ | _01208_;
	assign _02445_ = io_in[9] & ~_02444_;
	assign _02446_ = _01247_ | io_in[8];
	assign _02447_ = _02446_ | _02096_;
	assign _02448_ = io_in[10] & ~_02447_;
	assign _02449_ = _02319_ | io_in[7];
	assign _02451_ = _02449_ | _01208_;
	assign _02452_ = _02451_ | io_in[9];
	assign _02453_ = _06310_ & ~_02452_;
	assign _02454_ = _00178_ | _02207_;
	assign _02455_ = _02454_ | io_in[8];
	assign _02456_ = _02455_ | io_in[10];
	assign _02457_ = _01985_ & ~_02456_;
	assign _02458_ = _00360_ | _02207_;
	assign _02459_ = _02458_ | io_in[9];
	assign _02460_ = _02459_ | io_in[10];
	assign _02462_ = _01985_ & ~_02460_;
	assign _02463_ = _00900_ | _02207_;
	assign _02464_ = _02463_ | io_in[8];
	assign _02465_ = _02464_ | io_in[9];
	assign _02466_ = _06310_ & ~_02465_;
	assign _02467_ = _00373_ | io_in[6];
	assign _02468_ = _02467_ | io_in[7];
	assign _02469_ = _02468_ | io_in[9];
	assign _02470_ = _01985_ & ~_02469_;
	assign _02471_ = _07378_ | io_in[5];
	assign _02473_ = _02471_ | _02207_;
	assign _02474_ = _02473_ | _01208_;
	assign _02475_ = _02474_ | _02096_;
	assign _02476_ = _06310_ & ~_02475_;
	assign _02477_ = _01983_ | _06310_;
	assign _02478_ = io_in[11] & ~_02477_;
	assign _02479_ = _01864_ | _02207_;
	assign _02480_ = _02479_ | io_in[8];
	assign _02481_ = _02480_ | io_in[9];
	assign _02482_ = io_in[10] & ~_02481_;
	assign _02484_ = _01024_ | io_in[6];
	assign _02485_ = _02484_ | io_in[7];
	assign _02486_ = _02485_ | io_in[9];
	assign _02487_ = io_in[10] & ~_02486_;
	assign _02488_ = _07075_ | io_in[6];
	assign _02489_ = _02488_ | io_in[7];
	assign _02490_ = _02489_ | _01208_;
	assign _02491_ = _02490_ | io_in[9];
	assign _02492_ = _06310_ & ~_02491_;
	assign _02493_ = _01361_ | _02096_;
	assign _02495_ = _02493_ | io_in[10];
	assign _02496_ = _01985_ & ~_02495_;
	assign _02497_ = _00010_ | _03759_;
	assign _02498_ = _02497_ | io_in[8];
	assign _02499_ = _02498_ | io_in[9];
	assign _02500_ = io_in[10] & ~_02499_;
	assign _02501_ = _01006_ | io_in[6];
	assign _02502_ = _02501_ | io_in[8];
	assign _02503_ = _02502_ | io_in[9];
	assign _02504_ = io_in[11] & ~_02503_;
	assign _02506_ = _01672_ | io_in[7];
	assign _02507_ = _02506_ | _02096_;
	assign _02508_ = io_in[11] & ~_02507_;
	assign _02509_ = _05889_ | _03094_;
	assign _02510_ = _02207_ & ~_02509_;
	assign _02511_ = _01307_ | _02207_;
	assign _02512_ = _02511_ | _01208_;
	assign _02513_ = _02512_ | io_in[9];
	assign _02514_ = io_in[11] & ~_02513_;
	assign _02515_ = _02308_ | io_in[7];
	assign _02517_ = _02515_ | io_in[8];
	assign _02518_ = _02096_ & ~_02517_;
	assign _02519_ = _00971_ | io_in[6];
	assign _02520_ = _02519_ | io_in[7];
	assign _02521_ = _02520_ | _01208_;
	assign _02522_ = _02521_ | io_in[9];
	assign _02523_ = io_in[10] & ~_02522_;
	assign _02524_ = _02772_ | io_in[6];
	assign _02525_ = _02524_ | io_in[7];
	assign _02526_ = _02525_ | io_in[8];
	assign _02528_ = io_in[10] & ~_02526_;
	assign _02529_ = _00131_ | io_in[5];
	assign _02530_ = _02529_ | _03759_;
	assign _02531_ = _02530_ | io_in[7];
	assign _02532_ = _02531_ | _02096_;
	assign _02533_ = _02532_ | _06310_;
	assign _02534_ = _01985_ & ~_02533_;
	assign _02535_ = _07186_ | _03759_;
	assign _02536_ = _02535_ | io_in[7];
	assign _02537_ = _02536_ | _01208_;
	assign _02540_ = _02537_ | io_in[9];
	assign _02541_ = io_in[11] & ~_02540_;
	assign _02542_ = _04923_ & ~_01985_;
	assign _02543_ = _03992_ | io_in[5];
	assign _02544_ = _02543_ | _03759_;
	assign _02545_ = _02544_ | _02207_;
	assign _02546_ = _02545_ | io_in[8];
	assign _02547_ = _02546_ | io_in[9];
	assign _02548_ = io_in[10] & ~_02547_;
	assign _02549_ = _07410_ | _03759_;
	assign _02551_ = _02549_ | io_in[7];
	assign _02552_ = _02551_ | _01208_;
	assign _02553_ = _06310_ & ~_02552_;
	assign _02554_ = _02553_ & ~io_in[11];
	assign _02555_ = _07271_ | io_in[6];
	assign _02556_ = _02555_ | _01208_;
	assign _02557_ = _02556_ | io_in[9];
	assign _02558_ = io_in[10] & ~_02557_;
	assign _02559_ = _01632_ | io_in[8];
	assign _02560_ = _02559_ | io_in[9];
	assign _02562_ = io_in[10] & ~_02560_;
	assign _02563_ = _00540_ | _01208_;
	assign _02564_ = _02563_ | io_in[9];
	assign _02565_ = _02564_ | io_in[10];
	assign _02566_ = _01985_ & ~_02565_;
	assign _02567_ = _00360_ | _03759_;
	assign _02568_ = _02567_ | io_in[7];
	assign _02569_ = _02568_ | io_in[10];
	assign _02570_ = io_in[11] & ~_02569_;
	assign _02571_ = _01007_ | _03759_;
	assign _02573_ = _02571_ | io_in[7];
	assign _02574_ = _02573_ | _01208_;
	assign _02575_ = _06310_ & ~_02574_;
	assign _02576_ = _01416_ | io_in[7];
	assign _02577_ = _02576_ | _01208_;
	assign _02578_ = _02577_ | _02096_;
	assign _02579_ = _02578_ | _06310_;
	assign _02580_ = _01985_ & ~_02579_;
	assign _02581_ = _01505_ | io_in[8];
	assign _02582_ = _02581_ | _02096_;
	assign _02584_ = io_in[10] & ~_02582_;
	assign _02585_ = _01642_ | _03759_;
	assign _02586_ = _02585_ | io_in[7];
	assign _02587_ = _02586_ | io_in[10];
	assign _02588_ = io_in[11] & ~_02587_;
	assign _02589_ = _01215_ | _01208_;
	assign _02590_ = _02589_ | _02096_;
	assign _02591_ = io_in[10] & ~_02590_;
	assign _02592_ = _00986_ | io_in[7];
	assign _02593_ = _02592_ | _01208_;
	assign _02595_ = _02593_ | io_in[9];
	assign _02596_ = io_in[11] & ~_02595_;
	assign _02597_ = _01024_ | _02207_;
	assign _02598_ = _02597_ | io_in[8];
	assign _02599_ = io_in[11] & ~_02598_;
	assign _02600_ = _01910_ | io_in[8];
	assign _02601_ = io_in[10] & ~_02600_;
	assign _02602_ = _01817_ | io_in[7];
	assign _02603_ = _02602_ | _01208_;
	assign _02604_ = _02603_ | io_in[9];
	assign _02606_ = io_in[10] & ~_02604_;
	assign _02607_ = _00694_ | _01208_;
	assign _02608_ = _02607_ | io_in[9];
	assign _02609_ = _02608_ | io_in[10];
	assign _02610_ = _01985_ & ~_02609_;
	assign _02611_ = _06143_ | io_in[8];
	assign _02612_ = _02611_ | _02096_;
	assign _02613_ = io_in[10] & ~_02612_;
	assign _02614_ = _01595_ | io_in[7];
	assign _02615_ = _02614_ | _06310_;
	assign _02617_ = io_in[11] & ~_02615_;
	assign _02618_ = _06532_ | _03094_;
	assign _02619_ = _02618_ | _03759_;
	assign _02620_ = _02619_ | io_in[7];
	assign _02621_ = _02620_ | _01208_;
	assign _02622_ = _01985_ & ~_02621_;
	assign _02623_ = _01138_ | _02207_;
	assign _02624_ = _02623_ | _01208_;
	assign _02625_ = _02624_ | _06310_;
	assign _02626_ = _01985_ & ~_02625_;
	assign _02628_ = _07343_ | _02207_;
	assign _02629_ = _02628_ | _01208_;
	assign _02630_ = _02629_ | _02096_;
	assign _02631_ = _02630_ | _06310_;
	assign _02632_ = _01985_ & ~_02631_;
	assign _02633_ = _01203_ | io_in[8];
	assign _02634_ = io_in[10] & ~_02633_;
	assign _02635_ = _04458_ | _03094_;
	assign _02636_ = _02635_ | _02207_;
	assign _02637_ = io_in[11] & ~_02636_;
	assign _02639_ = _01710_ | io_in[7];
	assign _02640_ = _02639_ | _01208_;
	assign _02641_ = io_in[11] & ~_02640_;
	assign _02642_ = _00010_ | _03094_;
	assign _02643_ = _02642_ | io_in[6];
	assign _02644_ = _02643_ | _02207_;
	assign _02645_ = io_in[11] & ~_02644_;
	assign _02646_ = _01334_ | io_in[8];
	assign _02647_ = _02646_ | _02096_;
	assign _02648_ = io_in[11] & ~_02647_;
	assign _02651_ = _06609_ | io_in[6];
	assign _02652_ = _02651_ | _02207_;
	assign _02653_ = _02096_ & ~_02652_;
	assign _02654_ = _01438_ | io_in[6];
	assign _02655_ = _02654_ | _02207_;
	assign _02656_ = _02655_ | _01208_;
	assign _02657_ = _02656_ | _02096_;
	assign _02658_ = _01985_ & ~_02657_;
	assign _02659_ = _04990_ | _03759_;
	assign _02660_ = _02659_ | _06310_;
	assign _02662_ = io_in[11] & ~_02660_;
	assign _02663_ = _01483_ | io_in[5];
	assign _02664_ = _02663_ | _03759_;
	assign _02665_ = _02664_ | io_in[7];
	assign _02666_ = _02665_ | io_in[8];
	assign _02667_ = _02666_ | io_in[9];
	assign _02668_ = io_in[11] & ~_02667_;
	assign _02669_ = _07086_ | _02207_;
	assign _02670_ = _02669_ | io_in[9];
	assign _02671_ = _02670_ | io_in[10];
	assign _02673_ = _01985_ & ~_02671_;
	assign _02674_ = _01870_ | _03759_;
	assign _02675_ = _02674_ | io_in[7];
	assign _02676_ = _02675_ | io_in[8];
	assign _02677_ = _02676_ | io_in[9];
	assign _02678_ = _06310_ & ~_02677_;
	assign _02679_ = _01299_ | io_in[8];
	assign _02680_ = io_in[9] & ~_02679_;
	assign _02681_ = _00458_ | _01208_;
	assign _02682_ = _02681_ | _02096_;
	assign _02684_ = _02682_ | _06310_;
	assign _02685_ = _01985_ & ~_02684_;
	assign _02686_ = _01878_ | io_in[5];
	assign _02687_ = _02686_ | _03759_;
	assign _02688_ = _02687_ | _02207_;
	assign _02689_ = _02688_ | _02096_;
	assign _02690_ = _02689_ | _06310_;
	assign _02691_ = _01985_ & ~_02690_;
	assign _02692_ = _07383_ | io_in[6];
	assign _02693_ = _02692_ | _02207_;
	assign _02695_ = _02693_ | io_in[8];
	assign _02696_ = _02695_ | io_in[9];
	assign _02697_ = io_in[10] & ~_02696_;
	assign _02698_ = _01537_ | _03759_;
	assign _02699_ = _02698_ | _01208_;
	assign _02700_ = _02699_ | io_in[9];
	assign _02701_ = io_in[11] & ~_02700_;
	assign _02702_ = _01617_ | _01208_;
	assign _02703_ = _02096_ & ~_02702_;
	assign _02704_ = _07359_ | _02096_;
	assign _02706_ = _02704_ | io_in[10];
	assign _02707_ = io_in[11] & ~_02706_;
	assign _02708_ = _01786_ | io_in[7];
	assign _02709_ = _02708_ | io_in[9];
	assign _02710_ = _01985_ & ~_02709_;
	assign _02711_ = _04103_ | io_in[6];
	assign _02712_ = _02711_ | io_in[8];
	assign _02713_ = _02712_ | io_in[10];
	assign _02714_ = _01985_ & ~_02713_;
	assign _02715_ = _01547_ | io_in[7];
	assign _02717_ = _02715_ | _01208_;
	assign _02718_ = _02717_ | io_in[9];
	assign _02719_ = _06310_ & ~_02718_;
	assign _02720_ = _07392_ | _03759_;
	assign _02721_ = _02720_ | _02207_;
	assign _02722_ = _02721_ | io_in[8];
	assign _02723_ = _02722_ | _02096_;
	assign _02724_ = _06310_ & ~_02723_;
	assign _02725_ = _02549_ | _02207_;
	assign _02726_ = _02725_ | io_in[10];
	assign _02728_ = io_in[11] & ~_02726_;
	assign _02729_ = _01483_ | io_in[7];
	assign _02730_ = _02729_ | io_in[8];
	assign _02731_ = io_in[10] & ~_02730_;
	assign _02732_ = _01647_ | _02207_;
	assign _02733_ = _02096_ & ~_02732_;
	assign _02734_ = _01422_ | io_in[7];
	assign _02735_ = _02734_ | _01208_;
	assign _02736_ = io_in[11] & ~_02735_;
	assign _02737_ = _07255_ | io_in[8];
	assign _02739_ = _02737_ | _02096_;
	assign _02740_ = _02739_ | io_in[10];
	assign _02741_ = _01985_ & ~_02740_;
	assign _02742_ = _00439_ | io_in[7];
	assign _02743_ = _02742_ | io_in[8];
	assign _02744_ = _02743_ | io_in[10];
	assign _02745_ = _01985_ & ~_02744_;
	assign _02746_ = _06243_ | _01208_;
	assign _02747_ = _02746_ | io_in[9];
	assign _02748_ = _02747_ | io_in[10];
	assign _02750_ = _01985_ & ~_02748_;
	assign _02751_ = _07499_ | _07422_;
	assign _02752_ = _02751_ | _03759_;
	assign _02753_ = _02752_ | io_in[8];
	assign _02754_ = _02753_ | _02096_;
	assign _02755_ = io_in[11] & ~_02754_;
	assign _02756_ = _01013_ | _03759_;
	assign _02757_ = _02756_ | io_in[8];
	assign _02758_ = _02757_ | io_in[10];
	assign _02759_ = _01985_ & ~_02758_;
	assign _02762_ = _01138_ | io_in[8];
	assign _02763_ = _02762_ | io_in[9];
	assign _02764_ = io_in[10] & ~_02763_;
	assign _02765_ = _01434_ | _01208_;
	assign _02766_ = _02765_ | _02096_;
	assign _02767_ = _06310_ & ~_02766_;
	assign _02768_ = _07289_ | _03094_;
	assign _02769_ = _02207_ & ~_02768_;
	assign _02770_ = _02751_ | io_in[6];
	assign _02771_ = _02770_ | io_in[7];
	assign _02773_ = _02771_ | _02096_;
	assign _02774_ = _02773_ | _06310_;
	assign _02775_ = _01985_ & ~_02774_;
	assign _02776_ = _01289_ | _06310_;
	assign _02777_ = _01985_ & ~_02776_;
	assign _02778_ = _01031_ | io_in[4];
	assign _02779_ = _02778_ | io_in[5];
	assign _02780_ = _02779_ | _03759_;
	assign _02781_ = _02780_ | io_in[7];
	assign _02782_ = _02781_ | _01208_;
	assign _02784_ = _02782_ | _02096_;
	assign _02785_ = io_in[10] & ~_02784_;
	assign _02786_ = _01214_ | io_in[6];
	assign _02787_ = _02786_ | io_in[7];
	assign _02788_ = _02787_ | io_in[10];
	assign _02789_ = io_in[11] & ~_02788_;
	assign _02790_ = _01038_ | _02207_;
	assign _02791_ = _02790_ | _01208_;
	assign _02792_ = _06310_ & ~_02791_;
	assign _02793_ = _07410_ | _03094_;
	assign _02795_ = _02793_ | _03759_;
	assign _02796_ = _02795_ | _02096_;
	assign _02797_ = io_in[10] & ~_02796_;
	assign _02798_ = _06853_ | _03094_;
	assign _02799_ = _02798_ | _02207_;
	assign _02800_ = _02799_ | io_in[8];
	assign _02801_ = io_in[9] & ~_02800_;
	assign _02802_ = _01066_ | _02207_;
	assign _02803_ = _02802_ | io_in[8];
	assign _02804_ = _02803_ | io_in[9];
	assign _02806_ = _02804_ | _06310_;
	assign _02807_ = _01985_ & ~_02806_;
	assign _02808_ = _00274_ | io_in[6];
	assign _02809_ = _02808_ | _02207_;
	assign _02810_ = _02809_ | io_in[8];
	assign _02811_ = _02810_ | _02096_;
	assign _02812_ = io_in[11] & ~_02811_;
	assign _02813_ = _01982_ | io_in[6];
	assign _02814_ = _02813_ | _02207_;
	assign _02815_ = _02814_ | io_in[8];
	assign _02817_ = _02815_ | io_in[9];
	assign _02818_ = io_in[11] & ~_02817_;
	assign _02819_ = _06864_ | _03759_;
	assign _02820_ = _02819_ | io_in[8];
	assign _02821_ = _02820_ | _02096_;
	assign _02822_ = _06310_ & ~_02821_;
	assign _02823_ = _01025_ | io_in[7];
	assign _02824_ = _02823_ | io_in[8];
	assign _02825_ = _01985_ & ~_02824_;
	assign _02826_ = _02489_ | io_in[8];
	assign _02828_ = _02826_ | io_in[9];
	assign _02829_ = io_in[10] & ~_02828_;
	assign _02830_ = _01541_ | io_in[7];
	assign _02831_ = _02830_ | io_in[8];
	assign _02832_ = _02831_ | io_in[10];
	assign _02833_ = _01985_ & ~_02832_;
	assign _02834_ = _02437_ | io_in[7];
	assign _02835_ = _02834_ | _02096_;
	assign _02836_ = _06310_ & ~_02835_;
	assign _02837_ = _04978_ | io_in[8];
	assign _02839_ = _02837_ | io_in[9];
	assign _02840_ = io_in[10] & ~_02839_;
	assign _02841_ = _01029_ | io_in[7];
	assign _02842_ = _02841_ | _01208_;
	assign _02843_ = io_in[9] & ~_02842_;
	assign _02844_ = _02843_ & ~io_in[10];
	assign _02845_ = _01991_ | _02096_;
	assign _02846_ = _01985_ & ~_02845_;
	assign _02847_ = _01456_ | io_in[6];
	assign _02848_ = _02847_ | _01208_;
	assign _02850_ = _06310_ & ~_02848_;
	assign _02851_ = _01757_ | _02207_;
	assign _02852_ = _02851_ | _01208_;
	assign _02853_ = _02852_ | _06310_;
	assign _02854_ = _01985_ & ~_02853_;
	assign _02855_ = _03260_ | io_in[5];
	assign _02856_ = _02855_ | io_in[6];
	assign _02857_ = _02856_ | _02207_;
	assign _02858_ = _02857_ | _06310_;
	assign _02859_ = io_in[11] & ~_02858_;
	assign _02861_ = _01842_ | _02096_;
	assign _02862_ = io_in[10] & ~_02861_;
	assign _02863_ = _01112_ | io_in[8];
	assign _02864_ = _02863_ | io_in[9];
	assign _02865_ = io_in[11] & ~_02864_;
	assign _02866_ = _07367_ | _03094_;
	assign _02867_ = _02866_ | _02207_;
	assign _02868_ = _02867_ | _01208_;
	assign _02869_ = io_in[10] & ~_02868_;
	assign _02870_ = ~(io_in[5] & io_in[0]);
	assign _02873_ = _02870_ | _03759_;
	assign _02874_ = _02873_ | _02096_;
	assign _02875_ = _02874_ | io_in[10];
	assign _02876_ = io_in[11] & ~_02875_;
	assign _02877_ = _01931_ | io_in[9];
	assign _02878_ = _02877_ | io_in[10];
	assign _02879_ = _01985_ & ~_02878_;
	assign _02880_ = _02751_ | _02207_;
	assign _02881_ = _02880_ | io_in[9];
	assign _02882_ = _02881_ | io_in[10];
	assign _02884_ = _01985_ & ~_02882_;
	assign _02885_ = _01154_ | _02096_;
	assign _02886_ = io_in[10] & ~_02885_;
	assign _02887_ = ~(_03049_ & _06310_);
	assign _02888_ = _01985_ & ~_02887_;
	assign _02889_ = _02073_ | _01208_;
	assign _02890_ = _02096_ & ~_02889_;
	assign _02891_ = _00998_ | _02207_;
	assign _02892_ = _02891_ | _06310_;
	assign _02893_ = io_in[11] & ~_02892_;
	assign _02895_ = _00484_ | _02207_;
	assign _02896_ = _02895_ | _02096_;
	assign _02897_ = _02896_ | io_in[10];
	assign _02898_ = io_in[11] & ~_02897_;
	assign _02899_ = _04302_ | io_in[5];
	assign _02900_ = _02899_ | io_in[6];
	assign _02901_ = _02900_ | _02207_;
	assign _02902_ = _02901_ | _01208_;
	assign _02903_ = io_in[11] & ~_02902_;
	assign _02904_ = _01202_ | _02207_;
	assign _02906_ = _02904_ | _01208_;
	assign _02907_ = _02906_ | _02096_;
	assign _02908_ = _06310_ & ~_02907_;
	assign _02909_ = _07376_ | io_in[7];
	assign _02910_ = _02909_ | io_in[8];
	assign _02911_ = io_in[10] & ~_02910_;
	assign _02912_ = _02971_ | _03759_;
	assign _02913_ = _02912_ | _02207_;
	assign _02914_ = _02913_ | _01208_;
	assign _02915_ = _02914_ | io_in[9];
	assign _02917_ = io_in[10] & ~_02915_;
	assign _02918_ = _01553_ | _02207_;
	assign _02919_ = _02918_ | io_in[8];
	assign _02920_ = _02919_ | io_in[9];
	assign _02921_ = io_in[10] & ~_02920_;
	assign _02922_ = _00985_ | _03759_;
	assign _02923_ = _02922_ | _01208_;
	assign _02924_ = _02923_ | io_in[9];
	assign _02925_ = io_in[10] & ~_02924_;
	assign _02926_ = _02756_ | io_in[7];
	assign _02928_ = _02926_ | _01208_;
	assign _02929_ = _02096_ & ~_02928_;
	assign _02930_ = _00246_ | io_in[5];
	assign _02931_ = _02930_ | _03759_;
	assign _02932_ = _02931_ | io_in[7];
	assign _02933_ = _02932_ | _06310_;
	assign _02934_ = io_in[11] & ~_02933_;
	assign _02935_ = _02982_ | _03759_;
	assign _02936_ = _02935_ | io_in[7];
	assign _02937_ = _02936_ | io_in[8];
	assign _02939_ = _02937_ | io_in[9];
	assign _02940_ = io_in[11] & ~_02939_;
	assign _02941_ = _01057_ | _03759_;
	assign _02942_ = _02941_ | _02207_;
	assign _02943_ = _02942_ | _01208_;
	assign _02944_ = _02943_ | _02096_;
	assign _02945_ = _02944_ | _06310_;
	assign _02946_ = _01985_ & ~_02945_;
	assign _02947_ = _01960_ | io_in[8];
	assign _02948_ = _02947_ | _02096_;
	assign _02950_ = _01985_ & ~_02948_;
	assign _02951_ = _01213_ | io_in[6];
	assign _02952_ = _02951_ | _02207_;
	assign _02953_ = _02952_ | _01208_;
	assign _02954_ = io_in[10] & ~_02953_;
	assign _02955_ = _06754_ | _03094_;
	assign _02956_ = _03759_ & ~_02955_;
	assign _02957_ = _04302_ | _01208_;
	assign _02958_ = _02957_ | io_in[9];
	assign _02959_ = _06310_ & ~_02958_;
	assign _02961_ = _03304_ | _03759_;
	assign _02962_ = _02961_ | io_in[7];
	assign _02963_ = _02962_ | io_in[8];
	assign _02964_ = _02963_ | io_in[9];
	assign _02965_ = io_in[10] & ~_02964_;
	assign _02966_ = _01334_ | _03759_;
	assign _02967_ = _02966_ | io_in[8];
	assign _02968_ = _02967_ | _02096_;
	assign _02969_ = io_in[10] & ~_02968_;
	assign _02970_ = _01757_ | io_in[6];
	assign _02972_ = _02970_ | io_in[7];
	assign _02973_ = _02972_ | _02096_;
	assign _02974_ = io_in[11] & ~_02973_;
	assign _02975_ = _04047_ | io_in[6];
	assign _02976_ = _02975_ | _02207_;
	assign _02977_ = _02976_ | _01208_;
	assign _02978_ = _02977_ | io_in[9];
	assign _02979_ = io_in[10] & ~_02978_;
	assign _02980_ = _03304_ | io_in[5];
	assign _02981_ = _02980_ | io_in[6];
	assign _02984_ = _02981_ | _02207_;
	assign _02985_ = _02984_ | io_in[8];
	assign _02986_ = _02985_ | io_in[9];
	assign _02987_ = io_in[10] & ~_02986_;
	assign _02988_ = _00414_ | io_in[7];
	assign _02989_ = _02988_ | io_in[8];
	assign _02990_ = _02989_ | _02096_;
	assign _02991_ = io_in[10] & ~_02990_;
	assign _02992_ = _07419_ | io_in[6];
	assign _02993_ = _02992_ | io_in[7];
	assign _02995_ = _02993_ | _01208_;
	assign _02996_ = _02995_ | io_in[9];
	assign _02997_ = io_in[10] & ~_02996_;
	assign _02998_ = _06754_ | io_in[6];
	assign _02999_ = _02998_ | io_in[7];
	assign _03000_ = _02999_ | io_in[8];
	assign _03001_ = _02096_ & ~_03000_;
	assign _03002_ = _07358_ | _03759_;
	assign _03003_ = _03002_ | io_in[7];
	assign _03004_ = _03003_ | _01208_;
	assign _03006_ = _03004_ | io_in[9];
	assign _03007_ = _01985_ & ~_03006_;
	assign _03008_ = _00010_ | io_in[6];
	assign _03009_ = _03008_ | _02207_;
	assign _03010_ = _03009_ | io_in[9];
	assign _03011_ = _01985_ & ~_03010_;
	assign _03012_ = ~(_00517_ & _06310_);
	assign _03013_ = _01985_ & ~_03012_;
	assign _03014_ = _01930_ | io_in[7];
	assign _03015_ = _03014_ | io_in[8];
	assign _03017_ = io_in[9] & ~_03015_;
	assign _03018_ = _02778_ | _03759_;
	assign _03019_ = _03018_ | _02207_;
	assign _03020_ = _03019_ | io_in[8];
	assign _03021_ = _03020_ | io_in[9];
	assign _03022_ = io_in[10] & ~_03021_;
	assign _03023_ = _01617_ | _02207_;
	assign _03024_ = io_in[10] & ~_03023_;
	assign _03025_ = _01814_ | _01208_;
	assign _03026_ = io_in[9] & ~_03025_;
	assign _03028_ = _01133_ | _02207_;
	assign _03029_ = _03028_ | _01208_;
	assign _03030_ = _03029_ | io_in[9];
	assign _03031_ = io_in[11] & ~_03030_;
	assign _03032_ = _02096_ & ~_02574_;
	assign _03033_ = _03149_ | _03094_;
	assign _03034_ = _03033_ | _02207_;
	assign _03035_ = _03034_ | io_in[9];
	assign _03036_ = _01985_ & ~_03035_;
	assign _03037_ = _01327_ | io_in[8];
	assign _03039_ = io_in[10] & ~_03037_;
	assign _03040_ = _01184_ | io_in[8];
	assign _03041_ = _03040_ | _02096_;
	assign _03042_ = io_in[10] & ~_03041_;
	assign _03043_ = _01184_ | _02207_;
	assign _03044_ = _03043_ | _01208_;
	assign _03045_ = _03044_ | _02096_;
	assign _03046_ = _01985_ & ~_03045_;
	assign _03047_ = _01089_ | io_in[8];
	assign _03048_ = io_in[9] & ~_03047_;
	assign _03050_ = _05989_ | io_in[7];
	assign _03051_ = _03050_ | _02096_;
	assign _03052_ = _06310_ & ~_03051_;
	assign _03053_ = _00246_ | _02207_;
	assign _03054_ = _03053_ | _01208_;
	assign _03055_ = _03054_ | _02096_;
	assign _03056_ = _06310_ & ~_03055_;
	assign _03057_ = _00986_ | io_in[5];
	assign _03058_ = _03057_ | io_in[6];
	assign _03059_ = _03058_ | _02207_;
	assign _03061_ = _03059_ | _02096_;
	assign _03062_ = io_in[11] & ~_03061_;
	assign _03063_ = _02313_ | io_in[9];
	assign _03064_ = io_in[11] & ~_03063_;
	assign _03065_ = _07412_ | io_in[7];
	assign _03066_ = _03065_ | _01208_;
	assign _03067_ = _03066_ | _02096_;
	assign _03068_ = _03067_ | _06310_;
	assign _03069_ = _01985_ & ~_03068_;
	assign _03070_ = _02770_ | _02207_;
	assign _03072_ = _03070_ | _01208_;
	assign _03073_ = _03072_ | _02096_;
	assign _03074_ = _06310_ & ~_03073_;
	assign _03075_ = _05989_ | io_in[5];
	assign _03076_ = _03075_ | io_in[6];
	assign _03077_ = _03076_ | _02096_;
	assign _03078_ = io_in[11] & ~_03077_;
	assign _03079_ = _00768_ | io_in[6];
	assign _03080_ = _03079_ | _02207_;
	assign _03081_ = _03080_ | io_in[8];
	assign _03083_ = io_in[9] & ~_03081_;
	assign _03084_ = _00720_ | io_in[6];
	assign _03085_ = _03084_ | io_in[7];
	assign _03086_ = _03085_ | io_in[8];
	assign _03087_ = _02096_ & ~_03086_;
	assign _03088_ = _02378_ | io_in[9];
	assign _03089_ = io_in[10] & ~_03088_;
	assign _03090_ = _00598_ | io_in[5];
	assign _03091_ = _03090_ | io_in[7];
	assign _03092_ = _03091_ | _01208_;
	assign _03095_ = _03092_ | _02096_;
	assign _03096_ = _03095_ | _06310_;
	assign _03097_ = _01985_ & ~_03096_;
	assign _03098_ = _01038_ | _01208_;
	assign _03099_ = _03098_ | io_in[9];
	assign _03100_ = io_in[11] & ~_03099_;
	assign _03101_ = _00531_ | _03759_;
	assign _03102_ = _03101_ | io_in[7];
	assign _03103_ = _03102_ | _06310_;
	assign _03104_ = io_in[11] & ~_03103_;
	assign _03106_ = _01596_ | _03094_;
	assign _03107_ = _03106_ | _02207_;
	assign _03108_ = _03107_ | io_in[8];
	assign _03109_ = _06310_ & ~_03108_;
	assign _03110_ = _01236_ | _02207_;
	assign _03111_ = _03110_ | io_in[9];
	assign _03112_ = _03111_ | io_in[10];
	assign _03113_ = io_in[11] & ~_03112_;
	assign _03114_ = _04990_ | _02207_;
	assign _03115_ = _03114_ | _06310_;
	assign _03117_ = io_in[11] & ~_03115_;
	assign _03118_ = _07335_ | io_in[6];
	assign _03119_ = _03118_ | io_in[7];
	assign _03120_ = _03119_ | _01208_;
	assign _03121_ = _03120_ | _02096_;
	assign _03122_ = _06310_ & ~_03121_;
	assign _03123_ = _03371_ | _01208_;
	assign _03124_ = _03123_ | io_in[9];
	assign _03125_ = io_in[10] & ~_03124_;
	assign _03126_ = _02870_ | _02207_;
	assign _03128_ = _03126_ | _02096_;
	assign _03129_ = _03128_ | io_in[10];
	assign _03130_ = io_in[11] & ~_03129_;
	assign _03131_ = _01260_ | _01208_;
	assign _03132_ = _03131_ | io_in[10];
	assign _03133_ = io_in[11] & ~_03132_;
	assign _03134_ = _00766_ | _03094_;
	assign _03135_ = io_in[6] & ~_03134_;
	assign _03136_ = _01809_ | io_in[8];
	assign _03137_ = _03136_ | io_in[9];
	assign _03139_ = io_in[11] & ~_03137_;
	assign _03140_ = _01213_ | _03759_;
	assign _03141_ = _03140_ | io_in[7];
	assign _03142_ = _03141_ | _01208_;
	assign _03143_ = io_in[10] & ~_03142_;
	assign _03144_ = _02619_ | _01208_;
	assign _03145_ = _03144_ | _02096_;
	assign _03146_ = _06310_ & ~_03145_;
	assign _03147_ = _01505_ | _02096_;
	assign _03148_ = _03147_ | io_in[10];
	assign _03150_ = io_in[11] & ~_03148_;
	assign _03151_ = _04901_ | _02207_;
	assign _03152_ = _03151_ | io_in[10];
	assign _03153_ = io_in[11] & ~_03152_;
	assign _03154_ = _00955_ | io_in[10];
	assign _03155_ = _01985_ & ~_03154_;
	assign _03156_ = _01001_ | io_in[7];
	assign _03157_ = _03156_ | _01208_;
	assign _03158_ = _03157_ | io_in[9];
	assign _03159_ = io_in[10] & ~_03158_;
	assign _03161_ = _00679_ | io_in[6];
	assign _03162_ = _03161_ | io_in[7];
	assign _03163_ = _03162_ | _02096_;
	assign _03164_ = _06310_ & ~_03163_;
	assign _03165_ = _07153_ | io_in[7];
	assign _03166_ = _03165_ | io_in[8];
	assign _03167_ = _03166_ | io_in[9];
	assign _03168_ = io_in[11] & ~_03167_;
	assign _03169_ = _07250_ | _02207_;
	assign _03170_ = _03169_ | io_in[8];
	assign _03172_ = _03170_ | _02096_;
	assign _03173_ = io_in[10] & ~_03172_;
	assign _03174_ = _01607_ | io_in[6];
	assign _03175_ = _03174_ | io_in[7];
	assign _03176_ = _03175_ | io_in[8];
	assign _03177_ = _03176_ | _02096_;
	assign _03178_ = io_in[11] & ~_03177_;
	assign _03179_ = _03747_ | io_in[7];
	assign _03180_ = _03179_ | _02096_;
	assign _03181_ = _06310_ & ~_03180_;
	assign _03183_ = _07362_ | _03759_;
	assign _03184_ = _03183_ | _01208_;
	assign _03185_ = _03184_ | io_in[9];
	assign _03186_ = io_in[10] & ~_03185_;
	assign _03187_ = _02018_ | io_in[5];
	assign _03188_ = _03187_ | io_in[6];
	assign _03189_ = _03188_ | _02207_;
	assign _03190_ = _03189_ | io_in[8];
	assign _03191_ = _03190_ | _02096_;
	assign _03192_ = _03191_ | io_in[10];
	assign _03194_ = io_in[11] & ~_03192_;
	assign _03195_ = _01758_ | _06310_;
	assign _03196_ = io_in[11] & ~_03195_;
	assign _03197_ = _01391_ | io_in[6];
	assign _03198_ = _03197_ | _02207_;
	assign _03199_ = _03198_ | io_in[9];
	assign _03200_ = io_in[10] & ~_03199_;
	assign _03201_ = _06531_ | io_in[8];
	assign _03202_ = _03201_ | io_in[9];
	assign _03203_ = io_in[10] & ~_03202_;
	assign _03206_ = _01983_ | _02207_;
	assign _03207_ = _03206_ | io_in[8];
	assign _03208_ = _03207_ | _02096_;
	assign _03209_ = io_in[10] & ~_03208_;
	assign _03210_ = _03054_ | io_in[9];
	assign _03211_ = io_in[10] & ~_03210_;
	assign _03212_ = _01322_ | io_in[7];
	assign _03213_ = _03212_ | _01208_;
	assign _03214_ = _03213_ | _02096_;
	assign _03215_ = _06310_ & ~_03214_;
	assign _03217_ = _07392_ | io_in[6];
	assign _03218_ = _03217_ | io_in[7];
	assign _03219_ = _03218_ | _06310_;
	assign _03220_ = io_in[11] & ~_03219_;
	assign _03221_ = _01636_ | _01208_;
	assign _03222_ = _03221_ | io_in[9];
	assign _03223_ = io_in[10] & ~_03222_;
	assign _03224_ = _07302_ | io_in[5];
	assign _03225_ = _03224_ | _03759_;
	assign _03226_ = _03225_ | io_in[7];
	assign _03228_ = _03226_ | _06310_;
	assign _03229_ = io_in[11] & ~_03228_;
	assign _03230_ = _02654_ | io_in[7];
	assign _03231_ = _03230_ | _01208_;
	assign _03232_ = _03231_ | io_in[10];
	assign _03233_ = io_in[11] & ~_03232_;
	assign _03234_ = _01251_ | io_in[9];
	assign _03235_ = _03234_ | io_in[10];
	assign _03236_ = _01985_ & ~_03235_;
	assign _03237_ = _04313_ | _02207_;
	assign _03239_ = _03237_ | io_in[10];
	assign _03240_ = io_in[11] & ~_03239_;
	assign _03241_ = _01195_ | _01208_;
	assign _03242_ = _03241_ | io_in[10];
	assign _03243_ = _01985_ & ~_03242_;
	assign _03244_ = _02982_ | io_in[6];
	assign _03245_ = _03244_ | io_in[7];
	assign _03246_ = _03245_ | io_in[8];
	assign _03247_ = _03246_ | _02096_;
	assign _03248_ = io_in[11] & ~_03247_;
	assign _03250_ = _02798_ | _03759_;
	assign _03251_ = _03250_ | io_in[8];
	assign _03252_ = io_in[10] & ~_03251_;
	assign _03253_ = _01850_ | io_in[7];
	assign _03254_ = _03253_ | io_in[8];
	assign _03255_ = io_in[9] & ~_03254_;
	assign _03256_ = _03027_ | _01208_;
	assign _03257_ = _03256_ | io_in[9];
	assign _03258_ = _03257_ | io_in[10];
	assign _03259_ = _01985_ & ~_03258_;
	assign _03261_ = _03259_ | _03255_;
	assign _03262_ = _03261_ | _03252_;
	assign _03263_ = _03262_ | _03248_;
	assign _03264_ = _03263_ | _03243_;
	assign _03265_ = _03264_ | _03240_;
	assign _03266_ = _03265_ | _03236_;
	assign _03267_ = _03266_ | _03233_;
	assign _03268_ = _03267_ | _03229_;
	assign _03269_ = _03268_ | _03223_;
	assign _03270_ = _03269_ | _03220_;
	assign _03272_ = _03270_ | _03215_;
	assign _03273_ = _03272_ | _03211_;
	assign _03274_ = _03273_ | _03209_;
	assign _03275_ = _03274_ | _03203_;
	assign _03276_ = _03275_ | _03200_;
	assign _03277_ = _03276_ | _03196_;
	assign _03278_ = _03277_ | _03194_;
	assign _03279_ = _03278_ | _03186_;
	assign _03280_ = _03279_ | _03181_;
	assign _03281_ = _03280_ | _03178_;
	assign _03283_ = _03281_ | _03173_;
	assign _03284_ = _03283_ | _03168_;
	assign _03285_ = _03284_ | _03164_;
	assign _03286_ = _03285_ | _03159_;
	assign _03287_ = _03286_ | _03155_;
	assign _03288_ = _03287_ | _03153_;
	assign _03289_ = _03288_ | _03150_;
	assign _03290_ = _03289_ | _03146_;
	assign _03291_ = _03290_ | _03143_;
	assign _03292_ = _03291_ | _03139_;
	assign _03294_ = _03292_ | _03135_;
	assign _03295_ = _03294_ | _03133_;
	assign _03296_ = _03295_ | _03130_;
	assign _03297_ = _03296_ | _03125_;
	assign _03298_ = _03297_ | _03122_;
	assign _03299_ = _03298_ | _03117_;
	assign _03300_ = _03299_ | _03113_;
	assign _03301_ = _03300_ | _03109_;
	assign _03302_ = _03301_ | _03104_;
	assign _03303_ = _03302_ | _03100_;
	assign _03305_ = _03303_ | _03097_;
	assign _03306_ = _03305_ | _03089_;
	assign _03307_ = _03306_ | _03087_;
	assign _03308_ = _03307_ | _03083_;
	assign _03309_ = _03308_ | _03078_;
	assign _03310_ = _03309_ | _03074_;
	assign _03311_ = _03310_ | _03069_;
	assign _03312_ = _03311_ | _03064_;
	assign _03313_ = _03312_ | _03062_;
	assign _03314_ = _03313_ | _03056_;
	assign _03317_ = _03314_ | _03052_;
	assign _03318_ = _03317_ | _03048_;
	assign _03319_ = _03318_ | _03046_;
	assign _03320_ = _03319_ | _03042_;
	assign _03321_ = _03320_ | _03039_;
	assign _03322_ = _03321_ | _03036_;
	assign _03323_ = _03322_ | _03032_;
	assign _03324_ = _03323_ | _03031_;
	assign _03325_ = _03324_ | _03026_;
	assign _03326_ = _03325_ | _03024_;
	assign _03328_ = _03326_ | _03022_;
	assign _03329_ = _03328_ | _03017_;
	assign _03330_ = _03329_ | _03013_;
	assign _03331_ = _03330_ | _03011_;
	assign _03332_ = _03331_ | _03007_;
	assign _03333_ = _03332_ | _03001_;
	assign _03334_ = _03333_ | _02997_;
	assign _03335_ = _03334_ | _02991_;
	assign _03336_ = _03335_ | _02987_;
	assign _03337_ = _03336_ | _02979_;
	assign _03339_ = _03337_ | _02974_;
	assign _03340_ = _03339_ | _02969_;
	assign _03341_ = _03340_ | _02965_;
	assign _03342_ = _03341_ | _02959_;
	assign _03343_ = _03342_ | _02956_;
	assign _03344_ = _03343_ | _02954_;
	assign _03345_ = _03344_ | _02950_;
	assign _03346_ = _03345_ | _02946_;
	assign _03347_ = _03346_ | _02940_;
	assign _03348_ = _03347_ | _02934_;
	assign _03350_ = _03348_ | _02929_;
	assign _03351_ = _03350_ | _02925_;
	assign _03352_ = _03351_ | _02921_;
	assign _03353_ = _03352_ | _02917_;
	assign _03354_ = _03353_ | _02911_;
	assign _03355_ = _03354_ | _02908_;
	assign _03356_ = _03355_ | _02903_;
	assign _03357_ = _03356_ | _02898_;
	assign _03358_ = _03357_ | _02893_;
	assign _03359_ = _03358_ | _02890_;
	assign _03361_ = _03359_ | _02888_;
	assign _03362_ = _03361_ | _02886_;
	assign _03363_ = _03362_ | _02884_;
	assign _03364_ = _03363_ | _02879_;
	assign _03365_ = _03364_ | _02876_;
	assign _03366_ = _03365_ | _02869_;
	assign _03367_ = _03366_ | _02865_;
	assign _03368_ = _03367_ | _02862_;
	assign _03369_ = _03368_ | _02859_;
	assign _03370_ = _03369_ | _02854_;
	assign _03372_ = _03370_ | _02850_;
	assign _03373_ = _03372_ | _02846_;
	assign _03374_ = _03373_ | _02844_;
	assign _03375_ = _03374_ | _02840_;
	assign _03376_ = _03375_ | _02836_;
	assign _03377_ = _03376_ | _02833_;
	assign _03378_ = _03377_ | _02829_;
	assign _03379_ = _03378_ | _02825_;
	assign _03380_ = _03379_ | _02822_;
	assign _03381_ = _03380_ | _02818_;
	assign _03383_ = _03381_ | _02812_;
	assign _03384_ = _03383_ | _02807_;
	assign _03385_ = _03384_ | _02801_;
	assign _03386_ = _03385_ | _02797_;
	assign _03387_ = _03386_ | _02792_;
	assign _03388_ = _03387_ | _02789_;
	assign _03389_ = _03388_ | _02785_;
	assign _03390_ = _03389_ | _02777_;
	assign _03391_ = _03390_ | _02775_;
	assign _03392_ = _03391_ | _02769_;
	assign _03394_ = _03392_ | _02767_;
	assign _03395_ = _03394_ | _02764_;
	assign _03396_ = _03395_ | _02759_;
	assign _03397_ = _03396_ | _02755_;
	assign _03398_ = _03397_ | _02750_;
	assign _03399_ = _03398_ | _02745_;
	assign _03400_ = _03399_ | _02741_;
	assign _03401_ = _03400_ | _02736_;
	assign _03402_ = _03401_ | _02733_;
	assign _03403_ = _03402_ | _02731_;
	assign _03405_ = _03403_ | _02728_;
	assign _03406_ = _03405_ | _02724_;
	assign _03407_ = _03406_ | _02719_;
	assign _03408_ = _03407_ | _02714_;
	assign _03409_ = _03408_ | _02710_;
	assign _03410_ = _03409_ | _02707_;
	assign _03411_ = _03410_ | _02703_;
	assign _03412_ = _03411_ | _02701_;
	assign _03413_ = _03412_ | _02697_;
	assign _03414_ = _03413_ | _02691_;
	assign _03416_ = _03414_ | _02685_;
	assign _03417_ = _03416_ | _02680_;
	assign _03418_ = _03417_ | _02678_;
	assign _03419_ = _03418_ | _02673_;
	assign _03420_ = _03419_ | _02668_;
	assign _03421_ = _03420_ | _02662_;
	assign _03422_ = _03421_ | _02658_;
	assign _03423_ = _03422_ | _02653_;
	assign _03424_ = _03423_ | _02648_;
	assign _03425_ = _03424_ | _02645_;
	assign _03428_ = _03425_ | _02641_;
	assign _03429_ = _03428_ | _02637_;
	assign _03430_ = _03429_ | _02634_;
	assign _03431_ = _03430_ | _02632_;
	assign _03432_ = _03431_ | _02626_;
	assign _03433_ = _03432_ | _02622_;
	assign _03434_ = _03433_ | _02617_;
	assign _03435_ = _03434_ | _02613_;
	assign _03436_ = _03435_ | _02610_;
	assign _03437_ = _03436_ | _02606_;
	assign _03439_ = _03437_ | _02601_;
	assign _03440_ = _03439_ | _02599_;
	assign _03441_ = _03440_ | _02596_;
	assign _03442_ = _03441_ | _02591_;
	assign _03443_ = _03442_ | _02588_;
	assign _03444_ = _03443_ | _02584_;
	assign _03445_ = _03444_ | _02580_;
	assign _03446_ = _03445_ | _02575_;
	assign _03447_ = _03446_ | _02570_;
	assign _03448_ = _03447_ | _02566_;
	assign _03450_ = _03448_ | _02562_;
	assign _03451_ = _03450_ | _02558_;
	assign _03452_ = _03451_ | _02554_;
	assign _03453_ = _03452_ | _02548_;
	assign _03454_ = _03453_ | _02542_;
	assign _03455_ = _03454_ | _02541_;
	assign _03456_ = _03455_ | _02534_;
	assign _03457_ = _03456_ | _02528_;
	assign _03458_ = _03457_ | _02523_;
	assign _03459_ = _03458_ | _02518_;
	assign _03461_ = _03459_ | _02514_;
	assign _03462_ = _03461_ | _02510_;
	assign _03463_ = _03462_ | _02508_;
	assign _03464_ = _03463_ | _02504_;
	assign _03465_ = _03464_ | _02500_;
	assign _03466_ = _03465_ | _02496_;
	assign _03467_ = _03466_ | _02492_;
	assign _03468_ = _03467_ | _02487_;
	assign _03469_ = _03468_ | _02482_;
	assign _03470_ = _03469_ | _02478_;
	assign _03472_ = _03470_ | _02476_;
	assign _03473_ = _03472_ | _02470_;
	assign _03474_ = _03473_ | _02466_;
	assign _03475_ = _03474_ | _02462_;
	assign _03476_ = _03475_ | _02457_;
	assign _03477_ = _03476_ | _02453_;
	assign _03478_ = _03477_ | _02448_;
	assign _03479_ = _03478_ | _02445_;
	assign _03480_ = _03479_ | _02441_;
	assign _03481_ = _03480_ | _02436_;
	assign _03483_ = _03481_ | _02433_;
	assign _03484_ = _03483_ | _02430_;
	assign _03485_ = _03484_ | _02424_;
	assign _03486_ = _03485_ | _02422_;
	assign _03487_ = _03486_ | _02420_;
	assign _03488_ = _03487_ | _02415_;
	assign _03489_ = _03488_ | _02411_;
	assign _03490_ = _03489_ | _02406_;
	assign _03491_ = _03490_ | _02400_;
	assign _03492_ = _03491_ | _02396_;
	assign _03494_ = _03492_ | _02392_;
	assign _03495_ = _03494_ | _02389_;
	assign _03496_ = _03495_ | _02385_;
	assign _03497_ = _03496_ | _02380_;
	assign _03498_ = _03497_ | _02377_;
	assign _03499_ = _03498_ | _02376_;
	assign _03500_ = _03499_ | _02371_;
	assign _03501_ = _03500_ | _02368_;
	assign _03502_ = _03501_ | _02364_;
	assign _03503_ = _03502_ | _02358_;
	assign _03505_ = _03503_ | _02354_;
	assign _03506_ = _03505_ | _02348_;
	assign _03507_ = _03506_ | _02343_;
	assign _03508_ = _03507_ | _02338_;
	assign _03509_ = _03508_ | _02337_;
	assign _03510_ = _03509_ | _02334_;
	assign _03511_ = _03510_ | _02332_;
	assign _03512_ = _03511_ | _02327_;
	assign _03513_ = _03512_ | _02322_;
	assign _03514_ = _03513_ | _02318_;
	assign _03516_ = _03514_ | _02311_;
	assign _03517_ = _03516_ | _02307_;
	assign _03518_ = _03517_ | _02303_;
	assign _03519_ = _03518_ | _02300_;
	assign _03520_ = _03519_ | _02298_;
	assign _03521_ = _03520_ | _02295_;
	assign _03522_ = _03521_ | _02290_;
	assign _03523_ = _03522_ | _02284_;
	assign _03524_ = _03523_ | _02281_;
	assign _03525_ = _03524_ | _02279_;
	assign _03527_ = _03525_ | _02278_;
	assign _03528_ = _03527_ | _02274_;
	assign _03529_ = _03528_ | _02269_;
	assign \mchip.val [3] = _03529_ | _02266_;
	assign _03530_ = _07368_ | _03094_;
	assign _03531_ = _03530_ | io_in[6];
	assign _03532_ = _02207_ & ~_03531_;
	assign _03533_ = _06509_ | io_in[5];
	assign _03534_ = _03533_ | _03759_;
	assign _03535_ = _03534_ | _02207_;
	assign _03538_ = _03535_ | _06310_;
	assign _03539_ = io_in[11] & ~_03538_;
	assign _03540_ = _07419_ | _02207_;
	assign _03541_ = _03540_ | io_in[9];
	assign _03542_ = _03541_ | io_in[10];
	assign _03543_ = _01985_ & ~_03542_;
	assign _03544_ = _01272_ | _01208_;
	assign _03545_ = _03544_ | io_in[9];
	assign _03546_ = _06310_ & ~_03545_;
	assign _03547_ = io_in[11] & ~_01882_;
	assign _03549_ = _00398_ | _03759_;
	assign _03550_ = _03549_ | io_in[7];
	assign _03551_ = _03550_ | _01208_;
	assign _03552_ = _03551_ | _02096_;
	assign _03553_ = _06310_ & ~_03552_;
	assign _03554_ = _02543_ | io_in[7];
	assign _03555_ = _03554_ | _01208_;
	assign _03556_ = _03555_ | io_in[9];
	assign _03557_ = io_in[10] & ~_03556_;
	assign _03558_ = _00679_ | _03759_;
	assign _03560_ = _03558_ | io_in[7];
	assign _03561_ = io_in[10] & ~_03560_;
	assign _03562_ = _07510_ | _03094_;
	assign _03563_ = _03562_ | io_in[9];
	assign _03564_ = io_in[11] & ~_03563_;
	assign _03565_ = _02350_ | _02207_;
	assign _03566_ = _03565_ | _01208_;
	assign _03567_ = _06310_ & ~_03566_;
	assign _03568_ = _03204_ | io_in[6];
	assign _03569_ = _03568_ | _02207_;
	assign _03571_ = _03569_ | _01208_;
	assign _03572_ = _03571_ | io_in[9];
	assign _03573_ = io_in[10] & ~_03572_;
	assign _03574_ = _01101_ | _02207_;
	assign _03575_ = _03574_ | io_in[8];
	assign _03576_ = io_in[9] & ~_03575_;
	assign _03577_ = _02351_ | _06310_;
	assign _03578_ = io_in[11] & ~_03577_;
	assign _03579_ = _01507_ | _02207_;
	assign _03580_ = _03579_ | _02096_;
	assign _03582_ = _06310_ & ~_03580_;
	assign _03583_ = _00972_ | io_in[6];
	assign _03584_ = _03583_ | _02207_;
	assign _03585_ = _03584_ | _01208_;
	assign _03586_ = io_in[10] & ~_03585_;
	assign _03587_ = _01272_ | io_in[7];
	assign _03588_ = _03587_ | _01208_;
	assign _03589_ = io_in[11] & ~_03588_;
	assign _03590_ = _04047_ | _03094_;
	assign _03591_ = _03590_ | _02207_;
	assign _03593_ = _03591_ | io_in[8];
	assign _03594_ = io_in[10] & ~_03593_;
	assign _03595_ = _01296_ | _03759_;
	assign _03596_ = _03595_ | io_in[7];
	assign _03597_ = _03596_ | _01208_;
	assign _03598_ = _03597_ | io_in[9];
	assign _03599_ = io_in[10] & ~_03598_;
	assign _03600_ = _00502_ | _02207_;
	assign _03601_ = _03600_ | io_in[8];
	assign _03602_ = _03601_ | io_in[9];
	assign _03604_ = io_in[11] & ~_03602_;
	assign _03605_ = _01080_ | io_in[8];
	assign _03606_ = _03605_ | io_in[9];
	assign _03607_ = _01985_ & ~_03606_;
	assign _03608_ = _00679_ | io_in[7];
	assign _03609_ = _03608_ | io_in[8];
	assign _03610_ = io_in[9] & ~_03609_;
	assign _03611_ = _00328_ | _03759_;
	assign _03612_ = _03611_ | _02207_;
	assign _03613_ = _03612_ | _01208_;
	assign _03615_ = _06310_ & ~_03613_;
	assign _03616_ = _02350_ | io_in[6];
	assign _03617_ = _03616_ | io_in[8];
	assign _03618_ = _02096_ & ~_03617_;
	assign _03619_ = _02922_ | _02207_;
	assign _03620_ = _03619_ | io_in[8];
	assign _03621_ = _02096_ & ~_03620_;
	assign _03622_ = _00173_ | _01208_;
	assign _03623_ = _03622_ | io_in[9];
	assign _03624_ = _03623_ | io_in[10];
	assign _03626_ = _01985_ & ~_03624_;
	assign _03627_ = _07419_ | _03759_;
	assign _03628_ = _03627_ | _01208_;
	assign _03629_ = _03628_ | _02096_;
	assign _03630_ = io_in[10] & ~_03629_;
	assign _03631_ = _00135_ | io_in[8];
	assign _03632_ = _02096_ & ~_03631_;
	assign _03633_ = _01406_ | io_in[8];
	assign _03634_ = _03633_ | _02096_;
	assign _03635_ = _06310_ & ~_03634_;
	assign _03637_ = _02539_ | _01208_;
	assign _03638_ = _03637_ | io_in[9];
	assign _03639_ = _03638_ | io_in[10];
	assign _03640_ = _01985_ & ~_03639_;
	assign _03641_ = _01251_ | _03759_;
	assign _03642_ = _03641_ | io_in[7];
	assign _03643_ = _03642_ | io_in[8];
	assign _03644_ = io_in[10] & ~_03643_;
	assign _03645_ = _00207_ & ~_01985_;
	assign _03646_ = _02698_ | _02207_;
	assign _03649_ = _03646_ | io_in[8];
	assign _03650_ = _03649_ | io_in[9];
	assign _03651_ = _06310_ & ~_03650_;
	assign _03652_ = _00709_ | _02207_;
	assign _03653_ = _03652_ | io_in[8];
	assign _03654_ = _03653_ | io_in[9];
	assign _03655_ = io_in[10] & ~_03654_;
	assign _03656_ = io_in[8] & ~_01573_;
	assign _03657_ = _01296_ | _02207_;
	assign _03658_ = _03657_ | io_in[9];
	assign _03660_ = _03658_ | io_in[10];
	assign _03661_ = _01985_ & ~_03660_;
	assign _03662_ = _01006_ | io_in[7];
	assign _03663_ = _03662_ | io_in[8];
	assign _03664_ = _03663_ | io_in[10];
	assign _03665_ = _01985_ & ~_03664_;
	assign _03666_ = io_in[10] & ~_01675_;
	assign _03667_ = _00632_ | io_in[8];
	assign _03668_ = _02096_ & ~_03667_;
	assign _03669_ = _01807_ | io_in[6];
	assign _03671_ = _03669_ | _02207_;
	assign _03672_ = _03671_ | io_in[9];
	assign _03673_ = _03672_ | io_in[10];
	assign _03674_ = _01985_ & ~_03673_;
	assign _03675_ = _02790_ | io_in[8];
	assign _03676_ = io_in[11] & ~_03675_;
	assign _03677_ = _02783_ | _02207_;
	assign _03678_ = _03677_ | _01208_;
	assign _03679_ = io_in[11] & ~_03678_;
	assign _03680_ = _02855_ | _03759_;
	assign _03682_ = _03680_ | io_in[8];
	assign _03683_ = _03682_ | _02096_;
	assign _03684_ = io_in[10] & ~_03683_;
	assign _03685_ = _01360_ | _03759_;
	assign _03686_ = _03685_ | io_in[7];
	assign _03687_ = io_in[10] & ~_03686_;
	assign _03688_ = _05456_ | io_in[6];
	assign _03689_ = _03688_ | io_in[7];
	assign _03690_ = _03689_ | _01208_;
	assign _03691_ = io_in[11] & ~_03690_;
	assign _03693_ = _02531_ | io_in[9];
	assign _03694_ = _03693_ | io_in[10];
	assign _03695_ = _01985_ & ~_03694_;
	assign _03696_ = _01469_ | _03759_;
	assign _03697_ = _03696_ | _01208_;
	assign _03698_ = _03697_ | _02096_;
	assign _03699_ = _01985_ & ~_03698_;
	assign _03700_ = io_in[11] & ~_03617_;
	assign _03701_ = _01348_ | io_in[9];
	assign _03702_ = io_in[11] & ~_03701_;
	assign _03704_ = _07410_ | io_in[7];
	assign _03705_ = _03704_ | io_in[8];
	assign _03706_ = _03705_ | io_in[10];
	assign _03707_ = _01985_ & ~_03706_;
	assign _03708_ = _01260_ | _06310_;
	assign _03709_ = io_in[11] & ~_03708_;
	assign _03710_ = _00566_ | io_in[7];
	assign _03711_ = _03710_ | _02096_;
	assign _03712_ = io_in[11] & ~_03711_;
	assign _03713_ = _00434_ | io_in[6];
	assign _03715_ = _03713_ | _02207_;
	assign _03716_ = _03715_ | io_in[8];
	assign _03717_ = _03716_ | io_in[9];
	assign _03718_ = io_in[11] & ~_03717_;
	assign _03719_ = _04103_ | _03759_;
	assign _03720_ = _03719_ | _02207_;
	assign _03721_ = _03720_ | _01208_;
	assign _03722_ = _03721_ | _02096_;
	assign _03723_ = _06310_ & ~_03722_;
	assign _03724_ = _07311_ | io_in[8];
	assign _03726_ = _03724_ | io_in[9];
	assign _03727_ = io_in[10] & ~_03726_;
	assign _03728_ = _05977_ | io_in[7];
	assign _03729_ = _03728_ | io_in[8];
	assign _03730_ = _03729_ | io_in[9];
	assign _03731_ = io_in[10] & ~_03730_;
	assign _03732_ = _01839_ | io_in[7];
	assign _03733_ = _03732_ | _02096_;
	assign _03734_ = _06310_ & ~_03733_;
	assign _03735_ = _00540_ | _02207_;
	assign _03737_ = _03735_ | _01208_;
	assign _03738_ = _03737_ | _02096_;
	assign _03739_ = _06310_ & ~_03738_;
	assign _03740_ = _06000_ | io_in[8];
	assign _03741_ = io_in[10] & ~_03740_;
	assign _03742_ = _00971_ | _03759_;
	assign _03743_ = _03742_ | io_in[8];
	assign _03744_ = _03743_ | io_in[9];
	assign _03745_ = _03744_ | io_in[10];
	assign _03746_ = _01985_ & ~_03745_;
	assign _03748_ = _00482_ | _03094_;
	assign _03749_ = _03748_ | _03759_;
	assign _03750_ = _03749_ | io_in[7];
	assign _03751_ = _03750_ | _02096_;
	assign _03752_ = _06310_ & ~_03751_;
	assign _03753_ = _01150_ | io_in[10];
	assign _03754_ = _01985_ & ~_03753_;
	assign _03755_ = _02793_ | _02207_;
	assign _03756_ = io_in[9] & ~_03755_;
	assign _03757_ = _00757_ | _03094_;
	assign _03760_ = _03757_ | io_in[6];
	assign _03761_ = _03760_ | io_in[7];
	assign _03762_ = _03761_ | _06310_;
	assign _03763_ = io_in[11] & ~_03762_;
	assign _03764_ = _07300_ | _03094_;
	assign _03765_ = _06310_ & ~_03764_;
	assign _03766_ = _01144_ | _01208_;
	assign _03767_ = _03766_ | _02096_;
	assign _03768_ = _06310_ & ~_03767_;
	assign _03769_ = _00368_ | io_in[6];
	assign _03771_ = _03769_ | _02207_;
	assign _03772_ = _03771_ | _01208_;
	assign _03773_ = _03772_ | io_in[9];
	assign _03774_ = io_in[10] & ~_03773_;
	assign _03775_ = _01392_ | _01208_;
	assign _03776_ = _01985_ & ~_03775_;
	assign _03777_ = _00759_ | _02207_;
	assign _03778_ = _03777_ | io_in[8];
	assign _03779_ = io_in[9] & ~_03778_;
	assign _03780_ = _01995_ | io_in[8];
	assign _03782_ = _03780_ | io_in[9];
	assign _03783_ = io_in[10] & ~_03782_;
	assign _03784_ = _01642_ | _01208_;
	assign _03785_ = _03784_ | io_in[9];
	assign _03786_ = io_in[10] & ~_03785_;
	assign _03787_ = _03558_ | _02096_;
	assign _03788_ = io_in[11] & ~_03787_;
	assign _03789_ = io_in[5] & ~_04845_;
	assign _03790_ = _02725_ | _01208_;
	assign _03791_ = _03790_ | _02096_;
	assign _03793_ = _06310_ & ~_03791_;
	assign _03794_ = _07283_ | io_in[5];
	assign _03795_ = _03794_ | io_in[6];
	assign _03796_ = _03795_ | _02207_;
	assign _03797_ = _03796_ | io_in[8];
	assign _03798_ = _03797_ | io_in[9];
	assign _03799_ = io_in[10] & ~_03798_;
	assign _03800_ = _07441_ & ~io_in[6];
	assign _03801_ = _00388_ | _03759_;
	assign _03802_ = _03801_ | io_in[7];
	assign _03804_ = _03802_ | io_in[8];
	assign _03805_ = _03804_ | io_in[9];
	assign _03806_ = io_in[11] & ~_03805_;
	assign _03807_ = _01506_ | io_in[9];
	assign _03808_ = io_in[11] & ~_03807_;
	assign _03809_ = _02752_ | _02207_;
	assign _03810_ = _03809_ | _01208_;
	assign _03811_ = io_in[10] & ~_03810_;
	assign _03812_ = _01894_ | _01208_;
	assign _03813_ = io_in[10] & ~_03812_;
	assign _03815_ = _01958_ | _03759_;
	assign _03816_ = _03815_ | _02207_;
	assign _03817_ = _03816_ | io_in[8];
	assign _03818_ = _03817_ | io_in[9];
	assign _03819_ = _06310_ & ~_03818_;
	assign _03820_ = _03725_ | io_in[6];
	assign _03821_ = _03820_ | _02207_;
	assign _03822_ = _03821_ | _01208_;
	assign _03823_ = _03822_ | io_in[9];
	assign _03824_ = io_in[11] & ~_03823_;
	assign _03826_ = _01430_ | _03094_;
	assign _03827_ = _03826_ | io_in[8];
	assign _03828_ = _03827_ | io_in[10];
	assign _03829_ = _01985_ & ~_03828_;
	assign _03830_ = _00472_ | _03094_;
	assign _03831_ = io_in[6] & ~_03830_;
	assign _03832_ = _00174_ | io_in[5];
	assign _03833_ = _03832_ | io_in[6];
	assign _03834_ = _03833_ | _02207_;
	assign _03835_ = _03834_ | _02096_;
	assign _03837_ = io_in[11] & ~_03835_;
	assign _03838_ = _00759_ | io_in[7];
	assign _03839_ = _03838_ | _02096_;
	assign _03840_ = _03839_ | _06310_;
	assign _03841_ = _01985_ & ~_03840_;
	assign _03842_ = _00694_ | _03094_;
	assign _03843_ = _03842_ | io_in[6];
	assign _03844_ = io_in[9] & ~_03843_;
	assign _03845_ = _03772_ | _02096_;
	assign _03846_ = _06310_ & ~_03845_;
	assign _03848_ = _02529_ | io_in[6];
	assign _03849_ = _03848_ | io_in[7];
	assign _03850_ = _03849_ | _02096_;
	assign _03851_ = _03850_ | _06310_;
	assign _03852_ = _01985_ & ~_03851_;
	assign _03853_ = _07273_ & ~_01985_;
	assign _03854_ = _01765_ | io_in[8];
	assign _03855_ = _03854_ | _02096_;
	assign _03856_ = _03855_ | io_in[10];
	assign _03857_ = _01985_ & ~_03856_;
	assign _03859_ = _01658_ | _02207_;
	assign _03860_ = _03859_ | io_in[8];
	assign _03861_ = _03860_ | io_in[9];
	assign _03862_ = _03861_ | io_in[10];
	assign _03863_ = io_in[11] & ~_03862_;
	assign _03864_ = _02982_ | _02207_;
	assign _03865_ = _03864_ | _01208_;
	assign _03866_ = _03865_ | _02096_;
	assign _03867_ = _03866_ | _06310_;
	assign _03868_ = _01985_ & ~_03867_;
	assign _03871_ = _07257_ | io_in[6];
	assign _03872_ = _03871_ | io_in[7];
	assign _03873_ = _03872_ | io_in[8];
	assign _03874_ = io_in[11] & ~_03873_;
	assign _03875_ = _01976_ | io_in[7];
	assign _03876_ = io_in[11] & ~_03875_;
	assign _03877_ = _01148_ | _03759_;
	assign _03878_ = _03877_ | _02207_;
	assign _03879_ = _03878_ | io_in[10];
	assign _03880_ = io_in[11] & ~_03879_;
	assign _03882_ = _01642_ | io_in[6];
	assign _03883_ = _03882_ | _02096_;
	assign _03884_ = _03883_ | io_in[10];
	assign _03885_ = _01985_ & ~_03884_;
	assign _03886_ = _03017_ & ~_01985_;
	assign _03887_ = _07435_ | _03759_;
	assign _03888_ = _03887_ | _06310_;
	assign _03889_ = io_in[11] & ~_03888_;
	assign _03890_ = _03493_ | io_in[6];
	assign _03891_ = _03890_ | _02207_;
	assign _03893_ = _03891_ | io_in[8];
	assign _03894_ = _03893_ | io_in[9];
	assign _03895_ = _03894_ | _06310_;
	assign _03896_ = _01985_ & ~_03895_;
	assign _03897_ = _07306_ | io_in[6];
	assign _03898_ = _03897_ | io_in[7];
	assign _03899_ = _03898_ | _06310_;
	assign _03900_ = io_in[11] & ~_03899_;
	assign _03901_ = _00497_ | _02096_;
	assign _03902_ = _03901_ | io_in[10];
	assign _03904_ = _01985_ & ~_03902_;
	assign _03905_ = _02324_ | io_in[8];
	assign _03906_ = _03905_ | io_in[9];
	assign _03907_ = io_in[11] & ~_03906_;
	assign _03908_ = _07378_ | _03759_;
	assign _03909_ = _03908_ | _02207_;
	assign _03910_ = _03909_ | _01208_;
	assign _03911_ = _06310_ & ~_03910_;
	assign _03912_ = _00281_ | _03759_;
	assign _03913_ = _03912_ | io_in[7];
	assign _03915_ = _03913_ | _01208_;
	assign _03916_ = _03915_ | io_in[10];
	assign _03917_ = io_in[11] & ~_03916_;
	assign _03918_ = _01538_ | _02207_;
	assign _03919_ = _03918_ | _01208_;
	assign _03920_ = _03919_ | io_in[9];
	assign _03921_ = io_in[11] & ~_03920_;
	assign _03922_ = _07436_ | _02207_;
	assign _03923_ = _03922_ | io_in[9];
	assign _03924_ = _06310_ & ~_03923_;
	assign _03926_ = _07313_ | _01208_;
	assign _03927_ = _03926_ | io_in[9];
	assign _03928_ = _06310_ & ~_03927_;
	assign _03929_ = _04912_ | _01208_;
	assign _03930_ = _03929_ | _02096_;
	assign _03931_ = io_in[10] & ~_03930_;
	assign _03932_ = _00407_ | io_in[6];
	assign _03933_ = _03932_ | io_in[7];
	assign _03934_ = _03933_ | _06310_;
	assign _03935_ = io_in[11] & ~_03934_;
	assign _03937_ = _04647_ | _03759_;
	assign _03938_ = _03937_ | _02207_;
	assign _03939_ = _03938_ | _01208_;
	assign _03940_ = _03939_ | io_in[9];
	assign _03941_ = io_in[10] & ~_03940_;
	assign _03942_ = _05456_ | _03759_;
	assign _03943_ = _03942_ | _01208_;
	assign _03944_ = io_in[9] & ~_03943_;
	assign _03945_ = _02798_ | io_in[7];
	assign _03946_ = _02096_ & ~_03945_;
	assign _03948_ = _07378_ | io_in[7];
	assign _03949_ = _03948_ | _01208_;
	assign _03950_ = _03949_ | io_in[9];
	assign _03951_ = io_in[10] & ~_03950_;
	assign _03952_ = _06864_ | _03094_;
	assign _03953_ = io_in[11] & ~_03952_;
	assign _03954_ = _07352_ | io_in[6];
	assign _03955_ = _03954_ | _02207_;
	assign _03956_ = _03955_ | _01208_;
	assign _03957_ = io_in[10] & ~_03956_;
	assign _03959_ = _03719_ | io_in[7];
	assign _03960_ = _03959_ | io_in[8];
	assign _03961_ = _06310_ & ~_03960_;
	assign _03962_ = _01334_ | _02207_;
	assign _03963_ = io_in[11] & ~_03962_;
	assign _03964_ = _01119_ | _01208_;
	assign _03965_ = _03964_ | io_in[9];
	assign _03966_ = io_in[10] & ~_03965_;
	assign _03967_ = _01038_ | _06310_;
	assign _03968_ = io_in[11] & ~_03967_;
	assign _03970_ = _02000_ | io_in[7];
	assign _03971_ = _03970_ | _02096_;
	assign _03972_ = _01985_ & ~_03971_;
	assign _03973_ = _02323_ | _02207_;
	assign _03974_ = _03973_ | io_in[8];
	assign _03975_ = _03974_ | io_in[9];
	assign _03976_ = io_in[11] & ~_03975_;
	assign _03977_ = _03908_ | io_in[7];
	assign _03978_ = _03977_ | _01208_;
	assign _03979_ = _03978_ | io_in[9];
	assign _03982_ = _01985_ & ~_03979_;
	assign _03983_ = _03583_ | io_in[7];
	assign _03984_ = _03983_ | _02096_;
	assign _03985_ = _03984_ | io_in[10];
	assign _03986_ = io_in[11] & ~_03985_;
	assign _03987_ = _06310_ & ~_02302_;
	assign _03988_ = _00987_ | io_in[6];
	assign _03989_ = _03988_ | _01208_;
	assign _03990_ = _03989_ | io_in[10];
	assign _03991_ = _01985_ & ~_03990_;
	assign _03993_ = _03090_ | _03759_;
	assign _03994_ = _03993_ | io_in[8];
	assign _03995_ = _03994_ | _02096_;
	assign _03996_ = _01985_ & ~_03995_;
	assign _03997_ = _03942_ | _02207_;
	assign _03998_ = _03997_ | _02096_;
	assign _03999_ = io_in[10] & ~_03998_;
	assign _04000_ = _00174_ | _03759_;
	assign _04001_ = _04000_ | io_in[7];
	assign _04002_ = _04001_ | _01208_;
	assign _04004_ = _04002_ | _02096_;
	assign _04005_ = _04004_ | _06310_;
	assign _04006_ = _01985_ & ~_04005_;
	assign _04007_ = _05278_ | _01208_;
	assign _04008_ = _04007_ | io_in[9];
	assign _04009_ = _04008_ | io_in[10];
	assign _04010_ = _01985_ & ~_04009_;
	assign _04011_ = _02471_ | _03759_;
	assign _04012_ = _04011_ | _02207_;
	assign _04013_ = _04012_ | io_in[8];
	assign _04015_ = _04013_ | io_in[9];
	assign _04016_ = io_in[10] & ~_04015_;
	assign _04017_ = _00658_ | _07422_;
	assign _04018_ = _04017_ | io_in[6];
	assign _04019_ = _04018_ | _02207_;
	assign _04020_ = _04019_ | io_in[8];
	assign _04021_ = _04020_ | _02096_;
	assign _04022_ = io_in[11] & ~_04021_;
	assign _04023_ = _03736_ | io_in[7];
	assign _04024_ = _04023_ | io_in[9];
	assign _04026_ = _04024_ | io_in[10];
	assign _04027_ = _01985_ & ~_04026_;
	assign _04028_ = _02809_ | io_in[9];
	assign _04029_ = _04028_ | io_in[10];
	assign _04030_ = _01985_ & ~_04029_;
	assign _04031_ = _03742_ | _02207_;
	assign _04032_ = _04031_ | io_in[8];
	assign _04033_ = _04032_ | _02096_;
	assign _04034_ = io_in[10] & ~_04033_;
	assign _04035_ = _07303_ | io_in[8];
	assign _04037_ = _04035_ | io_in[10];
	assign _04038_ = _01985_ & ~_04037_;
	assign _04039_ = _03230_ | io_in[8];
	assign _04040_ = io_in[9] & ~_04039_;
	assign _04041_ = _01046_ | _01208_;
	assign _04042_ = _04041_ | io_in[9];
	assign _04043_ = io_in[11] & ~_04042_;
	assign _04044_ = _01429_ | io_in[6];
	assign _04045_ = _04044_ | io_in[9];
	assign _04046_ = _04045_ | io_in[10];
	assign _04048_ = _01985_ & ~_04046_;
	assign _04049_ = _00131_ | _03094_;
	assign _04050_ = _04049_ | io_in[6];
	assign _04051_ = _04050_ | _02207_;
	assign _04052_ = _04051_ | _02096_;
	assign _04053_ = io_in[11] & ~_04052_;
	assign _04054_ = _01006_ | _03094_;
	assign _04055_ = _04054_ | _01208_;
	assign _04056_ = _01985_ & ~_04055_;
	assign _04057_ = _03977_ | io_in[8];
	assign _04059_ = io_in[9] & ~_04057_;
	assign _04060_ = _01651_ | io_in[7];
	assign _04061_ = _04060_ | io_in[8];
	assign _04062_ = io_in[10] & ~_04061_;
	assign _04063_ = _00374_ | io_in[7];
	assign _04064_ = _04063_ | _01208_;
	assign _04065_ = io_in[10] & ~_04064_;
	assign _04066_ = _00732_ | _03759_;
	assign _04067_ = _04066_ | io_in[7];
	assign _04068_ = _04067_ | _06310_;
	assign _04070_ = io_in[11] & ~_04068_;
	assign _04071_ = _02756_ | _01208_;
	assign _04072_ = _04071_ | io_in[10];
	assign _04073_ = io_in[11] & ~_04072_;
	assign _04074_ = _01039_ | _01208_;
	assign _04075_ = _06310_ & ~_04074_;
	assign _04076_ = io_in[10] & ~_02881_;
	assign _04077_ = _00493_ | io_in[6];
	assign _04078_ = _04077_ | io_in[7];
	assign _04079_ = _04078_ | _01208_;
	assign _04081_ = _04079_ | _02096_;
	assign _04082_ = _06310_ & ~_04081_;
	assign _04083_ = _04001_ | io_in[8];
	assign _04084_ = _04083_ | io_in[9];
	assign _04085_ = io_in[11] & ~_04084_;
	assign _04086_ = _07510_ | _02207_;
	assign _04087_ = _04086_ | _01208_;
	assign _04088_ = _04087_ | io_in[9];
	assign _04089_ = io_in[10] & ~_04088_;
	assign _04090_ = _02870_ | io_in[6];
	assign _04093_ = _04090_ | _02207_;
	assign _04094_ = _04093_ | _02096_;
	assign _04095_ = _06310_ & ~_04094_;
	assign _04096_ = _01730_ | io_in[7];
	assign _04097_ = _04096_ | io_in[8];
	assign _04098_ = io_in[11] & ~_04097_;
	assign _04099_ = _02847_ | _02096_;
	assign _04100_ = _01985_ & ~_04099_;
	assign _04101_ = _06310_ & ~_01566_;
	assign _04102_ = _02972_ | _01208_;
	assign _04104_ = io_in[9] & ~_04102_;
	assign _04105_ = _03057_ | _02207_;
	assign _04106_ = _04105_ | io_in[9];
	assign _04107_ = _06310_ & ~_04106_;
	assign _04108_ = _03627_ | io_in[7];
	assign _04109_ = io_in[10] & ~_04108_;
	assign _04110_ = _03809_ | _02096_;
	assign _04111_ = io_in[11] & ~_04110_;
	assign _04112_ = _01985_ & ~_02620_;
	assign _04113_ = _01215_ | io_in[7];
	assign _04115_ = _04113_ | io_in[8];
	assign _04116_ = _02096_ & ~_04115_;
	assign _04117_ = _00166_ | _03759_;
	assign _04118_ = _04117_ | io_in[8];
	assign _04119_ = _04118_ | _02096_;
	assign _04120_ = io_in[11] & ~_04119_;
	assign _04121_ = _00329_ | _01208_;
	assign _04122_ = _04121_ | _02096_;
	assign _04123_ = _06310_ & ~_04122_;
	assign _04124_ = _06609_ | _02207_;
	assign _04126_ = _04124_ | _06310_;
	assign _04127_ = io_in[11] & ~_04126_;
	assign _04128_ = _02813_ | io_in[9];
	assign _04129_ = io_in[10] & ~_04128_;
	assign _04130_ = _01985_ & ~_03251_;
	assign _04131_ = _07311_ | _02207_;
	assign _04132_ = _04131_ | io_in[8];
	assign _04133_ = _04132_ | io_in[9];
	assign _04134_ = io_in[11] & ~_04133_;
	assign _04135_ = _03680_ | io_in[7];
	assign _04137_ = _04135_ | _06310_;
	assign _04138_ = io_in[11] & ~_04137_;
	assign _04139_ = _01318_ | _02207_;
	assign _04140_ = _04139_ | _01208_;
	assign _04141_ = _01985_ & ~_04140_;
	assign _04142_ = _02998_ | _02207_;
	assign _04143_ = _04142_ | _02096_;
	assign _04144_ = _04143_ | _06310_;
	assign _04145_ = _01985_ & ~_04144_;
	assign _04146_ = _01067_ | io_in[9];
	assign _04148_ = _04146_ | io_in[10];
	assign _04149_ = io_in[11] & ~_04148_;
	assign _04150_ = _04513_ | io_in[6];
	assign _04151_ = _04150_ | _02207_;
	assign _04152_ = _04151_ | io_in[8];
	assign _04153_ = _04152_ | _02096_;
	assign _04154_ = _06310_ & ~_04153_;
	assign _04155_ = _03742_ | io_in[7];
	assign _04156_ = _04155_ | io_in[8];
	assign _04157_ = _04156_ | io_in[9];
	assign _04159_ = _01985_ & ~_04157_;
	assign _04160_ = _01541_ | _03094_;
	assign _04161_ = _04160_ | io_in[6];
	assign _04162_ = _02207_ & ~_04161_;
	assign _04163_ = _01226_ | _01208_;
	assign _04164_ = _04163_ | _02096_;
	assign _04165_ = _04164_ | _06310_;
	assign _04166_ = _01985_ & ~_04165_;
	assign _04167_ = _02285_ | _01208_;
	assign _04168_ = _04167_ | io_in[10];
	assign _04170_ = _01985_ & ~_04168_;
	assign _04171_ = _02778_ | io_in[7];
	assign _04172_ = _04171_ | io_in[8];
	assign _04173_ = _04172_ | _02096_;
	assign _04174_ = io_in[10] & ~_04173_;
	assign _04175_ = _02524_ | _01208_;
	assign _04176_ = _04175_ | _02096_;
	assign _04177_ = _01985_ & ~_04176_;
	assign _04178_ = _01042_ | io_in[6];
	assign _04179_ = _04178_ | _02207_;
	assign _04181_ = _04179_ | io_in[9];
	assign _04182_ = io_in[10] & ~_04181_;
	assign _04183_ = _03748_ | io_in[7];
	assign _04184_ = _04183_ | _01208_;
	assign _04185_ = _04184_ | io_in[9];
	assign _04186_ = io_in[10] & ~_04185_;
	assign _04187_ = _01732_ | _02096_;
	assign _04188_ = _01985_ & ~_04187_;
	assign _04189_ = _01013_ | io_in[8];
	assign _04190_ = _04189_ | io_in[9];
	assign _04192_ = _04190_ | io_in[10];
	assign _04193_ = _01985_ & ~_04192_;
	assign _04194_ = _00716_ | io_in[8];
	assign _04195_ = io_in[9] & ~_04194_;
	assign _04196_ = _00166_ | io_in[9];
	assign _04197_ = _04196_ | io_in[10];
	assign _04198_ = _01985_ & ~_04197_;
	assign _04199_ = _00391_ | _02207_;
	assign _04200_ = _04199_ | io_in[9];
	assign _04201_ = io_in[10] & ~_04200_;
	assign _04204_ = _03224_ | io_in[6];
	assign _04205_ = _04204_ | io_in[7];
	assign _04206_ = _04205_ | _01208_;
	assign _04207_ = _04206_ | _06310_;
	assign _04208_ = _01985_ & ~_04207_;
	assign _04209_ = _01195_ | io_in[7];
	assign _04210_ = _01985_ & ~_04209_;
	assign _04211_ = _00391_ | _03759_;
	assign _04212_ = _04211_ | io_in[7];
	assign _04213_ = _04212_ | io_in[8];
	assign _04215_ = _04213_ | _02096_;
	assign _04216_ = io_in[10] & ~_04215_;
	assign _04217_ = _03882_ | _01208_;
	assign _04218_ = _04217_ | _06310_;
	assign _04219_ = _01985_ & ~_04218_;
	assign _04220_ = _02479_ | _02096_;
	assign _04221_ = io_in[10] & ~_04220_;
	assign _04222_ = _01392_ | io_in[8];
	assign _04223_ = io_in[11] & ~_04222_;
	assign _04224_ = _04091_ | io_in[4];
	assign _04226_ = _04224_ | io_in[5];
	assign _04227_ = _04226_ | io_in[6];
	assign _04228_ = _04227_ | _01208_;
	assign _04229_ = _04228_ | io_in[10];
	assign _04230_ = io_in[11] & ~_04229_;
	assign _04231_ = _01200_ | _03759_;
	assign _04232_ = _04231_ | _01208_;
	assign _04233_ = _04232_ | io_in[9];
	assign _04234_ = io_in[10] & ~_04233_;
	assign _04235_ = _00889_ | io_in[7];
	assign _04237_ = _04235_ | _01208_;
	assign _04238_ = _04237_ | _02096_;
	assign _04239_ = _06310_ & ~_04238_;
	assign _04240_ = _01322_ | _01208_;
	assign _04241_ = _04240_ | _02096_;
	assign _04242_ = _04241_ | _06310_;
	assign _04243_ = _01985_ & ~_04242_;
	assign _04244_ = _00317_ | _03759_;
	assign _04245_ = _04244_ | _01208_;
	assign _04246_ = _04245_ | io_in[9];
	assign _04248_ = _04246_ | io_in[10];
	assign _04249_ = _01985_ & ~_04248_;
	assign _04250_ = _01386_ | _01208_;
	assign _04251_ = _04250_ | io_in[9];
	assign _04252_ = _06310_ & ~_04251_;
	assign _04253_ = _01283_ | io_in[8];
	assign _04254_ = io_in[9] & ~_04253_;
	assign _04255_ = _01879_ | io_in[8];
	assign _04256_ = _04255_ | _02096_;
	assign _04257_ = _04256_ | io_in[10];
	assign _04259_ = _01985_ & ~_04257_;
	assign _04260_ = _02976_ | _06310_;
	assign _04261_ = io_in[11] & ~_04260_;
	assign _04262_ = _01098_ | _01208_;
	assign _04263_ = _04262_ | _02096_;
	assign _04264_ = _06310_ & ~_04263_;
	assign _04265_ = _07280_ | _01208_;
	assign _04266_ = _04265_ | io_in[9];
	assign _04267_ = io_in[10] & ~_04266_;
	assign _04268_ = _07198_ | io_in[4];
	assign _04270_ = _04268_ | io_in[5];
	assign _04271_ = _04270_ | io_in[6];
	assign _04272_ = _04271_ | _02207_;
	assign _04273_ = _04272_ | _02096_;
	assign _04274_ = _04273_ | io_in[10];
	assign _04275_ = _01985_ & ~_04274_;
	assign _04276_ = _01335_ | io_in[8];
	assign _04277_ = _04276_ | _02096_;
	assign _04278_ = io_in[10] & ~_04277_;
	assign _04279_ = _03225_ | _02207_;
	assign _04281_ = _04279_ | _01208_;
	assign _04282_ = _04281_ | _02096_;
	assign _04283_ = _04282_ | _06310_;
	assign _04284_ = _01985_ & ~_04283_;
	assign _04285_ = io_in[11] & ~_02786_;
	assign _04286_ = _01631_ | io_in[7];
	assign _04287_ = _04286_ | _02096_;
	assign _04288_ = _01985_ & ~_04287_;
	assign _04289_ = _03802_ | _01208_;
	assign _04290_ = _04289_ | io_in[9];
	assign _04292_ = io_in[10] & ~_04290_;
	assign _04293_ = _07376_ | _02207_;
	assign _04294_ = _04293_ | io_in[8];
	assign _04295_ = _04294_ | _02096_;
	assign _04296_ = _06310_ & ~_04295_;
	assign _04297_ = _01135_ | _06310_;
	assign _04298_ = _01985_ & ~_04297_;
	assign _04299_ = _01058_ | _02207_;
	assign _04300_ = _04299_ | _01208_;
	assign _04301_ = _04300_ | _02096_;
	assign _04303_ = _04301_ | _06310_;
	assign _04304_ = _01985_ & ~_04303_;
	assign _04305_ = _02040_ | io_in[8];
	assign _04306_ = _04305_ | _02096_;
	assign _04307_ = io_in[10] & ~_04306_;
	assign _04308_ = _01068_ | _06310_;
	assign _04309_ = _01985_ & ~_04308_;
	assign _04310_ = _02484_ | _02207_;
	assign _04311_ = _04310_ | _02096_;
	assign _04312_ = io_in[10] & ~_04311_;
	assign _04315_ = _00985_ | io_in[6];
	assign _04316_ = _04315_ | io_in[9];
	assign _04317_ = _04316_ | io_in[10];
	assign _04318_ = _01985_ & ~_04317_;
	assign _04319_ = _01031_ | io_in[5];
	assign _04320_ = _04319_ | _03759_;
	assign _04321_ = _04320_ | io_in[7];
	assign _04322_ = _04321_ | io_in[8];
	assign _04323_ = _04322_ | io_in[9];
	assign _04324_ = io_in[10] & ~_04323_;
	assign _04326_ = _00198_ | io_in[5];
	assign _04327_ = _04326_ | _02207_;
	assign _04328_ = _04327_ | io_in[8];
	assign _04329_ = _04328_ | io_in[9];
	assign _04330_ = _01985_ & ~_04329_;
	assign _04331_ = _01215_ | io_in[8];
	assign _04332_ = io_in[10] & ~_04331_;
	assign _04333_ = _01175_ | io_in[9];
	assign _04334_ = _04333_ | _06310_;
	assign _04335_ = _01985_ & ~_04334_;
	assign _04337_ = io_in[11] & ~_01939_;
	assign _04338_ = _02029_ | io_in[5];
	assign _04339_ = _04338_ | _03759_;
	assign _04340_ = _04339_ | io_in[7];
	assign _04341_ = _04340_ | _06310_;
	assign _04342_ = io_in[11] & ~_04341_;
	assign _04343_ = _06000_ | io_in[9];
	assign _04344_ = io_in[11] & ~_04343_;
	assign _04345_ = _00987_ | io_in[7];
	assign _04346_ = _04345_ | io_in[9];
	assign _04348_ = _04346_ | io_in[10];
	assign _04349_ = _01985_ & ~_04348_;
	assign _04350_ = _07413_ | _02207_;
	assign _04351_ = _04350_ | _02096_;
	assign _04352_ = _04351_ | _06310_;
	assign _04353_ = _01985_ & ~_04352_;
	assign _04354_ = _00250_ | io_in[7];
	assign _04355_ = _04354_ | io_in[8];
	assign _04356_ = _04355_ | io_in[9];
	assign _04357_ = io_in[11] & ~_04356_;
	assign _04359_ = _07257_ | _03094_;
	assign _04360_ = _04359_ | _03759_;
	assign _04361_ = io_in[8] & ~_04360_;
	assign _04362_ = _01190_ | io_in[6];
	assign _04363_ = _04362_ | _02207_;
	assign _04364_ = _04363_ | _01208_;
	assign _04365_ = io_in[9] & ~_04364_;
	assign _04366_ = _03936_ | io_in[6];
	assign _04367_ = _04366_ | _02207_;
	assign _04368_ = _04367_ | io_in[9];
	assign _04370_ = io_in[11] & ~_04368_;
	assign _04371_ = _04044_ | _02207_;
	assign _04372_ = _04371_ | io_in[8];
	assign _04373_ = _04372_ | io_in[9];
	assign _04374_ = _06310_ & ~_04373_;
	assign _04375_ = _00501_ | io_in[6];
	assign _04376_ = _04375_ | _02207_;
	assign _04377_ = _04376_ | _01208_;
	assign _04378_ = _04377_ | io_in[9];
	assign _04379_ = io_in[10] & ~_04378_;
	assign _04381_ = _02778_ | io_in[6];
	assign _04382_ = _04381_ | _02207_;
	assign _04383_ = _04382_ | _01208_;
	assign _04384_ = _02096_ & ~_04383_;
	assign _04385_ = _01184_ | _02096_;
	assign _04386_ = _04385_ | io_in[10];
	assign _04387_ = io_in[11] & ~_04386_;
	assign _04388_ = _03315_ | io_in[7];
	assign _04389_ = _04388_ | _01208_;
	assign _04390_ = _04389_ | io_in[10];
	assign _04392_ = _01985_ & ~_04390_;
	assign _04393_ = _01698_ | io_in[6];
	assign _04394_ = _04393_ | _02207_;
	assign _04395_ = _04394_ | _01208_;
	assign _04396_ = _02096_ & ~_04395_;
	assign _04397_ = _07318_ | io_in[6];
	assign _04398_ = _04397_ | _02207_;
	assign _04399_ = _04398_ | io_in[8];
	assign _04400_ = _04399_ | _02096_;
	assign _04401_ = io_in[11] & ~_04400_;
	assign _04403_ = _03090_ | io_in[6];
	assign _04404_ = _04403_ | io_in[7];
	assign _04405_ = _04404_ | _01208_;
	assign _04406_ = io_in[10] & ~_04405_;
	assign _04407_ = _07436_ | io_in[7];
	assign _04408_ = _04407_ | io_in[8];
	assign _04409_ = io_in[10] & ~_04408_;
	assign _04410_ = _00169_ | io_in[7];
	assign _04411_ = _04410_ | io_in[8];
	assign _04412_ = _04411_ | _02096_;
	assign _04414_ = io_in[10] & ~_04412_;
	assign _04415_ = _07373_ | _01208_;
	assign _04416_ = _04415_ | _02096_;
	assign _04417_ = _04416_ | _06310_;
	assign _04418_ = _01985_ & ~_04417_;
	assign _04419_ = _01340_ | _02207_;
	assign _04420_ = _04419_ | io_in[8];
	assign _04421_ = _04420_ | _02096_;
	assign _04422_ = _04421_ | _06310_;
	assign _04423_ = _01985_ & ~_04422_;
	assign _04426_ = _00694_ | io_in[5];
	assign _04427_ = _04426_ | _03759_;
	assign _04428_ = _04427_ | io_in[7];
	assign _04429_ = _04428_ | _06310_;
	assign _04430_ = io_in[11] & ~_04429_;
	assign _04431_ = _00388_ | io_in[5];
	assign _04432_ = _04431_ | io_in[6];
	assign _04433_ = _04432_ | io_in[8];
	assign _04434_ = _04433_ | io_in[9];
	assign _04435_ = io_in[10] & ~_04434_;
	assign _04437_ = _07428_ | io_in[7];
	assign _04438_ = _04437_ | _02096_;
	assign _04439_ = io_in[10] & ~_04438_;
	assign _04440_ = _07403_ | io_in[7];
	assign _04441_ = _04440_ | _01208_;
	assign _04442_ = _04441_ | io_in[9];
	assign _04443_ = io_in[11] & ~_04442_;
	assign _04444_ = _03641_ | io_in[9];
	assign _04445_ = io_in[11] & ~_04444_;
	assign _04446_ = _00900_ | io_in[8];
	assign _04448_ = _04446_ | _02096_;
	assign _04449_ = io_in[10] & ~_04448_;
	assign _04450_ = _03748_ | io_in[6];
	assign _04451_ = _04450_ | io_in[8];
	assign _04452_ = _04451_ | _02096_;
	assign _04453_ = io_in[10] & ~_04452_;
	assign _04454_ = _05434_ | _01208_;
	assign _04455_ = _02096_ & ~_04454_;
	assign _04456_ = _01428_ | _01208_;
	assign _04457_ = _04456_ | io_in[9];
	assign _04459_ = _06310_ & ~_04457_;
	assign _04460_ = _03677_ | io_in[8];
	assign _04461_ = io_in[9] & ~_04460_;
	assign _04462_ = _03992_ | _03759_;
	assign _04463_ = _04462_ | io_in[7];
	assign _04464_ = _04463_ | io_in[8];
	assign _04465_ = _04464_ | _02096_;
	assign _04466_ = io_in[10] & ~_04465_;
	assign _04467_ = _01251_ | _02207_;
	assign _04468_ = _04467_ | _01208_;
	assign _04470_ = _02096_ & ~_04468_;
	assign _04471_ = _01225_ | io_in[7];
	assign _04472_ = _04471_ | _01208_;
	assign _04473_ = _04472_ | io_in[9];
	assign _04474_ = io_in[11] & ~_04473_;
	assign _04475_ = _01042_ | _02207_;
	assign _04476_ = _04475_ | _01208_;
	assign _04477_ = _04476_ | io_in[9];
	assign _04478_ = io_in[11] & ~_04477_;
	assign _04479_ = _01976_ | _02096_;
	assign _04481_ = io_in[11] & ~_04479_;
	assign _04482_ = _04235_ | io_in[8];
	assign _04483_ = _04482_ | io_in[9];
	assign _04484_ = io_in[10] & ~_04483_;
	assign _04485_ = _01982_ | io_in[7];
	assign _04486_ = _04485_ | _02096_;
	assign _04487_ = io_in[11] & ~_04486_;
	assign _04488_ = _00768_ | io_in[7];
	assign _04489_ = _04488_ | io_in[8];
	assign _04490_ = _04489_ | io_in[10];
	assign _04492_ = _01985_ & ~_04490_;
	assign _04493_ = _07389_ | _02207_;
	assign _04494_ = io_in[11] & ~_04493_;
	assign _04495_ = _04018_ | io_in[9];
	assign _04496_ = _04495_ | io_in[10];
	assign _04497_ = _01985_ & ~_04496_;
	assign _04498_ = _04017_ | _03759_;
	assign _04499_ = _04498_ | _02207_;
	assign _04500_ = _04499_ | _01208_;
	assign _04501_ = _04500_ | io_in[10];
	assign _04503_ = io_in[11] & ~_04501_;
	assign _04504_ = _01505_ | io_in[7];
	assign _04505_ = _04504_ | io_in[8];
	assign _04506_ = io_in[11] & ~_04505_;
	assign _04507_ = _05200_ | io_in[9];
	assign _04508_ = io_in[10] & ~_04507_;
	assign _04509_ = _06864_ | io_in[7];
	assign _04510_ = _04509_ | io_in[8];
	assign _04511_ = _04510_ | io_in[9];
	assign _04512_ = io_in[10] & ~_04511_;
	assign _04514_ = _00246_ | io_in[9];
	assign _04515_ = _04514_ | io_in[10];
	assign _04516_ = _01985_ & ~_04515_;
	assign _04517_ = _04516_ | _04512_;
	assign _04518_ = _04517_ | _04508_;
	assign _04519_ = _04518_ | _04506_;
	assign _04520_ = _04519_ | _04503_;
	assign _04521_ = _04520_ | _04497_;
	assign _04522_ = _04521_ | _04494_;
	assign _04523_ = _04522_ | _04492_;
	assign _04525_ = _04523_ | _04487_;
	assign _04526_ = _04525_ | _04484_;
	assign _04527_ = _04526_ | _04481_;
	assign _04528_ = _04527_ | _04478_;
	assign _04529_ = _04528_ | _04474_;
	assign _04530_ = _04529_ | _04470_;
	assign _04531_ = _04530_ | _04466_;
	assign _04532_ = _04531_ | _04461_;
	assign _04533_ = _04532_ | _04459_;
	assign _04534_ = _04533_ | _04455_;
	assign _04537_ = _04534_ | _04453_;
	assign _04538_ = _04537_ | _04449_;
	assign _04539_ = _04538_ | _04445_;
	assign _04540_ = _04539_ | _04443_;
	assign _04541_ = _04540_ | _04439_;
	assign _04542_ = _04541_ | _04435_;
	assign _04543_ = _04542_ | _04430_;
	assign _04544_ = _04543_ | _04423_;
	assign _04545_ = _04544_ | _04418_;
	assign _04546_ = _04545_ | _04414_;
	assign _04548_ = _04546_ | _04409_;
	assign _04549_ = _04548_ | _04406_;
	assign _04550_ = _04549_ | _04401_;
	assign _04551_ = _04550_ | _04396_;
	assign _04552_ = _04551_ | _04392_;
	assign _04553_ = _04552_ | _04387_;
	assign _04554_ = _04553_ | _04384_;
	assign _04555_ = _04554_ | _04379_;
	assign _04556_ = _04555_ | _04374_;
	assign _04557_ = _04556_ | _04370_;
	assign _04559_ = _04557_ | _04365_;
	assign _04560_ = _04559_ | _04361_;
	assign _04561_ = _04560_ | _04357_;
	assign _04562_ = _04561_ | _04353_;
	assign _04563_ = _04562_ | _04349_;
	assign _04564_ = _04563_ | _04344_;
	assign _04565_ = _04564_ | _04342_;
	assign _04566_ = _04565_ | _04337_;
	assign _04567_ = _04566_ | _04335_;
	assign _04568_ = _04567_ | _04332_;
	assign _04570_ = _04568_ | _04330_;
	assign _04571_ = _04570_ | _04324_;
	assign _04572_ = _04571_ | _04318_;
	assign _04573_ = _04572_ | _04312_;
	assign _04574_ = _04573_ | _04309_;
	assign _04575_ = _04574_ | _04307_;
	assign _04576_ = _04575_ | _04304_;
	assign _04577_ = _04576_ | _04298_;
	assign _04578_ = _04577_ | _04296_;
	assign _04579_ = _04578_ | _04292_;
	assign _04581_ = _04579_ | _04288_;
	assign _04582_ = _04581_ | _04285_;
	assign _04583_ = _04582_ | _04284_;
	assign _04584_ = _04583_ | _04278_;
	assign _04585_ = _04584_ | _04275_;
	assign _04586_ = _04585_ | _04267_;
	assign _04587_ = _04586_ | _07245_;
	assign _04588_ = _04587_ | _04264_;
	assign _04589_ = _04588_ | _04261_;
	assign _04590_ = _04589_ | _04259_;
	assign _04592_ = _04590_ | _04254_;
	assign _04593_ = _04592_ | _04252_;
	assign _04594_ = _04593_ | _04249_;
	assign _04595_ = _04594_ | _04243_;
	assign _04596_ = _04595_ | _04239_;
	assign _04597_ = _04596_ | _04234_;
	assign _04598_ = _04597_ | _04230_;
	assign _04599_ = _04598_ | _04223_;
	assign _04600_ = _04599_ | _04221_;
	assign _04601_ = _04600_ | _04219_;
	assign _04603_ = _04601_ | _04216_;
	assign _04604_ = _04603_ | _04210_;
	assign _04605_ = _04604_ | _04208_;
	assign _04606_ = _04605_ | _04201_;
	assign _04607_ = _04606_ | _04198_;
	assign _04608_ = _04607_ | _04195_;
	assign _04609_ = _04608_ | _04193_;
	assign _04610_ = _04609_ | _04188_;
	assign _04611_ = _04610_ | _04186_;
	assign _04612_ = _04611_ | _04182_;
	assign _04614_ = _04612_ | _04177_;
	assign _04615_ = _04614_ | _04174_;
	assign _04616_ = _04615_ | _04170_;
	assign _04617_ = _04616_ | _04166_;
	assign _04618_ = _04617_ | _03001_;
	assign _04619_ = _04618_ | _04162_;
	assign _04620_ = _04619_ | _04159_;
	assign _04621_ = _04620_ | _04154_;
	assign _04622_ = _04621_ | _04149_;
	assign _04623_ = _04622_ | _04145_;
	assign _04625_ = _04623_ | _04141_;
	assign _04626_ = _04625_ | _04138_;
	assign _04627_ = _04626_ | _02974_;
	assign _04628_ = _04627_ | _04134_;
	assign _04629_ = _04628_ | _04130_;
	assign _04630_ = _04629_ | _04129_;
	assign _04631_ = _04630_ | _04127_;
	assign _04632_ = _04631_ | _04123_;
	assign _04633_ = _04632_ | _04120_;
	assign _04634_ = _04633_ | _04116_;
	assign _04636_ = _04634_ | _04112_;
	assign _04637_ = _04636_ | _04111_;
	assign _04638_ = _04637_ | _04109_;
	assign _04639_ = _04638_ | _04107_;
	assign _04640_ = _04639_ | _04104_;
	assign _04641_ = _04640_ | _04101_;
	assign _04642_ = _04641_ | _04100_;
	assign _04643_ = _04642_ | _04098_;
	assign _04644_ = _04643_ | _04095_;
	assign _04645_ = _04644_ | _04089_;
	assign _04648_ = _04645_ | _04085_;
	assign _04649_ = _04648_ | _04082_;
	assign _04650_ = _04649_ | _04076_;
	assign _04651_ = _04650_ | _04075_;
	assign _04652_ = _04651_ | _04073_;
	assign _04653_ = _04652_ | _04070_;
	assign _04654_ = _04653_ | _04065_;
	assign _04655_ = _04654_ | _04062_;
	assign _04656_ = _04655_ | _04059_;
	assign _04657_ = _04656_ | _04056_;
	assign _04659_ = _04657_ | _04053_;
	assign _04660_ = _04659_ | _04048_;
	assign _04661_ = _04660_ | _04043_;
	assign _04662_ = _04661_ | _04040_;
	assign _04663_ = _04662_ | _04038_;
	assign _04664_ = _04663_ | _04034_;
	assign _04665_ = _04664_ | _04030_;
	assign _04666_ = _04665_ | _04027_;
	assign _04667_ = _04666_ | _04022_;
	assign _04668_ = _04667_ | _04016_;
	assign _04670_ = _04668_ | _04010_;
	assign _04671_ = _04670_ | _04006_;
	assign _04672_ = _04671_ | _03999_;
	assign _04673_ = _04672_ | _03996_;
	assign _04674_ = _04673_ | _03991_;
	assign _04675_ = _04674_ | _03987_;
	assign _04676_ = _04675_ | _03986_;
	assign _04677_ = _04676_ | _03982_;
	assign _04678_ = _04677_ | _03976_;
	assign _04679_ = _04678_ | _03972_;
	assign _04681_ = _04679_ | _03968_;
	assign _04682_ = _04681_ | _03966_;
	assign _04683_ = _04682_ | _03963_;
	assign _04684_ = _04683_ | _03961_;
	assign _04685_ = _04684_ | _03957_;
	assign _04686_ = _04685_ | _03953_;
	assign _04687_ = _04686_ | _03951_;
	assign _04688_ = _04687_ | _03946_;
	assign _04689_ = _04688_ | _03944_;
	assign _04690_ = _04689_ | _03941_;
	assign _04692_ = _04690_ | _03935_;
	assign _04693_ = _04692_ | _03931_;
	assign _04694_ = _04693_ | _03928_;
	assign _04695_ = _04694_ | _03924_;
	assign _04696_ = _04695_ | _03921_;
	assign _04697_ = _04696_ | _03917_;
	assign _04698_ = _04697_ | _03911_;
	assign _04699_ = _04698_ | _03907_;
	assign _04700_ = _04699_ | _03904_;
	assign _04701_ = _04700_ | _03900_;
	assign _04703_ = _04701_ | _03896_;
	assign _04704_ = _04703_ | _03889_;
	assign _04705_ = _04704_ | _03886_;
	assign _04706_ = _04705_ | _03885_;
	assign _04707_ = _04706_ | _03880_;
	assign _04708_ = _04707_ | _03876_;
	assign _04709_ = _04708_ | _03874_;
	assign _04710_ = _04709_ | _03868_;
	assign _04711_ = _04710_ | _03863_;
	assign _04712_ = _04711_ | _03857_;
	assign _04714_ = _04712_ | _03853_;
	assign _04715_ = _04714_ | _03852_;
	assign _04716_ = _04715_ | _03846_;
	assign _04717_ = _04716_ | _03844_;
	assign _04718_ = _04717_ | _03841_;
	assign _04719_ = _04718_ | _03837_;
	assign _04720_ = _04719_ | _03831_;
	assign _04721_ = _04720_ | _03829_;
	assign _04722_ = _04721_ | _03824_;
	assign _04723_ = _04722_ | _03819_;
	assign _04725_ = _04723_ | _03813_;
	assign _04726_ = _04725_ | _03811_;
	assign _04727_ = _04726_ | _03808_;
	assign _04728_ = _04727_ | _03806_;
	assign _04729_ = _04728_ | _03800_;
	assign _04730_ = _04729_ | _03799_;
	assign _04731_ = _04730_ | _03793_;
	assign _04732_ = _04731_ | _03789_;
	assign _04733_ = _04732_ | _03788_;
	assign _04734_ = _04733_ | _03786_;
	assign _04736_ = _04734_ | _03783_;
	assign _04737_ = _04736_ | _03779_;
	assign _04738_ = _04737_ | _03776_;
	assign _04739_ = _04738_ | _03774_;
	assign _04740_ = _04739_ | _03768_;
	assign _04741_ = _04740_ | _03765_;
	assign _04742_ = _04741_ | _03763_;
	assign _04743_ = _04742_ | _03756_;
	assign _04744_ = _04743_ | _03754_;
	assign _04745_ = _04744_ | _03752_;
	assign _04747_ = _04745_ | _03746_;
	assign _04748_ = _04747_ | _03741_;
	assign _04749_ = _04748_ | _03739_;
	assign _04750_ = _04749_ | _03734_;
	assign _04751_ = _04750_ | _03731_;
	assign _04752_ = _04751_ | _03727_;
	assign _04753_ = _04752_ | _03723_;
	assign _04754_ = _04753_ | _03718_;
	assign _04755_ = _04754_ | _03712_;
	assign _04756_ = _04755_ | _03709_;
	assign _04759_ = _04756_ | _03707_;
	assign _04760_ = _04759_ | _03702_;
	assign _04761_ = _04760_ | _03700_;
	assign _04762_ = _04761_ | _03699_;
	assign _04763_ = _04762_ | _03695_;
	assign _04764_ = _04763_ | _03691_;
	assign _04765_ = _04764_ | _03687_;
	assign _04766_ = _04765_ | _03684_;
	assign _04767_ = _04766_ | _03679_;
	assign _04768_ = _04767_ | _03676_;
	assign _04770_ = _04768_ | _03674_;
	assign _04771_ = _04770_ | _03668_;
	assign _04772_ = _04771_ | _03666_;
	assign _04773_ = _04772_ | _03665_;
	assign _04774_ = _04773_ | _03661_;
	assign _04775_ = _04774_ | _03656_;
	assign _04776_ = _04775_ | _03655_;
	assign _04777_ = _04776_ | _03651_;
	assign _04778_ = _04777_ | _02457_;
	assign _04779_ = _04778_ | _03645_;
	assign _04781_ = _04779_ | _03644_;
	assign _04782_ = _04781_ | _03640_;
	assign _04783_ = _04782_ | _03635_;
	assign _04784_ = _04783_ | _03632_;
	assign _04785_ = _04784_ | _03630_;
	assign _04786_ = _04785_ | _03626_;
	assign _04787_ = _04786_ | _03621_;
	assign _04788_ = _04787_ | _03618_;
	assign _04789_ = _04788_ | _03615_;
	assign _04790_ = _04789_ | _03610_;
	assign _04792_ = _04790_ | _03607_;
	assign _04793_ = _04792_ | _03604_;
	assign _04794_ = _04793_ | _03599_;
	assign _04795_ = _04794_ | _03594_;
	assign _04796_ = _04795_ | _03589_;
	assign _04797_ = _04796_ | _03586_;
	assign _04798_ = _04797_ | _03582_;
	assign _04799_ = _04798_ | _02327_;
	assign _04800_ = _04799_ | _03578_;
	assign _04801_ = _04800_ | _03576_;
	assign _04803_ = _04801_ | _03573_;
	assign _04804_ = _04803_ | _03567_;
	assign _04805_ = _04804_ | _03564_;
	assign _04806_ = _04805_ | _03561_;
	assign _04807_ = _04806_ | _03557_;
	assign _04808_ = _04807_ | _03553_;
	assign _04809_ = _04808_ | _03547_;
	assign _04810_ = _04809_ | _03546_;
	assign _04811_ = _04810_ | _03543_;
	assign _04812_ = _04811_ | _03539_;
	assign \mchip.val [2] = _04812_ | _03532_;
	assign _04814_ = _00247_ | io_in[8];
	assign _04815_ = _04814_ | _02096_;
	assign _04816_ = io_in[10] & ~_04815_;
	assign _04817_ = _00823_ | _03759_;
	assign _04818_ = _04817_ | io_in[8];
	assign _04819_ = _04818_ | _02096_;
	assign _04820_ = _04819_ | io_in[10];
	assign _04821_ = _01985_ & ~_04820_;
	assign _04822_ = _07252_ | io_in[8];
	assign _04824_ = _04822_ | io_in[9];
	assign _04825_ = io_in[10] & ~_04824_;
	assign _04826_ = _04231_ | io_in[7];
	assign _04827_ = _04826_ | io_in[8];
	assign _04828_ = _04827_ | io_in[9];
	assign _04829_ = io_in[11] & ~_04828_;
	assign _04830_ = _01496_ | io_in[6];
	assign _04831_ = _04830_ | io_in[7];
	assign _04832_ = _04831_ | _02096_;
	assign _04833_ = _04832_ | _06310_;
	assign _04835_ = _01985_ & ~_04833_;
	assign _04836_ = _01335_ | _02096_;
	assign _04837_ = io_in[11] & ~_04836_;
	assign _04838_ = _01469_ | io_in[7];
	assign _04839_ = _04838_ | io_in[8];
	assign _04840_ = io_in[9] & ~_04839_;
	assign _04841_ = _03002_ | _02207_;
	assign _04842_ = _04841_ | io_in[9];
	assign _04843_ = _06310_ & ~_04842_;
	assign _04844_ = _01596_ | _03759_;
	assign _04846_ = _04844_ | io_in[7];
	assign _04847_ = _04846_ | _01208_;
	assign _04848_ = _04847_ | io_in[9];
	assign _04849_ = io_in[10] & ~_04848_;
	assign _04850_ = _01411_ | _03759_;
	assign _04851_ = _04850_ | _02207_;
	assign _04852_ = _04851_ | _02096_;
	assign _04853_ = _06310_ & ~_04852_;
	assign _04854_ = _04403_ | _02207_;
	assign _04855_ = _04854_ | _01208_;
	assign _04857_ = _06310_ & ~_04855_;
	assign _04858_ = _03571_ | _06310_;
	assign _04859_ = _01985_ & ~_04858_;
	assign _04860_ = _07142_ | _02207_;
	assign _04861_ = _04860_ | io_in[9];
	assign _04862_ = io_in[11] & ~_04861_;
	assign _04863_ = _01781_ | _01208_;
	assign _04864_ = io_in[11] & ~_04863_;
	assign _04865_ = _01340_ | _03759_;
	assign _04866_ = _04865_ | io_in[7];
	assign _04869_ = _04866_ | _01208_;
	assign _04870_ = _04869_ | _02096_;
	assign _04871_ = _04870_ | io_in[10];
	assign _04872_ = _01985_ & ~_04871_;
	assign _04873_ = _01327_ | _02096_;
	assign _04874_ = io_in[10] & ~_04873_;
	assign _04875_ = _01017_ | _01208_;
	assign _04876_ = _04875_ | io_in[9];
	assign _04877_ = _04876_ | io_in[10];
	assign _04878_ = _01985_ & ~_04877_;
	assign _04880_ = _01985_ & ~_03257_;
	assign _04881_ = _04058_ | _02207_;
	assign _04882_ = _04881_ | _01208_;
	assign _04883_ = _02096_ & ~_04882_;
	assign _04884_ = _07259_ | io_in[5];
	assign _04885_ = _04884_ | io_in[6];
	assign _04886_ = _04885_ | _02207_;
	assign _04887_ = _04886_ | _06310_;
	assign _04888_ = io_in[11] & ~_04887_;
	assign _04889_ = _03018_ | io_in[7];
	assign _04891_ = _04889_ | io_in[8];
	assign _04892_ = _04891_ | _02096_;
	assign _04893_ = io_in[11] & ~_04892_;
	assign _04894_ = _03055_ | _06310_;
	assign _04895_ = _01985_ & ~_04894_;
	assign _04896_ = _03777_ | _01208_;
	assign _04897_ = _04896_ | io_in[9];
	assign _04898_ = io_in[10] & ~_04897_;
	assign _04899_ = _03237_ | io_in[8];
	assign _04900_ = _04899_ | io_in[10];
	assign _04902_ = _01985_ & ~_04900_;
	assign _04903_ = _05489_ | io_in[6];
	assign _04904_ = _04903_ | io_in[7];
	assign _04905_ = _04904_ | io_in[8];
	assign _04906_ = _04905_ | io_in[9];
	assign _04907_ = io_in[11] & ~_04906_;
	assign _04908_ = _01125_ | _03759_;
	assign _04909_ = _04908_ | _02207_;
	assign _04910_ = _04909_ | io_in[8];
	assign _04911_ = _04910_ | _02096_;
	assign _04913_ = _06310_ & ~_04911_;
	assign _04914_ = _06520_ | io_in[5];
	assign _04915_ = _04914_ | io_in[6];
	assign _04916_ = _04915_ | _06310_;
	assign _04917_ = io_in[11] & ~_04916_;
	assign _04918_ = _00317_ | _03094_;
	assign _04919_ = _04918_ | _01208_;
	assign _04920_ = _06310_ & ~_04919_;
	assign _04921_ = _02355_ | io_in[8];
	assign _04922_ = _04921_ | io_in[9];
	assign _04924_ = io_in[10] & ~_04922_;
	assign _04925_ = _03106_ | _01208_;
	assign _04926_ = _06310_ & ~_04925_;
	assign _04927_ = _01408_ | _01208_;
	assign _04928_ = io_in[10] & ~_04927_;
	assign _04929_ = _00245_ | io_in[6];
	assign _04930_ = _04929_ | io_in[7];
	assign _04931_ = _04930_ | _01208_;
	assign _04932_ = _04931_ | io_in[9];
	assign _04933_ = _04932_ | _06310_;
	assign _04935_ = _01985_ & ~_04933_;
	assign _04936_ = io_in[6] & ~_02768_;
	assign _04937_ = _02819_ | _02207_;
	assign _04938_ = _04937_ | _01208_;
	assign _04939_ = _02096_ & ~_04938_;
	assign _04940_ = _01985_ & ~_01159_;
	assign _04941_ = _01438_ | _02207_;
	assign _04942_ = _04941_ | _01208_;
	assign _04943_ = _04942_ | io_in[10];
	assign _04944_ = io_in[11] & ~_04943_;
	assign _04946_ = _01148_ | io_in[6];
	assign _04947_ = _04946_ | io_in[7];
	assign _04948_ = io_in[11] & ~_04947_;
	assign _04949_ = _03747_ | _02207_;
	assign _04950_ = _04949_ | io_in[8];
	assign _04951_ = io_in[10] & ~_04950_;
	assign _04952_ = _02813_ | io_in[7];
	assign _04953_ = _04952_ | _01208_;
	assign _04954_ = _04953_ | _02096_;
	assign _04955_ = _01985_ & ~_04954_;
	assign _04957_ = _01958_ | io_in[7];
	assign _04958_ = _04957_ | io_in[8];
	assign _04959_ = _04958_ | _02096_;
	assign _04960_ = io_in[11] & ~_04959_;
	assign _04961_ = _07402_ | _02207_;
	assign _04962_ = _04961_ | _02096_;
	assign _04963_ = _04962_ | io_in[10];
	assign _04964_ = io_in[11] & ~_04963_;
	assign _04965_ = _01451_ | _01208_;
	assign _04966_ = _04965_ | _02096_;
	assign _04968_ = _04966_ | _06310_;
	assign _04969_ = io_in[11] & ~_04968_;
	assign _04970_ = _01101_ | io_in[9];
	assign _04971_ = _04970_ | io_in[10];
	assign _04972_ = _01985_ & ~_04971_;
	assign _04973_ = _03736_ | _02207_;
	assign _04974_ = _04973_ | io_in[9];
	assign _04975_ = _04974_ | io_in[10];
	assign _04976_ = _01985_ & ~_04975_;
	assign _04977_ = _01807_ | _03094_;
	assign _04980_ = _04977_ | _02207_;
	assign _04981_ = _04980_ | _01208_;
	assign _04982_ = io_in[11] & ~_04981_;
	assign _04983_ = _04384_ & ~_06310_;
	assign _04984_ = _03993_ | _06310_;
	assign _04985_ = io_in[11] & ~_04984_;
	assign _04986_ = _01919_ | _03759_;
	assign _04987_ = _04986_ | _02207_;
	assign _04988_ = _04987_ | io_in[8];
	assign _04989_ = _04988_ | _02096_;
	assign _04991_ = io_in[10] & ~_04989_;
	assign _04992_ = _01380_ | io_in[7];
	assign _04993_ = _04992_ | io_in[8];
	assign _04994_ = _04993_ | _02096_;
	assign _04995_ = io_in[11] & ~_04994_;
	assign _04996_ = _01282_ | io_in[7];
	assign _04997_ = _04996_ | _01208_;
	assign _04998_ = _04997_ | _06310_;
	assign _04999_ = _01985_ & ~_04998_;
	assign _05000_ = _02956_ & ~io_in[7];
	assign _05002_ = io_in[9] & ~_01531_;
	assign _05003_ = _04908_ | io_in[7];
	assign _05004_ = _05003_ | _01208_;
	assign _05005_ = _05004_ | io_in[9];
	assign _05006_ = _05005_ | io_in[10];
	assign _05007_ = io_in[11] & ~_05006_;
	assign _05008_ = _01421_ | io_in[7];
	assign _05009_ = _05008_ | _06310_;
	assign _05010_ = io_in[11] & ~_05009_;
	assign _05011_ = _01886_ | _02096_;
	assign _05013_ = _05011_ | _06310_;
	assign _05014_ = _01985_ & ~_05013_;
	assign _05015_ = _04978_ | _02207_;
	assign _05016_ = _05015_ | _01208_;
	assign _05017_ = _02096_ & ~_05016_;
	assign _05018_ = _02905_ & ~_06310_;
	assign _05019_ = _03942_ | io_in[8];
	assign _05020_ = _05019_ | _02096_;
	assign _05021_ = io_in[10] & ~_05020_;
	assign _05022_ = _02272_ | _01208_;
	assign _05024_ = _05022_ | io_in[9];
	assign _05025_ = _05024_ | io_in[10];
	assign _05026_ = _01985_ & ~_05025_;
	assign _05027_ = _02501_ | _02207_;
	assign _05028_ = _05027_ | _01208_;
	assign _05029_ = _05028_ | io_in[9];
	assign _05030_ = io_in[10] & ~_05029_;
	assign _05031_ = _03526_ | _07422_;
	assign _05032_ = _05031_ | io_in[5];
	assign _05033_ = _05032_ | io_in[6];
	assign _05035_ = _05033_ | io_in[7];
	assign _05036_ = _05035_ | _06310_;
	assign _05037_ = io_in[11] & ~_05036_;
	assign _05038_ = _03891_ | _01208_;
	assign _05039_ = _05038_ | io_in[9];
	assign _05040_ = _05039_ | _06310_;
	assign _05041_ = _01985_ & ~_05040_;
	assign _05042_ = _00708_ | io_in[6];
	assign _05043_ = _05042_ | io_in[8];
	assign _05044_ = _05043_ | io_in[9];
	assign _05046_ = io_in[11] & ~_05044_;
	assign _05047_ = _02485_ | io_in[8];
	assign _05048_ = io_in[10] & ~_05047_;
	assign _05049_ = _00988_ | io_in[8];
	assign _05050_ = _05049_ | _02096_;
	assign _05051_ = _01985_ & ~_05050_;
	assign _05052_ = _04393_ | io_in[8];
	assign _05053_ = _05052_ | _02096_;
	assign _05054_ = _05053_ | io_in[10];
	assign _05055_ = _01985_ & ~_05054_;
	assign _05057_ = _02497_ | io_in[7];
	assign _05058_ = _05057_ | _02096_;
	assign _05059_ = io_in[11] & ~_05058_;
	assign _05060_ = _03908_ | _01208_;
	assign _05061_ = _05060_ | io_in[9];
	assign _05062_ = _06310_ & ~_05061_;
	assign _05063_ = _01348_ | _02207_;
	assign _05064_ = _05063_ | io_in[9];
	assign _05065_ = _06310_ & ~_05064_;
	assign _05066_ = _02312_ | _02207_;
	assign _05068_ = _05066_ | io_in[9];
	assign _05069_ = _05068_ | io_in[10];
	assign _05070_ = _01985_ & ~_05069_;
	assign _05071_ = _04155_ | io_in[9];
	assign _05072_ = io_in[10] & ~_05071_;
	assign _05073_ = _01977_ | _06310_;
	assign _05074_ = _01985_ & ~_05073_;
	assign _05075_ = _06643_ | _03094_;
	assign _05076_ = _05075_ | _03759_;
	assign _05077_ = _05076_ | _02207_;
	assign _05079_ = _05077_ | _01208_;
	assign _05080_ = _05079_ | _06310_;
	assign _05081_ = _01985_ & ~_05080_;
	assign _05082_ = _04059_ & ~_06310_;
	assign _05083_ = _01213_ | _03094_;
	assign _05084_ = _05083_ | io_in[7];
	assign _05085_ = _05084_ | _06310_;
	assign _05086_ = io_in[11] & ~_05085_;
	assign _05087_ = _07358_ | _03094_;
	assign _05088_ = io_in[7] & ~_05087_;
	assign _05091_ = _07289_ | _03759_;
	assign _05092_ = _05091_ | _02207_;
	assign _05093_ = _05092_ | _02096_;
	assign _05094_ = _05093_ | io_in[10];
	assign _05095_ = io_in[11] & ~_05094_;
	assign _05096_ = _07335_ | _03094_;
	assign _05097_ = _05096_ | _03759_;
	assign _05098_ = _05097_ | _02207_;
	assign _05099_ = _02096_ & ~_05098_;
	assign _05100_ = _07358_ | io_in[6];
	assign _05102_ = _05100_ | _02207_;
	assign _05103_ = _05102_ | io_in[8];
	assign _05104_ = _05103_ | _02096_;
	assign _05105_ = io_in[10] & ~_05104_;
	assign _05106_ = _00559_ | _03759_;
	assign _05107_ = _05106_ | _02207_;
	assign _05108_ = _05107_ | _01208_;
	assign _05109_ = _05108_ | io_in[9];
	assign _05110_ = io_in[11] & ~_05109_;
	assign _05111_ = _01003_ | _01208_;
	assign _05113_ = _02096_ & ~_05111_;
	assign _05114_ = _02567_ | _02207_;
	assign _05115_ = _05114_ | _06310_;
	assign _05116_ = io_in[11] & ~_05115_;
	assign _05117_ = _00878_ | _03094_;
	assign _05118_ = _05117_ | io_in[7];
	assign _05119_ = _05118_ | io_in[9];
	assign _05120_ = io_in[10] & ~_05119_;
	assign _05121_ = _04440_ | io_in[8];
	assign _05122_ = io_in[9] & ~_05121_;
	assign _05124_ = _03749_ | _02207_;
	assign _05125_ = _05124_ | io_in[8];
	assign _05126_ = io_in[11] & ~_05125_;
	assign _05127_ = _01758_ | _02096_;
	assign _05128_ = io_in[11] & ~_05127_;
	assign _05129_ = _00439_ | _03759_;
	assign _05130_ = _05129_ | _02096_;
	assign _05131_ = _05130_ | io_in[10];
	assign _05132_ = io_in[11] & ~_05131_;
	assign _05133_ = _01652_ | _02207_;
	assign _05135_ = _05133_ | _01208_;
	assign _05136_ = _05135_ | _02096_;
	assign _05137_ = _06310_ & ~_05136_;
	assign _05138_ = _01871_ | io_in[7];
	assign _05139_ = _05138_ | _01208_;
	assign _05140_ = io_in[11] & ~_05139_;
	assign _05141_ = _03057_ | _03759_;
	assign _05142_ = _05141_ | io_in[8];
	assign _05143_ = _05142_ | io_in[9];
	assign _05144_ = io_in[10] & ~_05143_;
	assign _05146_ = _01538_ | io_in[8];
	assign _05147_ = _05146_ | io_in[10];
	assign _05148_ = _01985_ & ~_05147_;
	assign _05149_ = _01026_ | _06310_;
	assign _05150_ = _01985_ & ~_05149_;
	assign _05151_ = _01079_ | io_in[7];
	assign _05152_ = _05151_ | io_in[8];
	assign _05153_ = _05152_ | _02096_;
	assign _05154_ = io_in[10] & ~_05153_;
	assign _05155_ = _02798_ | io_in[6];
	assign _05157_ = _05155_ | _02096_;
	assign _05158_ = _01985_ & ~_05157_;
	assign _05159_ = _00383_ | _07422_;
	assign _05160_ = _05159_ | _03759_;
	assign _05161_ = _05160_ | _02207_;
	assign _05162_ = _05161_ | _02096_;
	assign _05163_ = _05162_ | io_in[10];
	assign _05164_ = _01985_ & ~_05163_;
	assign _05165_ = _01128_ | io_in[9];
	assign _05166_ = _05165_ | io_in[10];
	assign _05168_ = io_in[11] & ~_05166_;
	assign _05169_ = _00449_ | io_in[7];
	assign _05170_ = _01985_ & ~_05169_;
	assign _05171_ = _01112_ | io_in[9];
	assign _05172_ = _01985_ & ~_05171_;
	assign _05173_ = _03160_ | _03759_;
	assign _05174_ = _05173_ | _02207_;
	assign _05175_ = _05174_ | _01208_;
	assign _05176_ = _05175_ | _02096_;
	assign _05177_ = _06310_ & ~_05176_;
	assign _05179_ = _00900_ | _01208_;
	assign _05180_ = _05179_ | _02096_;
	assign _05181_ = _06310_ & ~_05180_;
	assign _05182_ = _01758_ | io_in[8];
	assign _05183_ = io_in[11] & ~_05182_;
	assign _05184_ = _04105_ | io_in[8];
	assign _05185_ = _05184_ | _02096_;
	assign _05186_ = io_in[10] & ~_05185_;
	assign _05187_ = _01139_ | _01208_;
	assign _05188_ = _06310_ & ~_05187_;
	assign _05190_ = _02971_ | _03094_;
	assign _05191_ = _05190_ | _03759_;
	assign _05192_ = _05191_ | io_in[7];
	assign _05193_ = _05192_ | _06310_;
	assign _05194_ = io_in[11] & ~_05193_;
	assign _05195_ = _06720_ | _03094_;
	assign _05196_ = _05195_ | io_in[6];
	assign _05197_ = _02207_ & ~_05196_;
	assign _05198_ = _01125_ | _02207_;
	assign _05199_ = _05198_ | _01208_;
	assign _05202_ = _05199_ | _02096_;
	assign _05203_ = _05202_ | _06310_;
	assign _05204_ = io_in[11] & ~_05203_;
	assign _05205_ = _05027_ | _06310_;
	assign _05206_ = io_in[11] & ~_05205_;
	assign _05207_ = _04117_ | _02207_;
	assign _05208_ = _05207_ | _01208_;
	assign _05209_ = _05208_ | _02096_;
	assign _05210_ = _06310_ & ~_05209_;
	assign _05211_ = _00981_ | _01208_;
	assign _05213_ = _05211_ | _06310_;
	assign _05214_ = _01985_ & ~_05213_;
	assign _05215_ = _01856_ | io_in[7];
	assign _05216_ = _05215_ | _01208_;
	assign _05217_ = io_in[10] & ~_05216_;
	assign _05218_ = _04865_ | io_in[8];
	assign _05219_ = _05218_ | io_in[9];
	assign _05220_ = _05219_ | io_in[10];
	assign _05221_ = _01985_ & ~_05220_;
	assign _05222_ = _01445_ | io_in[8];
	assign _05224_ = _05222_ | io_in[9];
	assign _05225_ = io_in[11] & ~_05224_;
	assign _05226_ = _02571_ | _01208_;
	assign _05227_ = _05226_ | _02096_;
	assign _05228_ = _05227_ | _06310_;
	assign _05229_ = _01985_ & ~_05228_;
	assign _05230_ = _02040_ | _02207_;
	assign _05231_ = _05230_ | _01208_;
	assign _05232_ = _05231_ | _02096_;
	assign _05233_ = _06310_ & ~_05232_;
	assign _05235_ = _02218_ | _03759_;
	assign _05236_ = _05235_ | _02207_;
	assign _05237_ = _05236_ | io_in[8];
	assign _05238_ = _05237_ | _02096_;
	assign _05239_ = _05238_ | io_in[10];
	assign _05240_ = _01985_ & ~_05239_;
	assign _05241_ = _06720_ | _03759_;
	assign _05242_ = _05241_ | io_in[7];
	assign _05243_ = _05242_ | io_in[8];
	assign _05244_ = _05243_ | io_in[9];
	assign _05246_ = _06310_ & ~_05244_;
	assign _05247_ = _03549_ | _02207_;
	assign _05248_ = _05247_ | io_in[8];
	assign _05249_ = _05248_ | io_in[9];
	assign _05250_ = io_in[10] & ~_05249_;
	assign _05251_ = _07356_ | _03094_;
	assign _05252_ = _05251_ | io_in[7];
	assign _05253_ = _05252_ | io_in[8];
	assign _05254_ = _05253_ | _02096_;
	assign _05255_ = io_in[10] & ~_05254_;
	assign _05257_ = _01849_ | io_in[5];
	assign _05258_ = _05257_ | _02207_;
	assign _05259_ = _05258_ | io_in[8];
	assign _05260_ = _05259_ | _02096_;
	assign _05261_ = io_in[10] & ~_05260_;
	assign _05262_ = _05241_ | _02207_;
	assign _05263_ = _05262_ | _02096_;
	assign _05264_ = _05263_ | _06310_;
	assign _05265_ = _01985_ & ~_05264_;
	assign _05266_ = _00709_ | io_in[6];
	assign _05268_ = _05266_ | io_in[7];
	assign _05269_ = _05268_ | _01208_;
	assign _05270_ = _05269_ | io_in[9];
	assign _05271_ = io_in[10] & ~_05270_;
	assign _05272_ = _01251_ | _01208_;
	assign _05273_ = _05272_ | io_in[10];
	assign _05274_ = _01985_ & ~_05273_;
	assign _05275_ = _01578_ | _02096_;
	assign _05276_ = io_in[10] & ~_05275_;
	assign _05277_ = _00757_ | io_in[5];
	assign _05279_ = _05277_ | io_in[6];
	assign _05280_ = _05279_ | io_in[7];
	assign _05281_ = _05280_ | _01208_;
	assign _05282_ = _05281_ | _02096_;
	assign _05283_ = _05282_ | _06310_;
	assign _05284_ = _01985_ & ~_05283_;
	assign _05285_ = _03912_ | _02207_;
	assign _05286_ = io_in[11] & ~_05285_;
	assign _05287_ = _01856_ | io_in[8];
	assign _05288_ = _05287_ | io_in[10];
	assign _05290_ = _01985_ & ~_05288_;
	assign _05291_ = _00336_ | _03759_;
	assign _05292_ = _05291_ | _02207_;
	assign _05293_ = _05292_ | io_in[8];
	assign _05294_ = _05293_ | io_in[9];
	assign _05295_ = io_in[11] & ~_05294_;
	assign _05296_ = _05159_ | io_in[6];
	assign _05297_ = _05296_ | _02207_;
	assign _05298_ = _05297_ | io_in[8];
	assign _05299_ = _05298_ | _02096_;
	assign _05301_ = io_in[10] & ~_05299_;
	assign _05302_ = _04580_ | _03759_;
	assign _05303_ = _05302_ | io_in[7];
	assign _05304_ = _05303_ | io_in[8];
	assign _05305_ = _05304_ | io_in[9];
	assign _05306_ = io_in[11] & ~_05305_;
	assign _05307_ = _00131_ | _02207_;
	assign _05308_ = _05307_ | _01208_;
	assign _05309_ = _05308_ | _02096_;
	assign _05310_ = _05309_ | _06310_;
	assign _05313_ = io_in[11] & ~_05310_;
	assign _05314_ = _04276_ | io_in[9];
	assign _05315_ = io_in[10] & ~_05314_;
	assign _05316_ = _01362_ | _01208_;
	assign _05317_ = io_in[10] & ~_05316_;
	assign _05318_ = _05100_ | io_in[7];
	assign _05319_ = _05318_ | _01208_;
	assign _05320_ = _05319_ | io_in[9];
	assign _05321_ = io_in[10] & ~_05320_;
	assign _05322_ = _00232_ | _02207_;
	assign _05324_ = _05322_ | _01208_;
	assign _05325_ = _05324_ | io_in[9];
	assign _05326_ = io_in[10] & ~_05325_;
	assign _05327_ = _03632_ & ~_01985_;
	assign _05328_ = _03183_ | io_in[7];
	assign _05329_ = _05328_ | io_in[9];
	assign _05330_ = io_in[10] & ~_05329_;
	assign _05331_ = _01698_ | io_in[7];
	assign _05332_ = _05331_ | io_in[8];
	assign _05333_ = _05332_ | io_in[10];
	assign _05335_ = _01985_ & ~_05333_;
	assign _05336_ = _04228_ | io_in[9];
	assign _05337_ = io_in[11] & ~_05336_;
	assign _05338_ = _01568_ | io_in[7];
	assign _05339_ = _05338_ | _01208_;
	assign _05340_ = _05339_ | io_in[10];
	assign _05341_ = io_in[11] & ~_05340_;
	assign _05342_ = _00521_ | _03759_;
	assign _05343_ = _05342_ | io_in[7];
	assign _05344_ = _05343_ | _06310_;
	assign _05346_ = io_in[11] & ~_05344_;
	assign _05347_ = _02852_ | _02096_;
	assign _05348_ = _06310_ & ~_05347_;
	assign _05349_ = _01434_ | io_in[7];
	assign _05350_ = _05349_ | io_in[9];
	assign _05351_ = io_in[10] & ~_05350_;
	assign _05352_ = _00120_ | io_in[6];
	assign _05353_ = _05352_ | io_in[7];
	assign _05354_ = _05353_ | io_in[8];
	assign _05355_ = _05354_ | _02096_;
	assign _05357_ = _05355_ | io_in[10];
	assign _05358_ = io_in[11] & ~_05357_;
	assign _05359_ = _01058_ | io_in[6];
	assign _05360_ = _05359_ | io_in[7];
	assign _05361_ = _05360_ | _01208_;
	assign _05362_ = _05361_ | io_in[9];
	assign _05363_ = _05362_ | io_in[10];
	assign _05364_ = io_in[11] & ~_05363_;
	assign _05365_ = _01046_ | io_in[8];
	assign _05366_ = _05365_ | _02096_;
	assign _05368_ = io_in[10] & ~_05366_;
	assign _05369_ = _02272_ | io_in[8];
	assign _05370_ = _05369_ | _02096_;
	assign _05371_ = _05370_ | io_in[10];
	assign _05372_ = _01985_ & ~_05371_;
	assign _05373_ = _01685_ | io_in[6];
	assign _05374_ = _05373_ | io_in[8];
	assign _05375_ = _05374_ | io_in[9];
	assign _05376_ = io_in[11] & ~_05375_;
	assign _05377_ = _02576_ | io_in[9];
	assign _05379_ = io_in[10] & ~_05377_;
	assign _05380_ = _01607_ | io_in[5];
	assign _05381_ = _05380_ | _02207_;
	assign _05382_ = _05381_ | io_in[9];
	assign _05383_ = _05382_ | io_in[10];
	assign _05384_ = _01985_ & ~_05383_;
	assign _05385_ = _02751_ | _03094_;
	assign _05386_ = io_in[7] & ~_05385_;
	assign _05387_ = _02458_ | _01208_;
	assign _05388_ = _05387_ | _02096_;
	assign _05390_ = _06310_ & ~_05388_;
	assign _05391_ = _07186_ | _02207_;
	assign _05392_ = _05391_ | io_in[9];
	assign _05393_ = _05392_ | io_in[10];
	assign _05394_ = _01985_ & ~_05393_;
	assign _05395_ = _04389_ | io_in[9];
	assign _05396_ = io_in[11] & ~_05395_;
	assign _05397_ = _01321_ | io_in[7];
	assign _05398_ = _05397_ | io_in[8];
	assign _05399_ = _05398_ | _02096_;
	assign _05401_ = io_in[11] & ~_05399_;
	assign _05402_ = _01195_ | _02207_;
	assign _05403_ = _05402_ | io_in[8];
	assign _05404_ = io_in[10] & ~_05403_;
	assign _05405_ = _01220_ | io_in[7];
	assign _05406_ = _05405_ | io_in[8];
	assign _05407_ = _05406_ | io_in[9];
	assign _05408_ = io_in[10] & ~_05407_;
	assign _05409_ = _01578_ | io_in[9];
	assign _05410_ = io_in[11] & ~_05409_;
	assign _05412_ = _04012_ | _01208_;
	assign _05413_ = _06310_ & ~_05412_;
	assign _05414_ = io_in[9] & ~_01004_;
	assign _05415_ = _03590_ | io_in[6];
	assign _05416_ = _05415_ | io_in[8];
	assign _05417_ = _05416_ | io_in[9];
	assign _05418_ = io_in[10] & ~_05417_;
	assign _05419_ = _02860_ | _03759_;
	assign _05420_ = _05419_ | io_in[7];
	assign _05421_ = _05420_ | _01208_;
	assign _05424_ = _05421_ | io_in[9];
	assign _05425_ = _01985_ & ~_05424_;
	assign _05426_ = _01387_ | io_in[8];
	assign _05427_ = _05426_ | _02096_;
	assign _05428_ = io_in[10] & ~_05427_;
	assign _05429_ = _01921_ | _06310_;
	assign _05430_ = io_in[11] & ~_05429_;
	assign _05431_ = _02373_ | io_in[6];
	assign _05432_ = _05431_ | io_in[7];
	assign _05433_ = _05432_ | _02096_;
	assign _05435_ = io_in[11] & ~_05433_;
	assign _05436_ = _05411_ | io_in[6];
	assign _05437_ = _05436_ | io_in[8];
	assign _05438_ = _05437_ | _02096_;
	assign _05439_ = io_in[10] & ~_05438_;
	assign _05440_ = _03641_ | _02207_;
	assign _05441_ = io_in[8] & ~_05440_;
	assign _05442_ = _01720_ | io_in[6];
	assign _05443_ = _05442_ | _02207_;
	assign _05444_ = _05443_ | io_in[8];
	assign _05446_ = _02096_ & ~_05444_;
	assign _05447_ = _00684_ | _03759_;
	assign _05448_ = _05447_ | io_in[7];
	assign _05449_ = _05448_ | io_in[9];
	assign _05450_ = io_in[11] & ~_05449_;
	assign _05451_ = _04978_ | _03759_;
	assign _05452_ = _05451_ | _02207_;
	assign _05453_ = _05452_ | io_in[9];
	assign _05454_ = io_in[11] & ~_05453_;
	assign _05455_ = _05191_ | io_in[9];
	assign _05457_ = io_in[10] & ~_05455_;
	assign _05458_ = _01190_ | io_in[7];
	assign _05459_ = _05458_ | io_in[8];
	assign _05460_ = _05459_ | io_in[9];
	assign _05461_ = _01985_ & ~_05460_;
	assign _05462_ = _03960_ | io_in[9];
	assign _05463_ = io_in[11] & ~_05462_;
	assign _05464_ = _03882_ | io_in[8];
	assign _05465_ = _05464_ | _02096_;
	assign _05466_ = _05465_ | io_in[10];
	assign _05468_ = _01985_ & ~_05466_;
	assign _05469_ = _01828_ | io_in[10];
	assign _05470_ = io_in[11] & ~_05469_;
	assign _05471_ = _01439_ | _02207_;
	assign _05472_ = _05471_ | io_in[9];
	assign _05473_ = io_in[11] & ~_05472_;
	assign _05474_ = _02324_ | io_in[7];
	assign _05475_ = _05474_ | _01208_;
	assign _05476_ = io_in[11] & ~_05475_;
	assign _05477_ = _02786_ | _01208_;
	assign _05479_ = _05477_ | _02096_;
	assign _05480_ = _06310_ & ~_05479_;
	assign _05481_ = io_in[10] & ~_03247_;
	assign _05482_ = _02285_ | io_in[6];
	assign _05483_ = _05482_ | _02207_;
	assign _05484_ = _05483_ | _01208_;
	assign _05485_ = _01985_ & ~_05484_;
	assign _05486_ = _03080_ | _01208_;
	assign _05487_ = _05486_ | io_in[9];
	assign _05488_ = io_in[10] & ~_05487_;
	assign _05490_ = _04398_ | _01208_;
	assign _05491_ = _05490_ | io_in[9];
	assign _05492_ = io_in[11] & ~_05491_;
	assign _05493_ = _00504_ | io_in[6];
	assign _05494_ = _05493_ | _01208_;
	assign _05495_ = _05494_ | io_in[9];
	assign _05496_ = _05495_ | io_in[10];
	assign _05497_ = _01985_ & ~_05496_;
	assign _05498_ = _07250_ | io_in[7];
	assign _05499_ = _05498_ | _01208_;
	assign _05501_ = _05499_ | _02096_;
	assign _05502_ = _05501_ | _06310_;
	assign _05503_ = _01985_ & ~_05502_;
	assign _05504_ = _01438_ | io_in[5];
	assign _05505_ = _05504_ | io_in[6];
	assign _05506_ = _05505_ | io_in[7];
	assign _05507_ = _05506_ | _01208_;
	assign _05508_ = io_in[9] & ~_05507_;
	assign _05509_ = _00636_ | io_in[10];
	assign _05510_ = io_in[11] & ~_05509_;
	assign _05512_ = _00175_ | io_in[7];
	assign _05513_ = _05512_ | _02096_;
	assign _05514_ = _05513_ | io_in[10];
	assign _05515_ = io_in[11] & ~_05514_;
	assign _05516_ = _04993_ | io_in[9];
	assign _05517_ = io_in[10] & ~_05516_;
	assign _05518_ = _02524_ | _02207_;
	assign _05519_ = _06310_ & ~_05518_;
	assign _05520_ = _02642_ | _02096_;
	assign _05521_ = io_in[11] & ~_05520_;
	assign _05523_ = _04912_ | _02096_;
	assign _05524_ = io_in[11] & ~_05523_;
	assign _05525_ = _04226_ | _03759_;
	assign _05526_ = _05525_ | io_in[8];
	assign _05527_ = _05526_ | io_in[9];
	assign _05528_ = _05527_ | io_in[10];
	assign _05529_ = _01985_ & ~_05528_;
	assign _05530_ = _05500_ | _03759_;
	assign _05531_ = _05530_ | io_in[7];
	assign _05532_ = _05531_ | io_in[8];
	assign _05535_ = _05532_ | _02096_;
	assign _05536_ = io_in[10] & ~_05535_;
	assign _05537_ = _01175_ | _02207_;
	assign _05538_ = _05537_ | io_in[8];
	assign _05539_ = _05538_ | io_in[10];
	assign _05540_ = _01985_ & ~_05539_;
	assign _05541_ = _00415_ | io_in[7];
	assign _05542_ = _05541_ | io_in[8];
	assign _05543_ = _05542_ | io_in[9];
	assign _05544_ = io_in[11] & ~_05543_;
	assign _05546_ = _02471_ | io_in[6];
	assign _05547_ = _05546_ | _06310_;
	assign _05548_ = io_in[11] & ~_05547_;
	assign _05549_ = _05493_ | io_in[7];
	assign _05550_ = _05549_ | _06310_;
	assign _05551_ = io_in[11] & ~_05550_;
	assign _05552_ = _00694_ | _03759_;
	assign _05553_ = _05552_ | _02207_;
	assign _05554_ = _05553_ | _01208_;
	assign _05555_ = _05554_ | io_in[9];
	assign _05557_ = io_in[10] & ~_05555_;
	assign _05558_ = _02891_ | io_in[9];
	assign _05559_ = io_in[10] & ~_05558_;
	assign _05560_ = _03977_ | io_in[9];
	assign _05561_ = _05560_ | io_in[10];
	assign _05562_ = _01985_ & ~_05561_;
	assign _05563_ = _00375_ | io_in[9];
	assign _05564_ = io_in[10] & ~_05563_;
	assign _05565_ = _00979_ | _02207_;
	assign _05566_ = _05565_ | _06310_;
	assign _05568_ = io_in[11] & ~_05566_;
	assign _05569_ = _01361_ | _02207_;
	assign _05570_ = _05569_ | _01208_;
	assign _05571_ = io_in[11] & ~_05570_;
	assign _05572_ = _01730_ | _01208_;
	assign _05573_ = _05572_ | _02096_;
	assign _05574_ = _05573_ | _06310_;
	assign _05575_ = _01985_ & ~_05574_;
	assign _05576_ = _01470_ | io_in[7];
	assign _05577_ = _05576_ | _02096_;
	assign _05579_ = _05577_ | _06310_;
	assign _05580_ = _01985_ & ~_05579_;
	assign _05581_ = _02708_ | io_in[8];
	assign _05582_ = _05581_ | io_in[9];
	assign _05583_ = io_in[10] & ~_05582_;
	assign _05584_ = _07031_ | io_in[6];
	assign _05585_ = _05584_ | io_in[7];
	assign _05586_ = _05585_ | io_in[8];
	assign _05587_ = _05586_ | io_in[9];
	assign _05588_ = io_in[11] & ~_05587_;
	assign _05590_ = _01306_ | io_in[7];
	assign _05591_ = _05590_ | _06310_;
	assign _05592_ = io_in[11] & ~_05591_;
	assign _05593_ = _01246_ | _01208_;
	assign _05594_ = _05593_ | io_in[10];
	assign _05595_ = io_in[11] & ~_05594_;
	assign _05596_ = _01404_ | _03094_;
	assign _05597_ = _05596_ | _03759_;
	assign _05598_ = _05597_ | _02096_;
	assign _05599_ = io_in[11] & ~_05598_;
	assign _05601_ = _02505_ | _03759_;
	assign _05602_ = _05601_ | io_in[7];
	assign _05603_ = _05602_ | _01208_;
	assign _05604_ = _05603_ | io_in[9];
	assign _05605_ = io_in[10] & ~_05604_;
	assign _05606_ = _02096_ & ~_02953_;
	assign _05607_ = _01175_ | io_in[8];
	assign _05608_ = _05607_ | _02096_;
	assign _05609_ = _05608_ | io_in[10];
	assign _05610_ = io_in[11] & ~_05609_;
	assign _05612_ = _01059_ | _02207_;
	assign _05613_ = _05612_ | io_in[8];
	assign _05614_ = _05613_ | _02096_;
	assign _05615_ = _05614_ | _06310_;
	assign _05616_ = _01985_ & ~_05615_;
	assign _05617_ = _01360_ | io_in[7];
	assign _05618_ = _05617_ | io_in[8];
	assign _05619_ = _05618_ | _02096_;
	assign _05620_ = io_in[10] & ~_05619_;
	assign _05621_ = _01391_ | _02207_;
	assign _05623_ = _05621_ | _01208_;
	assign _05624_ = _06310_ & ~_05623_;
	assign _05625_ = _03315_ | io_in[8];
	assign _05626_ = _05625_ | _02096_;
	assign _05627_ = _05626_ | io_in[10];
	assign _05628_ = _01985_ & ~_05627_;
	assign _05629_ = _02386_ | _02207_;
	assign _05630_ = _05629_ | io_in[8];
	assign _05631_ = _05630_ | _02096_;
	assign _05632_ = _06310_ & ~_05631_;
	assign _05634_ = _05451_ | io_in[7];
	assign _05635_ = _05634_ | _01208_;
	assign _05636_ = _05635_ | _02096_;
	assign _05637_ = _01985_ & ~_05636_;
	assign _05638_ = _02971_ | io_in[6];
	assign _05639_ = _05638_ | _02207_;
	assign _05640_ = _05639_ | io_in[9];
	assign _05641_ = _05640_ | io_in[10];
	assign _05642_ = _01985_ & ~_05641_;
	assign _05643_ = _01666_ | io_in[7];
	assign _05646_ = _05643_ | _01208_;
	assign _05647_ = _05646_ | _02096_;
	assign _05648_ = _06310_ & ~_05647_;
	assign _05649_ = _07352_ | _02207_;
	assign _05650_ = _05649_ | _01208_;
	assign _05651_ = _05650_ | _02096_;
	assign _05652_ = _05651_ | _06310_;
	assign _05653_ = _01985_ & ~_05652_;
	assign _05654_ = _01650_ | io_in[8];
	assign _05655_ = _05654_ | io_in[9];
	assign _05657_ = io_in[11] & ~_05655_;
	assign _05658_ = _05447_ | io_in[8];
	assign _05659_ = _05658_ | _02096_;
	assign _05660_ = io_in[10] & ~_05659_;
	assign _05661_ = _01042_ | _03094_;
	assign _05662_ = _05661_ | _03759_;
	assign _05663_ = _05662_ | io_in[7];
	assign _05664_ = io_in[11] & ~_05663_;
	assign _05665_ = _02970_ | _02207_;
	assign _05666_ = _05665_ | io_in[8];
	assign _05668_ = _05666_ | io_in[9];
	assign _05669_ = io_in[10] & ~_05668_;
	assign _05670_ = _05755_ | io_in[8];
	assign _05671_ = _05670_ | _02096_;
	assign _05672_ = io_in[10] & ~_05671_;
	assign _05673_ = _01580_ | io_in[8];
	assign _05674_ = io_in[11] & ~_05673_;
	assign _05675_ = _04437_ | _06310_;
	assign _05676_ = io_in[11] & ~_05675_;
	assign _05677_ = _02976_ | io_in[8];
	assign _05679_ = _05677_ | _02096_;
	assign _05680_ = io_in[11] & ~_05679_;
	assign _05681_ = _06310_ & ~_02393_;
	assign _05682_ = _01486_ | io_in[9];
	assign _05683_ = io_in[10] & ~_05682_;
	assign _05684_ = _03127_ | _02207_;
	assign _05685_ = _05684_ | io_in[8];
	assign _05686_ = _05685_ | io_in[9];
	assign _05687_ = io_in[10] & ~_05686_;
	assign _05688_ = _06754_ | io_in[7];
	assign _05690_ = _05688_ | io_in[8];
	assign _05691_ = _05690_ | _02096_;
	assign _05692_ = io_in[11] & ~_05691_;
	assign _05693_ = ~(_05478_ & io_in[9]);
	assign _05694_ = io_in[10] & ~_05693_;
	assign _05695_ = _01534_ | _01208_;
	assign _05696_ = _05695_ | _02096_;
	assign _05697_ = _05696_ | _06310_;
	assign _05698_ = _01985_ & ~_05697_;
	assign _05699_ = _01404_ | _03759_;
	assign _05701_ = _05699_ | io_in[7];
	assign _05702_ = _05701_ | io_in[8];
	assign _05703_ = _05702_ | _02096_;
	assign _05704_ = io_in[10] & ~_05703_;
	assign _05705_ = _01334_ | io_in[5];
	assign _05706_ = _05705_ | _03759_;
	assign _05707_ = _05706_ | _01208_;
	assign _05708_ = _05707_ | _02096_;
	assign _05709_ = _01985_ & ~_05708_;
	assign _05710_ = _05585_ | _01208_;
	assign _05712_ = _05710_ | _02096_;
	assign _05713_ = _06310_ & ~_05712_;
	assign _05714_ = _04289_ | _02096_;
	assign _05715_ = _06310_ & ~_05714_;
	assign _05716_ = _01181_ | _02096_;
	assign _05717_ = _01985_ & ~_05716_;
	assign _05718_ = _00988_ | io_in[7];
	assign _05719_ = _05718_ | _01208_;
	assign _05720_ = _05719_ | io_in[10];
	assign _05721_ = io_in[11] & ~_05720_;
	assign _05723_ = _01251_ | _02096_;
	assign _05724_ = _06310_ & ~_05723_;
	assign _05725_ = _02005_ | io_in[9];
	assign _05726_ = _05725_ | io_in[10];
	assign _05727_ = _01985_ & ~_05726_;
	assign _05728_ = _04058_ | io_in[7];
	assign _05729_ = _05728_ | io_in[8];
	assign _05730_ = _05729_ | io_in[9];
	assign _05731_ = io_in[10] & ~_05730_;
	assign _05732_ = _05278_ | _02207_;
	assign _05734_ = _05732_ | io_in[8];
	assign _05735_ = _05734_ | _02096_;
	assign _05736_ = io_in[11] & ~_05735_;
	assign _05737_ = _02535_ | _02207_;
	assign _05738_ = _05737_ | _06310_;
	assign _05739_ = io_in[11] & ~_05738_;
	assign _05740_ = _05739_ | _05736_;
	assign _05741_ = _05740_ | _05731_;
	assign _05742_ = _05741_ | _05727_;
	assign _05743_ = _05742_ | _05724_;
	assign _05745_ = _05743_ | _05721_;
	assign _05746_ = _05745_ | _05717_;
	assign _05747_ = _05746_ | _05715_;
	assign _05748_ = _05747_ | _05713_;
	assign _05749_ = _05748_ | _05709_;
	assign _05750_ = _05749_ | _05704_;
	assign _05751_ = _05750_ | _05698_;
	assign _05752_ = _05751_ | _05694_;
	assign _05753_ = _05752_ | _05692_;
	assign _05754_ = _05753_ | _05687_;
	assign _05757_ = _05754_ | _05683_;
	assign _05758_ = _05757_ | _05681_;
	assign _05759_ = _05758_ | _05680_;
	assign _05760_ = _05759_ | _05676_;
	assign _05761_ = _05760_ | _05674_;
	assign _05762_ = _05761_ | _05672_;
	assign _05763_ = _05762_ | _05669_;
	assign _05764_ = _05763_ | _05664_;
	assign _05765_ = _05764_ | _05660_;
	assign _05766_ = _05765_ | _05657_;
	assign _05768_ = _05766_ | _05653_;
	assign _05769_ = _05768_ | _05648_;
	assign _05770_ = _05769_ | _05642_;
	assign _05771_ = _05770_ | _05637_;
	assign _05772_ = _05771_ | _05632_;
	assign _05773_ = _05772_ | _05628_;
	assign _05774_ = _05773_ | _05624_;
	assign _05775_ = _05774_ | _05620_;
	assign _05776_ = _05775_ | _05616_;
	assign _05777_ = _05776_ | _05610_;
	assign _05779_ = _05777_ | _05606_;
	assign _05780_ = _05779_ | _05605_;
	assign _05781_ = _05780_ | _07357_;
	assign _05782_ = _05781_ | _05599_;
	assign _05783_ = _05782_ | _05595_;
	assign _05784_ = _05783_ | _05592_;
	assign _05785_ = _05784_ | _05588_;
	assign _05786_ = _05785_ | _05583_;
	assign _05787_ = _05786_ | _05580_;
	assign _05788_ = _05787_ | _05575_;
	assign _05790_ = _05788_ | _05571_;
	assign _05791_ = _05790_ | _05568_;
	assign _05792_ = _05791_ | _05564_;
	assign _05793_ = _05792_ | _03130_;
	assign _05794_ = _05793_ | _05562_;
	assign _05795_ = _05794_ | _05559_;
	assign _05796_ = _05795_ | _03125_;
	assign _05797_ = _05796_ | _01909_;
	assign _05798_ = _05797_ | _05557_;
	assign _05799_ = _05798_ | _05551_;
	assign _05801_ = _05799_ | _05548_;
	assign _05802_ = _05801_ | _05544_;
	assign _05803_ = _05802_ | _05540_;
	assign _05804_ = _05803_ | _05536_;
	assign _05805_ = _05804_ | _05529_;
	assign _05806_ = _05805_ | _05524_;
	assign _05807_ = _05806_ | _05521_;
	assign _05808_ = _05807_ | _05519_;
	assign _05809_ = _05808_ | _05517_;
	assign _05810_ = _05809_ | _05515_;
	assign _05812_ = _05810_ | _05510_;
	assign _05813_ = _05812_ | _05508_;
	assign _05814_ = _05813_ | _05503_;
	assign _05815_ = _05814_ | _05497_;
	assign _05816_ = _05815_ | _05492_;
	assign _05817_ = _05816_ | _05488_;
	assign _05818_ = _05817_ | _05485_;
	assign _05819_ = _05818_ | _05481_;
	assign _05820_ = _05819_ | _05480_;
	assign _05821_ = _05820_ | _05476_;
	assign _05823_ = _05821_ | _05473_;
	assign _05824_ = _05823_ | _05470_;
	assign _05825_ = _05824_ | _05468_;
	assign _05826_ = _05825_ | _05463_;
	assign _05827_ = _05826_ | _05461_;
	assign _05828_ = _05827_ | _05457_;
	assign _05829_ = _05828_ | _05454_;
	assign _05830_ = _05829_ | _05450_;
	assign _05831_ = _05830_ | _05446_;
	assign _05832_ = _05831_ | _05441_;
	assign _05834_ = _05832_ | _05439_;
	assign _05835_ = _05834_ | _05435_;
	assign _05836_ = _05835_ | _05430_;
	assign _05837_ = _05836_ | _05428_;
	assign _05838_ = _05837_ | _05425_;
	assign _05839_ = _05838_ | _05418_;
	assign _05840_ = _05839_ | _05414_;
	assign _05841_ = _05840_ | _05413_;
	assign _05842_ = _05841_ | _05410_;
	assign _05843_ = _05842_ | _05408_;
	assign _05845_ = _05843_ | _05404_;
	assign _05846_ = _05845_ | _05401_;
	assign _05847_ = _05846_ | _05396_;
	assign _05848_ = _05847_ | _05394_;
	assign _05849_ = _05848_ | _05390_;
	assign _05850_ = _05849_ | _05386_;
	assign _05851_ = _05850_ | _05384_;
	assign _05852_ = _05851_ | _05379_;
	assign _05853_ = _05852_ | _05376_;
	assign _05854_ = _05853_ | _05372_;
	assign _05856_ = _05854_ | _05368_;
	assign _05857_ = _05856_ | _05364_;
	assign _05858_ = _05857_ | _05358_;
	assign _05859_ = _05858_ | _05351_;
	assign _05860_ = _05859_ | _05348_;
	assign _05861_ = _05860_ | _05346_;
	assign _05862_ = _05861_ | _05341_;
	assign _05863_ = _05862_ | _05337_;
	assign _05864_ = _05863_ | _05335_;
	assign _05865_ = _05864_ | _05330_;
	assign _05868_ = _05865_ | _05327_;
	assign _05869_ = _05868_ | _05326_;
	assign _05870_ = _05869_ | _05321_;
	assign _05871_ = _05870_ | _05317_;
	assign _05872_ = _05871_ | _05315_;
	assign _05873_ = _05872_ | _05313_;
	assign _05874_ = _05873_ | _05306_;
	assign _05875_ = _05874_ | _05301_;
	assign _05876_ = _05875_ | _05295_;
	assign _05877_ = _05876_ | _05290_;
	assign _05879_ = _05877_ | _05286_;
	assign _05880_ = _05879_ | _02395_;
	assign _05881_ = _05880_ | _05284_;
	assign _05882_ = _05881_ | _05276_;
	assign _05883_ = _05882_ | _05274_;
	assign _05884_ = _05883_ | _05271_;
	assign _05885_ = _05884_ | _05265_;
	assign _05886_ = _05885_ | _05261_;
	assign _05887_ = _05886_ | _05255_;
	assign _05888_ = _05887_ | _05250_;
	assign _05890_ = _05888_ | _05246_;
	assign _05891_ = _05890_ | _05240_;
	assign _05892_ = _05891_ | _05233_;
	assign _05893_ = _05892_ | _05229_;
	assign _05894_ = _05893_ | _05225_;
	assign _05895_ = _05894_ | _05221_;
	assign _05896_ = _05895_ | _05217_;
	assign _05897_ = _05896_ | _05214_;
	assign _05898_ = _05897_ | _05210_;
	assign _05899_ = _05898_ | _05206_;
	assign _05901_ = _05899_ | _05204_;
	assign _05902_ = _05901_ | _05197_;
	assign _05903_ = _05902_ | _05194_;
	assign _05904_ = _05903_ | _05188_;
	assign _05905_ = _05904_ | _05186_;
	assign _05906_ = _05905_ | _05183_;
	assign _05907_ = _05906_ | _05181_;
	assign _05908_ = _05907_ | _05177_;
	assign _05909_ = _05908_ | _05172_;
	assign _05910_ = _05909_ | _05170_;
	assign _05912_ = _05910_ | _05168_;
	assign _05913_ = _05912_ | _05164_;
	assign _05914_ = _05913_ | _05158_;
	assign _05915_ = _05914_ | _05154_;
	assign _05916_ = _05915_ | _05150_;
	assign _05917_ = _05916_ | _05148_;
	assign _05918_ = _05917_ | _05144_;
	assign _05919_ = _05918_ | _05140_;
	assign _05920_ = _05919_ | _05137_;
	assign _05921_ = _05920_ | _05132_;
	assign _05923_ = _05921_ | _05128_;
	assign _05924_ = _05923_ | _05126_;
	assign _05925_ = _05924_ | _05122_;
	assign _05926_ = _05925_ | _05120_;
	assign _05927_ = _05926_ | _05116_;
	assign _05928_ = _05927_ | _05113_;
	assign _05929_ = _05928_ | _05110_;
	assign _05930_ = _05929_ | _05105_;
	assign _05931_ = _05930_ | _05099_;
	assign _05932_ = _05931_ | _05095_;
	assign _05934_ = _05932_ | _05088_;
	assign _05935_ = _05934_ | _05086_;
	assign _05936_ = _05935_ | _05082_;
	assign _05937_ = _05936_ | _05081_;
	assign _05938_ = _05937_ | _05074_;
	assign _05939_ = _05938_ | _05072_;
	assign _05940_ = _05939_ | _05070_;
	assign _05941_ = _05940_ | _05065_;
	assign _05942_ = _05941_ | _05062_;
	assign _05943_ = _05942_ | _05059_;
	assign _05945_ = _05943_ | _01394_;
	assign _05946_ = _05945_ | _05055_;
	assign _05947_ = _05946_ | _05051_;
	assign _05948_ = _05947_ | _05048_;
	assign _05949_ = _05948_ | _05046_;
	assign _05950_ = _05949_ | _05041_;
	assign _05951_ = _05950_ | _02384_;
	assign _05952_ = _05951_ | _05037_;
	assign _05953_ = _05952_ | _05030_;
	assign _05954_ = _05953_ | _05026_;
	assign _05956_ = _05954_ | _05021_;
	assign _05957_ = _05956_ | _05018_;
	assign _05958_ = _05957_ | _05017_;
	assign _05959_ = _05958_ | _05014_;
	assign _05960_ = _05959_ | _05010_;
	assign _05961_ = _05960_ | _03739_;
	assign _05962_ = _05961_ | _05007_;
	assign _05963_ = _05962_ | _05002_;
	assign _05964_ = _05963_ | _05000_;
	assign _05965_ = _05964_ | _04999_;
	assign _05967_ = _05965_ | _04995_;
	assign _05968_ = _05967_ | _04991_;
	assign _05969_ = _05968_ | _04985_;
	assign _05970_ = _05969_ | _04983_;
	assign _05971_ = _05970_ | _04982_;
	assign _05972_ = _05971_ | _04976_;
	assign _05973_ = _05972_ | _04972_;
	assign _05974_ = _05973_ | _04969_;
	assign _05975_ = _05974_ | _04964_;
	assign _05976_ = _05975_ | _04960_;
	assign _05979_ = _05976_ | _04955_;
	assign _05980_ = _05979_ | _04951_;
	assign _05981_ = _05980_ | _04948_;
	assign _05982_ = _05981_ | _04944_;
	assign _05983_ = _05982_ | _04940_;
	assign _05984_ = _05983_ | _04939_;
	assign _05985_ = _05984_ | _04936_;
	assign _05986_ = _05985_ | _04935_;
	assign _05987_ = _05986_ | _04928_;
	assign _05988_ = _05987_ | _04926_;
	assign _05990_ = _05988_ | _04924_;
	assign _05991_ = _05990_ | _03644_;
	assign _05992_ = _05991_ | _02843_;
	assign _05993_ = _05992_ | _04920_;
	assign _05994_ = _05993_ | _04917_;
	assign _05995_ = _05994_ | _04913_;
	assign _05996_ = _05995_ | _04907_;
	assign _05997_ = _05996_ | _04902_;
	assign _05998_ = _05997_ | _04898_;
	assign _05999_ = _05998_ | _04895_;
	assign _06001_ = _05999_ | _04893_;
	assign _06002_ = _06001_ | _04888_;
	assign _06003_ = _06002_ | _04883_;
	assign _06004_ = _06003_ | _04880_;
	assign _06005_ = _06004_ | _04878_;
	assign _06006_ = _06005_ | _04874_;
	assign _06007_ = _06006_ | _04872_;
	assign _06008_ = _06007_ | _04864_;
	assign _06009_ = _06008_ | _04862_;
	assign _06010_ = _06009_ | _04859_;
	assign _06012_ = _06010_ | _04857_;
	assign _06013_ = _06012_ | _04853_;
	assign _06014_ = _06013_ | _04849_;
	assign _06015_ = _06014_ | _04843_;
	assign _06016_ = _06015_ | _04840_;
	assign _06017_ = _06016_ | _04837_;
	assign _06018_ = _06017_ | _04835_;
	assign _06019_ = _06018_ | _04829_;
	assign _06020_ = _06019_ | _04825_;
	assign _06021_ = _06020_ | _04821_;
	assign \mchip.val [1] = _06021_ | _04816_;
	assign _06023_ = _04524_ | io_in[6];
	assign _06024_ = _06023_ | _02207_;
	assign _06025_ = _06024_ | io_in[8];
	assign _06026_ = io_in[11] & ~_06025_;
	assign _06027_ = io_in[11] & ~_03014_;
	assign _06028_ = io_in[7] & ~_03830_;
	assign _06029_ = _06509_ | io_in[6];
	assign _06030_ = _06029_ | io_in[8];
	assign _06031_ = _06030_ | _02096_;
	assign _06033_ = _06031_ | io_in[10];
	assign _06034_ = _01985_ & ~_06033_;
	assign _06035_ = _00585_ | _03759_;
	assign _06036_ = _06035_ | _02207_;
	assign _06037_ = _06036_ | _06310_;
	assign _06038_ = io_in[11] & ~_06037_;
	assign _06039_ = _02618_ | _02207_;
	assign _06040_ = _06039_ | _01208_;
	assign _06041_ = _06040_ | io_in[9];
	assign _06042_ = io_in[10] & ~_06041_;
	assign _06044_ = _01931_ | _02096_;
	assign _06045_ = _06310_ & ~_06044_;
	assign _06046_ = _01360_ | _01208_;
	assign _06047_ = _06046_ | io_in[9];
	assign _06048_ = io_in[10] & ~_06047_;
	assign _06049_ = _01277_ | io_in[7];
	assign _06050_ = _06049_ | io_in[9];
	assign _06051_ = _06310_ & ~_06050_;
	assign _06052_ = _02296_ | _02096_;
	assign _06053_ = _06052_ | _06310_;
	assign _06055_ = _01985_ & ~_06053_;
	assign _06056_ = _05075_ | io_in[6];
	assign _06057_ = _01208_ & ~_06056_;
	assign _06058_ = _03197_ | _01208_;
	assign _06059_ = _02096_ & ~_06058_;
	assign _06060_ = _02012_ | _02207_;
	assign _06061_ = _06060_ | io_in[9];
	assign _06062_ = _06061_ | _06310_;
	assign _06063_ = _01985_ & ~_06062_;
	assign _06064_ = _01507_ | io_in[7];
	assign _06066_ = _06064_ | io_in[8];
	assign _06067_ = io_in[10] & ~_06066_;
	assign _06068_ = _02771_ | io_in[8];
	assign _06069_ = io_in[11] & ~_06068_;
	assign _06070_ = _01990_ | io_in[6];
	assign _06071_ = _06070_ | _02207_;
	assign _06072_ = _06071_ | _02096_;
	assign _06073_ = _01985_ & ~_06072_;
	assign _06074_ = _01006_ | io_in[5];
	assign _06075_ = _06074_ | io_in[6];
	assign _06077_ = _06075_ | _02207_;
	assign _06078_ = _06077_ | io_in[9];
	assign _06079_ = io_in[10] & ~_06078_;
	assign _06080_ = _05003_ | io_in[9];
	assign _06081_ = _06080_ | io_in[10];
	assign _06082_ = io_in[11] & ~_06081_;
	assign _06083_ = _01485_ | io_in[6];
	assign _06084_ = _06083_ | io_in[7];
	assign _06085_ = _06084_ | _01208_;
	assign _06086_ = _06085_ | _02096_;
	assign _06089_ = _06086_ | _06310_;
	assign _06090_ = _01985_ & ~_06089_;
	assign _06091_ = _01225_ | io_in[8];
	assign _06092_ = _06091_ | io_in[10];
	assign _06093_ = _01985_ & ~_06092_;
	assign _06094_ = _02096_ & ~_02552_;
	assign _06095_ = _01919_ | _02207_;
	assign _06096_ = _06095_ | _06310_;
	assign _06097_ = io_in[11] & ~_06096_;
	assign _06098_ = _03887_ | _02096_;
	assign _06100_ = io_in[11] & ~_06098_;
	assign _06101_ = _04978_ | _01208_;
	assign _06102_ = _06101_ | io_in[9];
	assign _06103_ = _01985_ & ~_06102_;
	assign _06104_ = _05411_ | _03094_;
	assign _06105_ = _06104_ | _03759_;
	assign _06106_ = io_in[11] & ~_06105_;
	assign _06107_ = _01547_ | _01208_;
	assign _06108_ = _06107_ | io_in[9];
	assign _06109_ = io_in[10] & ~_06108_;
	assign _06111_ = _04513_ | _03759_;
	assign _06112_ = _06111_ | _02207_;
	assign _06113_ = _06112_ | io_in[9];
	assign _06114_ = io_in[11] & ~_06113_;
	assign _06115_ = _00768_ | io_in[5];
	assign _06116_ = _06115_ | io_in[6];
	assign _06117_ = _06116_ | _02207_;
	assign _06118_ = _06117_ | _02096_;
	assign _06119_ = io_in[10] & ~_06118_;
	assign _06120_ = _07075_ | io_in[5];
	assign _06122_ = _06120_ | _03759_;
	assign _06123_ = _06122_ | _06310_;
	assign _06124_ = io_in[11] & ~_06123_;
	assign _06125_ = _07257_ | _03759_;
	assign _06126_ = _06125_ | io_in[7];
	assign _06127_ = _06126_ | io_in[8];
	assign _06128_ = io_in[10] & ~_06127_;
	assign _06129_ = _02018_ | _03759_;
	assign _06130_ = _06129_ | io_in[7];
	assign _06131_ = _06130_ | _01208_;
	assign _06133_ = _06131_ | _02096_;
	assign _06134_ = _06133_ | _06310_;
	assign _06135_ = io_in[11] & ~_06134_;
	assign _06136_ = _02756_ | io_in[9];
	assign _06137_ = _06310_ & ~_06136_;
	assign _06138_ = _00660_ | io_in[6];
	assign _06139_ = _06138_ | io_in[7];
	assign _06140_ = _06139_ | _01208_;
	assign _06141_ = _06140_ | io_in[9];
	assign _06142_ = io_in[11] & ~_06141_;
	assign _06144_ = _00743_ | _03759_;
	assign _06145_ = _06144_ | _02207_;
	assign _06146_ = _06145_ | _01208_;
	assign _06147_ = _06146_ | _02096_;
	assign _06148_ = _06147_ | _06310_;
	assign _06149_ = _01985_ & ~_06148_;
	assign _06150_ = _00773_ | _03759_;
	assign _06151_ = _06150_ | io_in[7];
	assign _06152_ = _06151_ | io_in[8];
	assign _06153_ = _06152_ | io_in[9];
	assign _06155_ = io_in[11] & ~_06153_;
	assign _06156_ = _07265_ | io_in[8];
	assign _06157_ = _06156_ | io_in[10];
	assign _06158_ = _01985_ & ~_06157_;
	assign _06159_ = _06310_ & ~_00460_;
	assign _06160_ = _05482_ | _02096_;
	assign _06161_ = _06310_ & ~_06160_;
	assign _06162_ = _02417_ | _01208_;
	assign _06163_ = _01985_ & ~_06162_;
	assign _06164_ = _06853_ | io_in[8];
	assign _06166_ = _06164_ | _02096_;
	assign _06167_ = _06166_ | io_in[10];
	assign _06168_ = _01985_ & ~_06167_;
	assign _06169_ = io_in[8] & ~_01581_;
	assign _06170_ = _01006_ | _03759_;
	assign _06171_ = _06170_ | io_in[7];
	assign _06172_ = _06171_ | io_in[9];
	assign _06173_ = io_in[11] & ~_06172_;
	assign _06174_ = _02725_ | io_in[8];
	assign _06175_ = io_in[11] & ~_06174_;
	assign _06177_ = _04826_ | io_in[9];
	assign _06178_ = io_in[10] & ~_06177_;
	assign _06179_ = _03725_ | io_in[7];
	assign _06180_ = _06179_ | io_in[8];
	assign _06181_ = _06180_ | io_in[10];
	assign _06182_ = _01985_ & ~_06181_;
	assign _06183_ = _01360_ | io_in[8];
	assign _06184_ = _06183_ | _02096_;
	assign _06185_ = io_in[11] & ~_06184_;
	assign _06186_ = io_in[10] & ~_05597_;
	assign _06188_ = _02000_ | _02207_;
	assign _06189_ = _06188_ | _01208_;
	assign _06190_ = _01985_ & ~_06189_;
	assign _06191_ = _01157_ | io_in[7];
	assign _06192_ = io_in[11] & ~_06191_;
	assign _06193_ = _00812_ | io_in[5];
	assign _06194_ = _06193_ | io_in[6];
	assign _06195_ = _06194_ | _02207_;
	assign _06196_ = _06195_ | io_in[8];
	assign _06197_ = _06196_ | io_in[9];
	assign _06200_ = io_in[10] & ~_06197_;
	assign _06201_ = _02096_ & ~_02412_;
	assign _06202_ = _05129_ | io_in[7];
	assign _06203_ = _06202_ | _01208_;
	assign _06204_ = _02096_ & ~_06203_;
	assign _06205_ = _01818_ | _02207_;
	assign _06206_ = _06205_ | _02096_;
	assign _06207_ = _06206_ | io_in[10];
	assign _06208_ = io_in[11] & ~_06207_;
	assign _06209_ = _01184_ | _01208_;
	assign _06211_ = _06209_ | _02096_;
	assign _06212_ = _06310_ & ~_06211_;
	assign _06213_ = _05359_ | _01208_;
	assign _06214_ = _06213_ | _02096_;
	assign _06215_ = _06214_ | _06310_;
	assign _06216_ = io_in[11] & ~_06215_;
	assign _06217_ = _04325_ | _02096_;
	assign _06218_ = _06310_ & ~_06217_;
	assign _06219_ = _03728_ | _06310_;
	assign _06220_ = io_in[11] & ~_06219_;
	assign _06222_ = _01746_ | _01208_;
	assign _06223_ = io_in[9] & ~_06222_;
	assign _06224_ = _01985_ & ~_01508_;
	assign _06225_ = _02720_ | io_in[8];
	assign _06226_ = _06225_ | io_in[9];
	assign _06227_ = io_in[10] & ~_06226_;
	assign _06228_ = _01386_ | io_in[8];
	assign _06229_ = io_in[10] & ~_06228_;
	assign _06230_ = _01790_ | _02096_;
	assign _06231_ = _06230_ | io_in[10];
	assign _06233_ = _01985_ & ~_06231_;
	assign _06234_ = _01725_ | _06310_;
	assign _06235_ = io_in[11] & ~_06234_;
	assign _06236_ = _00900_ | io_in[7];
	assign _06237_ = _06236_ | _01208_;
	assign _06238_ = _06237_ | _06310_;
	assign _06239_ = _01985_ & ~_06238_;
	assign _06240_ = _01985_ & ~_02481_;
	assign _06241_ = _07430_ & ~_06310_;
	assign _06242_ = _01745_ | io_in[7];
	assign _06244_ = _06242_ | _02096_;
	assign _06245_ = _01985_ & ~_06244_;
	assign _06246_ = _00724_ | io_in[7];
	assign _06247_ = _06246_ | _02096_;
	assign _06248_ = _01985_ & ~_06247_;
	assign _06249_ = _02694_ | _06310_;
	assign _06250_ = io_in[11] & ~_06249_;
	assign _06251_ = _01985_ & ~_03222_;
	assign _06252_ = _03936_ | _02207_;
	assign _06253_ = _06252_ | io_in[8];
	assign _06255_ = io_in[10] & ~_06253_;
	assign _06256_ = _04509_ | io_in[9];
	assign _06257_ = _06256_ | io_in[10];
	assign _06258_ = _01985_ & ~_06257_;
	assign _06259_ = _06509_ | _03759_;
	assign _06260_ = _06259_ | _02207_;
	assign _06261_ = _06260_ | _01208_;
	assign _06262_ = _06261_ | io_in[9];
	assign _06263_ = io_in[10] & ~_06262_;
	assign _06264_ = _00632_ | _01208_;
	assign _06266_ = _06264_ | io_in[9];
	assign _06267_ = io_in[11] & ~_06266_;
	assign _06268_ = _03662_ | _01208_;
	assign _06269_ = _06268_ | _02096_;
	assign _06270_ = _06269_ | _06310_;
	assign _06271_ = _01985_ & ~_06270_;
	assign _06272_ = _04472_ | _02096_;
	assign _06273_ = _06310_ & ~_06272_;
	assign _06274_ = _04204_ | _02207_;
	assign _06275_ = _06274_ | io_in[8];
	assign _06277_ = _02096_ & ~_06275_;
	assign _06278_ = _04919_ | _06310_;
	assign _06279_ = _01985_ & ~_06278_;
	assign _06280_ = _01111_ | _01208_;
	assign _06281_ = _06280_ | io_in[9];
	assign _06282_ = io_in[11] & ~_06281_;
	assign _06283_ = _04428_ | _02096_;
	assign _06284_ = io_in[11] & ~_06283_;
	assign _06285_ = _03842_ | _03759_;
	assign _06286_ = _02096_ & ~_06285_;
	assign _06288_ = _05420_ | io_in[8];
	assign _06289_ = io_in[9] & ~_06288_;
	assign _06290_ = _00043_ | _07422_;
	assign _06291_ = _06290_ | io_in[6];
	assign _06292_ = _06291_ | io_in[7];
	assign _06293_ = _06292_ | io_in[8];
	assign _06294_ = _06293_ | _02096_;
	assign _06295_ = io_in[10] & ~_06294_;
	assign _06296_ = _03871_ | _02207_;
	assign _06297_ = _06296_ | io_in[8];
	assign _06299_ = _06297_ | _02096_;
	assign _06300_ = io_in[10] & ~_06299_;
	assign _06301_ = _00687_ | _03094_;
	assign _06302_ = _03759_ & ~_06301_;
	assign _06303_ = _01745_ | _01208_;
	assign _06304_ = _06303_ | io_in[10];
	assign _06305_ = _01985_ & ~_06304_;
	assign _06306_ = _03151_ | io_in[8];
	assign _06307_ = io_in[10] & ~_06306_;
	assign _06308_ = _00327_ & ~io_in[11];
	assign _06311_ = _07255_ | io_in[6];
	assign _06312_ = _06311_ | io_in[7];
	assign _06313_ = _01208_ & ~_06312_;
	assign _06314_ = _02727_ | _03759_;
	assign _06315_ = _06314_ | _02207_;
	assign _06316_ = _06315_ | io_in[8];
	assign _06317_ = _06316_ | io_in[9];
	assign _06318_ = io_in[11] & ~_06317_;
	assign _06319_ = _00439_ | _03094_;
	assign _06320_ = _06319_ | io_in[6];
	assign _06322_ = _06320_ | _06310_;
	assign _06323_ = io_in[11] & ~_06322_;
	assign _06324_ = _01306_ | _02207_;
	assign _06325_ = _06324_ | _01208_;
	assign _06326_ = _06325_ | _06310_;
	assign _06327_ = _01985_ & ~_06326_;
	assign _06328_ = _00998_ | _01208_;
	assign _06329_ = _06328_ | io_in[9];
	assign _06330_ = io_in[10] & ~_06329_;
	assign _06331_ = _02551_ | io_in[8];
	assign _06333_ = _06331_ | _02096_;
	assign _06334_ = io_in[10] & ~_06333_;
	assign _06335_ = _02381_ | io_in[9];
	assign _06336_ = _06310_ & ~_06335_;
	assign _06337_ = _00933_ | io_in[6];
	assign _06338_ = _06337_ | _02207_;
	assign _06339_ = _06338_ | _01208_;
	assign _06340_ = _06339_ | _02096_;
	assign _06341_ = _06340_ | _06310_;
	assign _06342_ = _01985_ & ~_06341_;
	assign _06344_ = _00245_ | io_in[7];
	assign _06345_ = _06344_ | _01208_;
	assign _06346_ = _06345_ | _02096_;
	assign _06347_ = _06346_ | io_in[10];
	assign _06348_ = _01985_ & ~_06347_;
	assign _06349_ = _04446_ | io_in[9];
	assign _06350_ = _06310_ & ~_06349_;
	assign _06351_ = io_in[1] | ~io_in[4];
	assign _06352_ = _06351_ | _03759_;
	assign _06353_ = _06352_ | _01208_;
	assign _06355_ = _06353_ | io_in[9];
	assign _06356_ = _06355_ | io_in[10];
	assign _06357_ = _01985_ & ~_06356_;
	assign _06358_ = _04268_ | _03094_;
	assign _06359_ = _06358_ | _03759_;
	assign _06360_ = _06359_ | io_in[7];
	assign _06361_ = io_in[10] & ~_06360_;
	assign _06362_ = _01522_ | io_in[9];
	assign _06363_ = io_in[11] & ~_06362_;
	assign _06364_ = _00625_ | io_in[8];
	assign _06366_ = _06364_ | _02096_;
	assign _06367_ = _06310_ & ~_06366_;
	assign _06368_ = _00649_ | _01208_;
	assign _06369_ = _06368_ | _02096_;
	assign _06370_ = _06310_ & ~_06369_;
	assign _06371_ = _02808_ | _01208_;
	assign _06372_ = _06371_ | io_in[10];
	assign _06373_ = io_in[11] & ~_06372_;
	assign _06374_ = _04362_ | io_in[8];
	assign _06375_ = io_in[11] & ~_06374_;
	assign _06377_ = _04362_ | io_in[7];
	assign _06378_ = _02096_ & ~_06377_;
	assign _06379_ = _01809_ | _01208_;
	assign _06380_ = _06379_ | _02096_;
	assign _06381_ = _06380_ | _06310_;
	assign _06382_ = _01985_ & ~_06381_;
	assign _06383_ = _02096_ & ~_01619_;
	assign _06384_ = _06310_ & ~_03649_;
	assign _06385_ = _01105_ | io_in[7];
	assign _06386_ = _06385_ | _06310_;
	assign _06388_ = io_in[11] & ~_06386_;
	assign _06389_ = _01839_ | io_in[8];
	assign _06390_ = io_in[11] & ~_06389_;
	assign _06391_ = _01914_ | _01208_;
	assign _06392_ = _06391_ | io_in[9];
	assign _06393_ = io_in[10] & ~_06392_;
	assign _06394_ = _04973_ | io_in[8];
	assign _06395_ = _06394_ | _02096_;
	assign _06396_ = io_in[10] & ~_06395_;
	assign _06397_ = _03592_ | io_in[6];
	assign _06399_ = _06397_ | io_in[8];
	assign _06400_ = _06399_ | _02096_;
	assign _06401_ = _06400_ | io_in[10];
	assign _06402_ = _01985_ & ~_06401_;
	assign _06403_ = _07271_ | io_in[7];
	assign _06404_ = _06403_ | io_in[8];
	assign _06405_ = _06404_ | io_in[9];
	assign _06406_ = io_in[10] & ~_06405_;
	assign _06407_ = _01406_ | _01208_;
	assign _06408_ = _01985_ & ~_06407_;
	assign _06410_ = _01601_ | io_in[8];
	assign _06411_ = _06410_ | io_in[9];
	assign _06412_ = io_in[11] & ~_06411_;
	assign _06413_ = _07257_ | io_in[7];
	assign _06414_ = _06413_ | io_in[8];
	assign _06415_ = _06414_ | io_in[9];
	assign _06416_ = io_in[11] & ~_06415_;
	assign _06417_ = _01501_ | _01208_;
	assign _06418_ = _06417_ | _02096_;
	assign _06419_ = _06310_ & ~_06418_;
	assign _06422_ = _02669_ | io_in[8];
	assign _06423_ = _06422_ | io_in[9];
	assign _06424_ = _01985_ & ~_06423_;
	assign _06425_ = _01277_ | _03759_;
	assign _06426_ = _06425_ | _01208_;
	assign _06427_ = _06426_ | _06310_;
	assign _06428_ = _01985_ & ~_06427_;
	assign _06429_ = _04326_ | _03759_;
	assign _06430_ = _06429_ | _02096_;
	assign _06431_ = _06430_ | io_in[10];
	assign _06433_ = _01985_ & ~_06431_;
	assign _06434_ = _03590_ | _03759_;
	assign _06435_ = _06434_ | _02207_;
	assign _06436_ = _06435_ | _06310_;
	assign _06437_ = _01985_ & ~_06436_;
	assign _06438_ = _02593_ | _02096_;
	assign _06439_ = _06310_ & ~_06438_;
	assign _06440_ = _01101_ | io_in[8];
	assign _06441_ = io_in[11] & ~_06440_;
	assign _06442_ = _01214_ | io_in[7];
	assign _06444_ = _06442_ | io_in[8];
	assign _06445_ = _01985_ & ~_06444_;
	assign _06446_ = _02344_ | io_in[8];
	assign _06447_ = _06446_ | _02096_;
	assign _06448_ = io_in[10] & ~_06447_;
	assign _06449_ = _02770_ | io_in[8];
	assign _06450_ = _06449_ | io_in[10];
	assign _06451_ = _01985_ & ~_06450_;
	assign _06452_ = _00227_ | io_in[7];
	assign _06453_ = _06452_ | io_in[8];
	assign _06455_ = _06453_ | io_in[9];
	assign _06456_ = io_in[10] & ~_06455_;
	assign _06457_ = _03304_ | _03094_;
	assign _06458_ = _06457_ | io_in[8];
	assign _06459_ = io_in[9] & ~_06458_;
	assign _06460_ = _01367_ | _01208_;
	assign _06461_ = _06460_ | _06310_;
	assign _06462_ = _01985_ & ~_06461_;
	assign _06463_ = _03887_ | _02207_;
	assign _06464_ = _06463_ | io_in[8];
	assign _06466_ = _02096_ & ~_06464_;
	assign _06467_ = _07257_ | _01208_;
	assign _06468_ = _06467_ | io_in[9];
	assign _06469_ = _06468_ | io_in[10];
	assign _06470_ = _01985_ & ~_06469_;
	assign _06471_ = _07153_ | _02207_;
	assign _06472_ = _06471_ | _02096_;
	assign _06473_ = _06310_ & ~_06472_;
	assign _06474_ = _04841_ | _01208_;
	assign _06475_ = io_in[9] & ~_06474_;
	assign _06477_ = _03002_ | _01208_;
	assign _06478_ = _06477_ | io_in[9];
	assign _06479_ = _01985_ & ~_06478_;
	assign _06480_ = _05705_ | _02207_;
	assign _06481_ = _06480_ | io_in[8];
	assign _06482_ = io_in[10] & ~_06481_;
	assign _06483_ = _05160_ | io_in[7];
	assign _06484_ = _06483_ | _02096_;
	assign _06485_ = _06484_ | _06310_;
	assign _06486_ = _01985_ & ~_06485_;
	assign _06488_ = _06290_ | _03759_;
	assign _06489_ = _06488_ | io_in[7];
	assign _06490_ = _06489_ | io_in[8];
	assign _06491_ = _06490_ | io_in[9];
	assign _06492_ = io_in[10] & ~_06491_;
	assign _06493_ = _01880_ | _02096_;
	assign _06494_ = _06310_ & ~_06493_;
	assign _06495_ = _03897_ | _02207_;
	assign _06496_ = _06495_ | _01208_;
	assign _06497_ = _02096_ & ~_06496_;
	assign _06499_ = _00010_ | _02207_;
	assign _06500_ = _06499_ | io_in[8];
	assign _06501_ = _06500_ | io_in[9];
	assign _06502_ = io_in[10] & ~_06501_;
	assign _06503_ = _07250_ | io_in[6];
	assign _06504_ = _06503_ | _02207_;
	assign _06505_ = _06504_ | _01208_;
	assign _06506_ = _02096_ & ~_06505_;
	assign _06507_ = _05789_ | _02207_;
	assign _06508_ = _06507_ | _01208_;
	assign _06510_ = _06508_ | io_in[10];
	assign _06511_ = io_in[11] & ~_06510_;
	assign _06512_ = _00250_ | io_in[5];
	assign _06513_ = _06512_ | _02207_;
	assign _06514_ = _06513_ | _06310_;
	assign _06515_ = io_in[11] & ~_06514_;
	assign _06516_ = _01698_ | _03094_;
	assign _06517_ = _06516_ | io_in[6];
	assign _06518_ = _06517_ | io_in[7];
	assign _06519_ = _06518_ | _06310_;
	assign _06521_ = io_in[11] & ~_06519_;
	assign _06522_ = _03757_ | io_in[7];
	assign _06523_ = _06522_ | io_in[8];
	assign _06524_ = _06523_ | io_in[9];
	assign _06525_ = io_in[10] & ~_06524_;
	assign _06526_ = _03696_ | _02207_;
	assign _06527_ = _06526_ | io_in[10];
	assign _06528_ = _01985_ & ~_06527_;
	assign _06529_ = _00988_ | io_in[9];
	assign _06530_ = _01985_ & ~_06529_;
	assign _06533_ = _02602_ | io_in[8];
	assign _06534_ = io_in[9] & ~_06533_;
	assign _06535_ = _00274_ | _03094_;
	assign _06536_ = _06535_ | io_in[7];
	assign _06537_ = _06536_ | _01208_;
	assign _06538_ = io_in[11] & ~_06537_;
	assign _06539_ = _01671_ | _02207_;
	assign _06540_ = _06539_ | io_in[8];
	assign _06541_ = _06540_ | io_in[9];
	assign _06542_ = io_in[10] & ~_06541_;
	assign _06544_ = _00239_ | io_in[7];
	assign _06545_ = _06544_ | _01208_;
	assign _06546_ = _06545_ | io_in[9];
	assign _06547_ = io_in[10] & ~_06546_;
	assign _06548_ = _00500_ | io_in[8];
	assign _06549_ = _06548_ | _02096_;
	assign _06550_ = _06549_ | io_in[10];
	assign _06551_ = _01985_ & ~_06550_;
	assign _06552_ = _01404_ | io_in[6];
	assign _06553_ = _06552_ | _02207_;
	assign _06555_ = _06553_ | _02096_;
	assign _06556_ = _06310_ & ~_06555_;
	assign _06557_ = io_in[10] & ~_04276_;
	assign _06558_ = _01985_ & ~_05361_;
	assign _06559_ = _05533_ | io_in[10];
	assign _06560_ = _01985_ & ~_06559_;
	assign _06561_ = _00178_ | _03759_;
	assign _06562_ = _06561_ | io_in[7];
	assign _06563_ = _06562_ | _01208_;
	assign _06564_ = _06563_ | _06310_;
	assign _06566_ = _01985_ & ~_06564_;
	assign _06567_ = _04431_ | _02207_;
	assign _06568_ = _06567_ | io_in[10];
	assign _06569_ = io_in[11] & ~_06568_;
	assign _06570_ = _05613_ | io_in[10];
	assign _06571_ = io_in[11] & ~_06570_;
	assign _06572_ = _02407_ | io_in[7];
	assign _06573_ = _06572_ | io_in[8];
	assign _06574_ = _06573_ | _02096_;
	assign _06575_ = io_in[10] & ~_06574_;
	assign _06577_ = _02018_ | io_in[6];
	assign _06578_ = _06577_ | io_in[7];
	assign _06579_ = _06578_ | _01208_;
	assign _06580_ = _06579_ | _02096_;
	assign _06581_ = _01985_ & ~_06580_;
	assign _06582_ = _03713_ | _01208_;
	assign _06583_ = _06582_ | io_in[9];
	assign _06584_ = _06583_ | io_in[10];
	assign _06585_ = _01985_ & ~_06584_;
	assign _06586_ = _00889_ | _03759_;
	assign _06588_ = _06586_ | _02207_;
	assign _06589_ = _06588_ | io_in[9];
	assign _06590_ = io_in[10] & ~_06589_;
	assign _06591_ = _04836_ | _06310_;
	assign _06592_ = _01985_ & ~_06591_;
	assign _06593_ = _01134_ | io_in[8];
	assign _06594_ = io_in[9] & ~_06593_;
	assign _06595_ = _00768_ | _01208_;
	assign _06596_ = _06595_ | io_in[9];
	assign _06597_ = _06596_ | io_in[10];
	assign _06599_ = _01985_ & ~_06597_;
	assign _06600_ = _05173_ | io_in[7];
	assign _06601_ = _06600_ | io_in[8];
	assign _06602_ = io_in[9] & ~_06601_;
	assign _06603_ = _01794_ | _02207_;
	assign _06604_ = io_in[10] & ~_06603_;
	assign _06605_ = _05042_ | io_in[7];
	assign _06606_ = _06605_ | io_in[8];
	assign _06607_ = _06606_ | io_in[9];
	assign _06608_ = io_in[11] & ~_06607_;
	assign _06610_ = _06243_ | _03094_;
	assign _06611_ = _02207_ & ~_06610_;
	assign _06612_ = _00496_ | io_in[6];
	assign _06613_ = _06612_ | _06310_;
	assign _06614_ = io_in[11] & ~_06613_;
	assign _06615_ = _02635_ | io_in[6];
	assign _06616_ = _02207_ & ~_06615_;
	assign _06617_ = _01657_ | _02207_;
	assign _06618_ = _06617_ | io_in[8];
	assign _06619_ = _06618_ | io_in[9];
	assign _06621_ = _06619_ | _06310_;
	assign _06622_ = _01985_ & ~_06621_;
	assign _06623_ = _01208_ & ~_06191_;
	assign _06624_ = _07142_ | io_in[5];
	assign _06625_ = _06624_ | io_in[6];
	assign _06626_ = _06625_ | io_in[7];
	assign _06627_ = _06626_ | _06310_;
	assign _06628_ = io_in[11] & ~_06627_;
	assign _06629_ = _05436_ | io_in[9];
	assign _06630_ = _06629_ | io_in[10];
	assign _06632_ = _01985_ & ~_06630_;
	assign _06633_ = _00547_ | _03759_;
	assign _06634_ = _06633_ | _02207_;
	assign _06635_ = _06634_ | io_in[8];
	assign _06636_ = _06635_ | _02096_;
	assign _06637_ = io_in[10] & ~_06636_;
	assign _06638_ = _06310_ & ~_04510_;
	assign _06639_ = _01431_ | io_in[9];
	assign _06640_ = io_in[10] & ~_06639_;
	assign _06641_ = _04901_ | io_in[8];
	assign _06644_ = _06641_ | _02096_;
	assign _06645_ = io_in[10] & ~_06644_;
	assign _06646_ = _06368_ | io_in[9];
	assign _06647_ = io_in[10] & ~_06646_;
	assign _06648_ = _07455_ | io_in[6];
	assign _06649_ = _06648_ | _02207_;
	assign _06650_ = _06649_ | _01208_;
	assign _06651_ = io_in[11] & ~_06650_;
	assign _06652_ = _06310_ & ~_05695_;
	assign _06653_ = _01736_ | io_in[7];
	assign _06655_ = _06653_ | io_in[8];
	assign _06656_ = io_in[10] & ~_06655_;
	assign _06657_ = _01985_ & ~_05136_;
	assign _06658_ = _03909_ | _02096_;
	assign _06659_ = io_in[11] & ~_06658_;
	assign _06660_ = _01214_ | _02207_;
	assign _06661_ = _06660_ | _01208_;
	assign _06662_ = io_in[10] & ~_06661_;
	assign _06663_ = _01637_ | _01208_;
	assign _06664_ = _06663_ | _02096_;
	assign _06666_ = _06310_ & ~_06664_;
	assign _06667_ = _05262_ | io_in[9];
	assign _06668_ = io_in[11] & ~_06667_;
	assign _06669_ = _06310_ & ~_04504_;
	assign _06670_ = _03608_ | _01208_;
	assign _06671_ = _06310_ & ~_06670_;
	assign _06672_ = _06290_ | io_in[5];
	assign _06673_ = _06672_ | _03759_;
	assign _06674_ = _06673_ | _02207_;
	assign _06675_ = _06674_ | _01208_;
	assign _06677_ = _01985_ & ~_06675_;
	assign _06678_ = _01651_ | _02207_;
	assign _06679_ = _06678_ | _02096_;
	assign _06680_ = _06310_ & ~_06679_;
	assign _06681_ = _06324_ | io_in[9];
	assign _06682_ = io_in[10] & ~_06681_;
	assign _06683_ = _02672_ | io_in[8];
	assign _06684_ = _06683_ | _02096_;
	assign _06685_ = _06684_ | io_in[10];
	assign _06686_ = _01985_ & ~_06685_;
	assign _06688_ = _01985_ & ~_05714_;
	assign _06689_ = io_in[11] & ~_07332_;
	assign _06690_ = _02285_ | io_in[5];
	assign _06691_ = _06690_ | io_in[7];
	assign _06692_ = _06691_ | io_in[8];
	assign _06693_ = _01985_ & ~_06692_;
	assign _06694_ = _01531_ | _06310_;
	assign _06695_ = _01985_ & ~_06694_;
	assign _06696_ = _04209_ | _01208_;
	assign _06697_ = io_in[10] & ~_06696_;
	assign _06699_ = io_in[11] & ~_05192_;
	assign _06700_ = _03535_ | io_in[8];
	assign _06701_ = _06700_ | _02096_;
	assign _06702_ = io_in[10] & ~_06701_;
	assign _06703_ = _05076_ | _02096_;
	assign _06704_ = _06310_ & ~_06703_;
	assign _06705_ = _04091_ | _03094_;
	assign _06706_ = _06705_ | io_in[6];
	assign _06707_ = _06706_ | _02207_;
	assign _06708_ = _06707_ | io_in[8];
	assign _06710_ = _06708_ | io_in[9];
	assign _06711_ = io_in[10] & ~_06710_;
	assign _06712_ = _00459_ | io_in[10];
	assign _06713_ = _01985_ & ~_06712_;
	assign _06714_ = _01411_ | _02207_;
	assign _06715_ = _06714_ | io_in[9];
	assign _06716_ = _06310_ & ~_06715_;
	assign _06717_ = _01017_ | io_in[5];
	assign _06718_ = _06717_ | _02207_;
	assign _06719_ = _06718_ | _02096_;
	assign _06721_ = io_in[11] & ~_06719_;
	assign _06722_ = _03260_ | _03759_;
	assign _06723_ = _06722_ | io_in[7];
	assign _06724_ = _06723_ | _01208_;
	assign _06725_ = _06724_ | _02096_;
	assign _06726_ = _01985_ & ~_06725_;
	assign _06727_ = _01234_ | io_in[7];
	assign _06728_ = _06727_ | _01208_;
	assign _06729_ = _06728_ | _06310_;
	assign _06730_ = _01985_ & ~_06729_;
	assign _06732_ = _02998_ | io_in[8];
	assign _06733_ = _06732_ | io_in[9];
	assign _06734_ = io_in[11] & ~_06733_;
	assign _06735_ = _01714_ | _03759_;
	assign _06736_ = _06735_ | io_in[8];
	assign _06737_ = _06736_ | io_in[9];
	assign _06738_ = io_in[11] & ~_06737_;
	assign _06739_ = _01902_ | io_in[8];
	assign _06740_ = io_in[11] & ~_06739_;
	assign _06741_ = _04047_ | io_in[5];
	assign _06743_ = _06741_ | _03759_;
	assign _06744_ = _06743_ | _02207_;
	assign _06745_ = _06744_ | _01208_;
	assign _06746_ = _06745_ | _02096_;
	assign _06747_ = _06310_ & ~_06746_;
	assign _06748_ = _01314_ | _02207_;
	assign _06749_ = _06748_ | _01208_;
	assign _06750_ = _06749_ | _02096_;
	assign _06751_ = _06750_ | _06310_;
	assign _06752_ = _01985_ & ~_06751_;
	assign _06755_ = _01735_ | io_in[6];
	assign _06756_ = _06755_ | _02207_;
	assign _06757_ = _06756_ | io_in[8];
	assign _06758_ = io_in[9] & ~_06757_;
	assign _06759_ = _03801_ | _01208_;
	assign _06760_ = _06759_ | _02096_;
	assign _06761_ = _06760_ | _06310_;
	assign _06762_ = _01985_ & ~_06761_;
	assign _06763_ = _04817_ | io_in[7];
	assign _06764_ = _06763_ | _01208_;
	assign _06766_ = _06764_ | _02096_;
	assign _06767_ = _06766_ | _06310_;
	assign _06768_ = _01985_ & ~_06767_;
	assign _06769_ = _01201_ | _02207_;
	assign _06770_ = _06769_ | _01208_;
	assign _06771_ = _06770_ | _02096_;
	assign _06772_ = io_in[10] & ~_06771_;
	assign _06773_ = _03188_ | io_in[7];
	assign _06774_ = _06773_ | io_in[8];
	assign _06775_ = _06774_ | _02096_;
	assign _06777_ = _06775_ | io_in[10];
	assign _06778_ = io_in[11] & ~_06777_;
	assign _06779_ = _04407_ | io_in[9];
	assign _06780_ = _01985_ & ~_06779_;
	assign _06781_ = _04382_ | _06310_;
	assign _06782_ = io_in[11] & ~_06781_;
	assign _06783_ = _06853_ | io_in[5];
	assign _06784_ = _06783_ | io_in[6];
	assign _06785_ = _06784_ | io_in[7];
	assign _06786_ = _06785_ | io_in[8];
	assign _06788_ = _06786_ | _02096_;
	assign _06789_ = io_in[11] & ~_06788_;
	assign _06790_ = _06442_ | io_in[9];
	assign _06791_ = _01985_ & ~_06790_;
	assign _06792_ = _01213_ | _02207_;
	assign _06793_ = _06792_ | io_in[9];
	assign _06794_ = io_in[11] & ~_06793_;
	assign _06795_ = _00599_ | io_in[7];
	assign _06796_ = _06795_ | _01208_;
	assign _06797_ = _06796_ | io_in[10];
	assign _06799_ = io_in[11] & ~_06797_;
	assign _06800_ = _07277_ & ~_06310_;
	assign _06801_ = _01376_ | _01208_;
	assign _06802_ = _06801_ | io_in[9];
	assign _06803_ = io_in[10] & ~_06802_;
	assign _06804_ = _02751_ | io_in[7];
	assign _06805_ = _06804_ | io_in[8];
	assign _06806_ = _06805_ | io_in[10];
	assign _06807_ = _01985_ & ~_06806_;
	assign _06808_ = _00235_ | _03759_;
	assign _06810_ = _06808_ | _02207_;
	assign _06811_ = _06810_ | io_in[8];
	assign _06812_ = _06811_ | _02096_;
	assign _06813_ = io_in[10] & ~_06812_;
	assign _06814_ = _00708_ | _03759_;
	assign _06815_ = _06814_ | io_in[7];
	assign _06816_ = _06815_ | _01208_;
	assign _06817_ = _06816_ | io_in[9];
	assign _06818_ = io_in[10] & ~_06817_;
	assign _06819_ = _06975_ | _03759_;
	assign _06821_ = _06819_ | _02207_;
	assign _06822_ = _06821_ | _02096_;
	assign _06823_ = _06822_ | io_in[10];
	assign _06824_ = io_in[11] & ~_06823_;
	assign _06825_ = _05031_ | io_in[6];
	assign _06826_ = _06825_ | _02207_;
	assign _06827_ = _06826_ | io_in[8];
	assign _06828_ = _06827_ | io_in[9];
	assign _06829_ = io_in[11] & ~_06828_;
	assign _06830_ = _07383_ | io_in[7];
	assign _06832_ = _06830_ | io_in[8];
	assign _06833_ = _06832_ | io_in[10];
	assign _06834_ = _01985_ & ~_06833_;
	assign _06835_ = _01878_ | io_in[7];
	assign _06836_ = _06835_ | _02096_;
	assign _06837_ = _06836_ | io_in[10];
	assign _06838_ = io_in[11] & ~_06837_;
	assign _06839_ = _00267_ | io_in[6];
	assign _06840_ = _06839_ | _02207_;
	assign _06841_ = _06840_ | _01208_;
	assign _06843_ = _06841_ | _02096_;
	assign _06844_ = _06843_ | _06310_;
	assign _06845_ = _01985_ & ~_06844_;
	assign _06846_ = _01086_ | _03759_;
	assign _06847_ = _06846_ | _02207_;
	assign _06848_ = _06847_ | _01208_;
	assign _06849_ = _06848_ | io_in[9];
	assign _06850_ = io_in[11] & ~_06849_;
	assign _06851_ = _04114_ | io_in[8];
	assign _06852_ = _06851_ | io_in[9];
	assign _06854_ = io_in[10] & ~_06852_;
	assign _06855_ = _04458_ | io_in[6];
	assign _06856_ = _06855_ | io_in[7];
	assign _06857_ = _06856_ | io_in[8];
	assign _06858_ = _02096_ & ~_06857_;
	assign _06859_ = _00729_ | _02207_;
	assign _06860_ = _06859_ | _01208_;
	assign _06861_ = _06860_ | io_in[9];
	assign _06862_ = io_in[11] & ~_06861_;
	assign _06863_ = _06483_ | io_in[10];
	assign _06866_ = io_in[11] & ~_06863_;
	assign _06867_ = _01469_ | _02207_;
	assign _06868_ = _06867_ | io_in[8];
	assign _06869_ = _06868_ | _02096_;
	assign _06870_ = _01985_ & ~_06869_;
	assign _06871_ = _05590_ | _02096_;
	assign _06872_ = io_in[10] & ~_06871_;
	assign _06873_ = _05352_ | _02207_;
	assign _06874_ = _06873_ | io_in[8];
	assign _06875_ = _06874_ | io_in[9];
	assign _06877_ = _06875_ | _06310_;
	assign _06878_ = _01985_ & ~_06877_;
	assign _06879_ = _07360_ | io_in[10];
	assign _06880_ = _01985_ & ~_06879_;
	assign _06881_ = _03558_ | io_in[8];
	assign _06882_ = io_in[9] & ~_06881_;
	assign _06883_ = _03685_ | _02207_;
	assign _06884_ = io_in[8] & ~_06883_;
	assign _06885_ = _07283_ | io_in[6];
	assign _06886_ = _06885_ | _02207_;
	assign _06888_ = _06886_ | io_in[8];
	assign _06889_ = _06888_ | _02096_;
	assign _06890_ = _06310_ & ~_06889_;
	assign _06891_ = _05629_ | io_in[10];
	assign _06892_ = _01985_ & ~_06891_;
	assign _06893_ = _06056_ | io_in[9];
	assign _06894_ = io_in[10] & ~_06893_;
	assign _06895_ = _07275_ | io_in[9];
	assign _06896_ = _06895_ | io_in[10];
	assign _06897_ = _01985_ & ~_06896_;
	assign _06899_ = _07301_ | _03759_;
	assign _06900_ = _06899_ | _01208_;
	assign _06901_ = _06900_ | io_in[9];
	assign _06902_ = _06901_ | io_in[10];
	assign _06903_ = _01985_ & ~_06902_;
	assign _06904_ = _06125_ | io_in[9];
	assign _06905_ = io_in[11] & ~_06904_;
	assign _06906_ = _00175_ | _02207_;
	assign _06907_ = _06906_ | io_in[8];
	assign _06908_ = _06907_ | _02096_;
	assign _06910_ = io_in[11] & ~_06908_;
	assign _06911_ = _07120_ | io_in[8];
	assign _06912_ = _06911_ | io_in[9];
	assign _06913_ = _01985_ & ~_06912_;
	assign _06914_ = _03033_ | _03759_;
	assign _06915_ = _06914_ | _02207_;
	assign _06916_ = _06915_ | io_in[8];
	assign _06917_ = io_in[10] & ~_06916_;
	assign _06918_ = _04272_ | io_in[8];
	assign _06919_ = _06918_ | io_in[9];
	assign _06921_ = _06310_ & ~_06919_;
	assign _06922_ = _03404_ | _03759_;
	assign _06923_ = _06922_ | _02207_;
	assign _06924_ = _06923_ | io_in[8];
	assign _06925_ = _06924_ | _02096_;
	assign _06926_ = io_in[11] & ~_06925_;
	assign _06927_ = _02629_ | _06310_;
	assign _06928_ = _01985_ & ~_06927_;
	assign _06929_ = _02555_ | io_in[7];
	assign _06930_ = _06929_ | _01208_;
	assign _06932_ = io_in[10] & ~_06930_;
	assign _06933_ = _00173_ | _03759_;
	assign _06934_ = _06933_ | _02207_;
	assign _06935_ = _06934_ | _01208_;
	assign _06936_ = _02096_ & ~_06935_;
	assign _06937_ = (io_in[11] ? _06936_ : _06932_);
	assign _06938_ = _06937_ | _06928_;
	assign _06939_ = _06938_ | _06926_;
	assign _06940_ = _06939_ | _06921_;
	assign _06941_ = _06940_ | _06917_;
	assign _06943_ = _06941_ | _06913_;
	assign _06944_ = _06943_ | _06910_;
	assign _06945_ = _06944_ | _06905_;
	assign _06946_ = _06945_ | _06903_;
	assign _06947_ = _06946_ | _06897_;
	assign _06948_ = _06947_ | _06894_;
	assign _06949_ = _06948_ | _06892_;
	assign _06950_ = _06949_ | _06890_;
	assign _06951_ = _06950_ | _06884_;
	assign _06952_ = _06951_ | _06882_;
	assign _06954_ = _06952_ | _06880_;
	assign _06955_ = _06954_ | _06878_;
	assign _06956_ = _06955_ | _06872_;
	assign _06957_ = _06956_ | _06870_;
	assign _06958_ = _06957_ | _06866_;
	assign _06959_ = _06958_ | _02553_;
	assign _06960_ = _06959_ | _06862_;
	assign _06961_ = _06960_ | _06858_;
	assign _06962_ = _06961_ | _06854_;
	assign _06963_ = _06962_ | _06850_;
	assign _06965_ = _06963_ | _06845_;
	assign _06966_ = _06965_ | _06838_;
	assign _06967_ = _06966_ | _06834_;
	assign _06968_ = _06967_ | _06829_;
	assign _06969_ = _06968_ | _06824_;
	assign _06970_ = _06969_ | _06818_;
	assign _06971_ = _06970_ | _06813_;
	assign _06972_ = _06971_ | _06807_;
	assign _06973_ = _06972_ | _06803_;
	assign _06974_ = _06973_ | _06800_;
	assign _06977_ = _06974_ | _06799_;
	assign _06978_ = _06977_ | _06794_;
	assign _06979_ = _06978_ | _06791_;
	assign _06980_ = _06979_ | _06789_;
	assign _06981_ = _06980_ | _06782_;
	assign _06982_ = _06981_ | _06780_;
	assign _06983_ = _06982_ | _06778_;
	assign _06984_ = _06983_ | _06772_;
	assign _06985_ = _06984_ | _06768_;
	assign _06986_ = _06985_ | _06762_;
	assign _06988_ = _06986_ | _06758_;
	assign _06989_ = _06988_ | _06752_;
	assign _06990_ = _06989_ | _06747_;
	assign _06991_ = _06990_ | _06740_;
	assign _06992_ = _06991_ | _06738_;
	assign _06993_ = _06992_ | _06734_;
	assign _06994_ = _06993_ | _06730_;
	assign _06995_ = _06994_ | _06726_;
	assign _06996_ = _06995_ | _06721_;
	assign _06997_ = _06996_ | _05524_;
	assign _06999_ = _06997_ | _06716_;
	assign _07000_ = _06999_ | _06713_;
	assign _07001_ = _07000_ | _06711_;
	assign _07002_ = _07001_ | _06704_;
	assign _07003_ = _07002_ | _06702_;
	assign _07004_ = _07003_ | _03087_;
	assign _07005_ = _07004_ | _06699_;
	assign _07006_ = _07005_ | _06697_;
	assign _07007_ = _07006_ | _06695_;
	assign _07008_ = _07007_ | _06693_;
	assign _07010_ = _07008_ | _06689_;
	assign _07011_ = _07010_ | _06688_;
	assign _07012_ = _07011_ | _06686_;
	assign _07013_ = _07012_ | _06682_;
	assign _07014_ = _07013_ | _06680_;
	assign _07015_ = _07014_ | _06677_;
	assign _07016_ = _07015_ | _06671_;
	assign _07017_ = _07016_ | _06669_;
	assign _07018_ = _07017_ | _06668_;
	assign _07019_ = _07018_ | _06666_;
	assign _07021_ = _07019_ | _01816_;
	assign _07022_ = _07021_ | _06662_;
	assign _07023_ = _07022_ | _06659_;
	assign _07024_ = _07023_ | _06657_;
	assign _07025_ = _07024_ | _06656_;
	assign _07026_ = _07025_ | _06652_;
	assign _07027_ = _07026_ | _06651_;
	assign _07028_ = _07027_ | _06647_;
	assign _07029_ = _07028_ | _06645_;
	assign _07030_ = _07029_ | _06640_;
	assign _07032_ = _07030_ | _06638_;
	assign _07033_ = _07032_ | _06637_;
	assign _07034_ = _07033_ | _06632_;
	assign _07035_ = _07034_ | _06628_;
	assign _07036_ = _07035_ | _06623_;
	assign _07037_ = _07036_ | _06622_;
	assign _07038_ = _07037_ | _06616_;
	assign _07039_ = _07038_ | _06614_;
	assign _07040_ = _07039_ | _06611_;
	assign _07041_ = _07040_ | _04111_;
	assign _07043_ = _07041_ | _06608_;
	assign _07044_ = _07043_ | _06604_;
	assign _07045_ = _07044_ | _06602_;
	assign _07046_ = _07045_ | _06599_;
	assign _07047_ = _07046_ | _06594_;
	assign _07048_ = _07047_ | _06592_;
	assign _07049_ = _07048_ | _01204_;
	assign _07050_ = _07049_ | _04101_;
	assign _07051_ = _07050_ | _06590_;
	assign _07052_ = _07051_ | _06585_;
	assign _07054_ = _07052_ | _06581_;
	assign _07055_ = _07054_ | _06575_;
	assign _07056_ = _07055_ | _06571_;
	assign _07057_ = _07056_ | _06569_;
	assign _07058_ = _07057_ | _06566_;
	assign _07059_ = _07058_ | _06560_;
	assign _07060_ = _07059_ | _06558_;
	assign _07061_ = _07060_ | _06557_;
	assign _07062_ = _07061_ | _06556_;
	assign _07063_ = _07062_ | _06551_;
	assign _07065_ = _07063_ | _06547_;
	assign _07066_ = _07065_ | _06542_;
	assign _07067_ = _07066_ | _01646_;
	assign _07068_ = _07067_ | _06538_;
	assign _07069_ = _07068_ | _06534_;
	assign _07070_ = _07069_ | _06530_;
	assign _07071_ = _07070_ | _06528_;
	assign _07072_ = _07071_ | _06525_;
	assign _07073_ = _07072_ | _06521_;
	assign _07074_ = _07073_ | _06515_;
	assign _07076_ = _07074_ | _06511_;
	assign _07077_ = _07076_ | _06506_;
	assign _07078_ = _07077_ | _06502_;
	assign _07079_ = _07078_ | _06497_;
	assign _07080_ = _07079_ | _06494_;
	assign _07081_ = _07080_ | _05284_;
	assign _07082_ = _07081_ | _06492_;
	assign _07083_ = _07082_ | _06486_;
	assign _07084_ = _07083_ | _06482_;
	assign _07085_ = _07084_ | _06479_;
	assign _07088_ = _07085_ | _06475_;
	assign _07089_ = _07088_ | _06473_;
	assign _07090_ = _07089_ | _06470_;
	assign _07091_ = _07090_ | _06466_;
	assign _07092_ = _07091_ | _06462_;
	assign _07093_ = _07092_ | _02792_;
	assign _07094_ = _07093_ | _06459_;
	assign _07095_ = _07094_ | _06456_;
	assign _07096_ = _07095_ | _06451_;
	assign _07097_ = _07096_ | _06448_;
	assign _07099_ = _07097_ | _06445_;
	assign _07100_ = _07099_ | _06441_;
	assign _07101_ = _07100_ | _06439_;
	assign _07102_ = _07101_ | _06437_;
	assign _07103_ = _07102_ | _06433_;
	assign _07104_ = _07103_ | _06428_;
	assign _07105_ = _07104_ | _06424_;
	assign _07106_ = _07105_ | _06419_;
	assign _07107_ = _07106_ | _06416_;
	assign _07108_ = _07107_ | _06412_;
	assign _07110_ = _07108_ | _06408_;
	assign _07111_ = _07110_ | _06406_;
	assign _07112_ = _07111_ | _06402_;
	assign _07113_ = _07112_ | _06396_;
	assign _07114_ = _07113_ | _06393_;
	assign _07115_ = _07114_ | _06390_;
	assign _07116_ = _07115_ | _06388_;
	assign _07117_ = _07116_ | _06384_;
	assign _07118_ = _07117_ | _06383_;
	assign _07119_ = _07118_ | _06382_;
	assign _07121_ = _07119_ | _06378_;
	assign _07122_ = _07121_ | _06375_;
	assign _07123_ = _07122_ | _06373_;
	assign _07124_ = _07123_ | _06370_;
	assign _07125_ = _07124_ | _06367_;
	assign _07126_ = _07125_ | _06363_;
	assign _07127_ = _07126_ | _06361_;
	assign _07128_ = _07127_ | _06357_;
	assign _07129_ = _07128_ | _03853_;
	assign _07130_ = _07129_ | _06350_;
	assign _07132_ = _07130_ | _06348_;
	assign _07133_ = _07132_ | _06342_;
	assign _07134_ = _07133_ | _06336_;
	assign _07135_ = _07134_ | _06334_;
	assign _07136_ = _07135_ | _06330_;
	assign _07137_ = _07136_ | _06327_;
	assign _07138_ = _07137_ | _06323_;
	assign _07139_ = _07138_ | _06318_;
	assign _07140_ = _07139_ | _06313_;
	assign _07141_ = _07140_ | _06308_;
	assign _07143_ = _07141_ | _06307_;
	assign _07144_ = _07143_ | _06305_;
	assign _07145_ = _07144_ | _06302_;
	assign _07146_ = _07145_ | _06300_;
	assign _07147_ = _07146_ | _06295_;
	assign _07148_ = _07147_ | _06289_;
	assign _07149_ = _07148_ | _06286_;
	assign _07150_ = _07149_ | _06284_;
	assign _07151_ = _07150_ | _06282_;
	assign _07152_ = _07151_ | _06279_;
	assign _07154_ = _07152_ | _06277_;
	assign _07155_ = _07154_ | _06273_;
	assign _07156_ = _07155_ | _06271_;
	assign _07157_ = _07156_ | _06267_;
	assign _07158_ = _07157_ | _06263_;
	assign _07159_ = _07158_ | _06258_;
	assign _07160_ = _07159_ | _06255_;
	assign _07161_ = _07160_ | _06251_;
	assign _07162_ = _07161_ | _06250_;
	assign _07163_ = _07162_ | _06248_;
	assign _07165_ = _07163_ | _06245_;
	assign _07166_ = _07165_ | _06241_;
	assign _07167_ = _07166_ | _06240_;
	assign _07168_ = _07167_ | _06239_;
	assign _07169_ = _07168_ | _03691_;
	assign _07170_ = _07169_ | _06235_;
	assign _07171_ = _07170_ | _06233_;
	assign _07172_ = _07171_ | _06229_;
	assign _07173_ = _07172_ | _06227_;
	assign _07174_ = _07173_ | _06224_;
	assign _07176_ = _07174_ | _06223_;
	assign _07177_ = _07176_ | _06220_;
	assign _07178_ = _07177_ | _06218_;
	assign _07179_ = _07178_ | _06216_;
	assign _07180_ = _07179_ | _06212_;
	assign _07181_ = _07180_ | _06208_;
	assign _07182_ = _07181_ | _06204_;
	assign _07183_ = _07182_ | _06201_;
	assign _07184_ = _07183_ | _06200_;
	assign _07185_ = _07184_ | _06192_;
	assign _07187_ = _07185_ | _06190_;
	assign _07188_ = _07187_ | _06186_;
	assign _07189_ = _07188_ | _06185_;
	assign _07190_ = _07189_ | _06182_;
	assign _07191_ = _07190_ | _06178_;
	assign _07192_ = _07191_ | _06175_;
	assign _07193_ = _07192_ | _06173_;
	assign _07194_ = _07193_ | _06169_;
	assign _07195_ = _07194_ | _06168_;
	assign _07196_ = _07195_ | _06163_;
	assign _07199_ = _07196_ | _06161_;
	assign _07200_ = _07199_ | _06159_;
	assign _07201_ = _07200_ | _06158_;
	assign _07202_ = _07201_ | _06155_;
	assign _07203_ = _07202_ | _06149_;
	assign _07204_ = _07203_ | _06142_;
	assign _07205_ = _07204_ | _06137_;
	assign _07206_ = _07205_ | _06135_;
	assign _07207_ = _07206_ | _06128_;
	assign _07208_ = _07207_ | _06124_;
	assign _07210_ = _07208_ | _06119_;
	assign _07211_ = _07210_ | _06114_;
	assign _07212_ = _07211_ | _06109_;
	assign _07213_ = _07212_ | _06106_;
	assign _07214_ = _07213_ | _06103_;
	assign _07215_ = _07214_ | _06100_;
	assign _07216_ = _07215_ | _06097_;
	assign _07217_ = _07216_ | _06094_;
	assign _07218_ = _07217_ | _06093_;
	assign _07219_ = _07218_ | _06090_;
	assign _07221_ = _07219_ | _06082_;
	assign _07222_ = _07221_ | _06079_;
	assign _07223_ = _07222_ | _06073_;
	assign _07224_ = _07223_ | _06069_;
	assign _07225_ = _07224_ | _06067_;
	assign _07226_ = _07225_ | _06063_;
	assign _07227_ = _07226_ | _06059_;
	assign _07228_ = _07227_ | _06057_;
	assign _07229_ = _07228_ | _06055_;
	assign _07230_ = _07229_ | _06051_;
	assign _07232_ = _07230_ | _06048_;
	assign _07233_ = _07232_ | _06045_;
	assign _07234_ = _07233_ | _06042_;
	assign _07235_ = _07234_ | _06038_;
	assign _07236_ = _07235_ | _06034_;
	assign _07237_ = _07236_ | _06028_;
	assign _07238_ = _07237_ | _06027_;
	assign \mchip.val [0] = _07238_ | _06026_;
	reg \mchip.io_out_reg[0] ;
	always @(posedge io_in[12]) \mchip.io_out_reg[0]  <= \mchip.val [0];
	assign \mchip.io_out [0] = \mchip.io_out_reg[0] ;
	reg \mchip.io_out_reg[1] ;
	always @(posedge io_in[12]) \mchip.io_out_reg[1]  <= \mchip.val [1];
	assign \mchip.io_out [1] = \mchip.io_out_reg[1] ;
	reg \mchip.io_out_reg[2] ;
	always @(posedge io_in[12]) \mchip.io_out_reg[2]  <= \mchip.val [2];
	assign \mchip.io_out [2] = \mchip.io_out_reg[2] ;
	reg \mchip.io_out_reg[3] ;
	always @(posedge io_in[12]) \mchip.io_out_reg[3]  <= \mchip.val [3];
	assign \mchip.io_out [3] = \mchip.io_out_reg[3] ;
	reg \mchip.io_out_reg[4] ;
	always @(posedge io_in[12]) \mchip.io_out_reg[4]  <= \mchip.val [4];
	assign \mchip.io_out [4] = \mchip.io_out_reg[4] ;
	reg \mchip.io_out_reg[5] ;
	always @(posedge io_in[12]) \mchip.io_out_reg[5]  <= \mchip.val [5];
	assign \mchip.io_out [5] = \mchip.io_out_reg[5] ;
	reg \mchip.io_out_reg[6] ;
	always @(posedge io_in[12]) \mchip.io_out_reg[6]  <= \mchip.val [6];
	assign \mchip.io_out [6] = \mchip.io_out_reg[6] ;
	assign io_out = {7'h00, \mchip.io_out [6:0]};
	assign \mchip.clock  = io_in[12];
	assign \mchip.io_in  = io_in[11:0];
	assign \mchip.io_out [11:7] = 5'h00;
	assign \mchip.reset  = io_in[13];
	assign \mchip.val [7] = 1'h0;
endmodule
module d11_gbailey_bfchip (
	io_in,
	io_out
);
	wire _0000_;
	wire _0001_;
	wire _0002_;
	wire _0003_;
	wire _0004_;
	wire _0005_;
	wire _0006_;
	wire _0007_;
	wire _0008_;
	wire _0009_;
	wire _0010_;
	wire _0011_;
	wire _0012_;
	wire _0013_;
	wire _0014_;
	wire _0015_;
	wire _0016_;
	wire _0017_;
	wire _0018_;
	wire _0019_;
	wire _0020_;
	wire _0021_;
	wire _0022_;
	wire _0023_;
	wire _0024_;
	wire _0025_;
	wire _0026_;
	wire _0027_;
	wire _0028_;
	wire _0029_;
	wire _0030_;
	wire _0031_;
	wire _0032_;
	wire _0033_;
	wire _0034_;
	wire _0035_;
	wire _0036_;
	wire _0037_;
	wire _0038_;
	wire _0039_;
	wire _0040_;
	wire _0041_;
	wire _0042_;
	wire _0043_;
	wire _0044_;
	wire _0045_;
	wire _0046_;
	wire _0047_;
	wire _0048_;
	wire _0049_;
	wire _0050_;
	wire _0051_;
	wire _0052_;
	wire _0053_;
	wire _0054_;
	wire _0055_;
	wire _0056_;
	wire _0057_;
	wire _0058_;
	wire _0059_;
	wire _0060_;
	wire _0061_;
	wire _0062_;
	wire _0063_;
	wire _0064_;
	wire _0065_;
	wire _0066_;
	wire _0067_;
	wire _0068_;
	wire _0069_;
	wire _0070_;
	wire _0071_;
	wire _0072_;
	wire _0073_;
	wire _0074_;
	wire _0075_;
	wire _0076_;
	wire _0077_;
	wire _0078_;
	wire _0079_;
	wire _0080_;
	wire _0081_;
	wire _0082_;
	wire _0083_;
	wire _0084_;
	wire _0085_;
	wire _0086_;
	wire _0087_;
	wire _0088_;
	wire _0089_;
	wire _0090_;
	wire _0091_;
	wire _0092_;
	wire _0093_;
	wire _0094_;
	wire _0095_;
	wire _0096_;
	wire _0097_;
	wire _0098_;
	wire _0099_;
	wire _0100_;
	wire _0101_;
	wire _0102_;
	wire _0103_;
	wire _0104_;
	wire _0105_;
	wire _0106_;
	wire _0107_;
	wire _0108_;
	wire _0109_;
	wire _0110_;
	wire _0111_;
	wire _0112_;
	wire _0113_;
	wire _0114_;
	wire _0115_;
	wire _0116_;
	wire _0117_;
	wire _0118_;
	wire _0119_;
	wire _0120_;
	wire _0121_;
	wire _0122_;
	wire _0123_;
	wire _0124_;
	wire _0125_;
	wire _0126_;
	wire _0127_;
	wire _0128_;
	wire _0129_;
	wire _0130_;
	wire _0131_;
	wire _0132_;
	wire _0133_;
	wire _0134_;
	wire _0135_;
	wire _0136_;
	wire _0137_;
	wire _0138_;
	wire _0139_;
	wire _0140_;
	wire _0141_;
	wire _0142_;
	wire _0143_;
	wire _0144_;
	wire _0145_;
	wire _0146_;
	wire _0147_;
	wire _0148_;
	wire _0149_;
	wire _0150_;
	wire _0151_;
	wire _0152_;
	wire _0153_;
	wire _0154_;
	wire _0155_;
	wire _0156_;
	wire _0157_;
	wire _0158_;
	wire _0159_;
	wire _0160_;
	wire _0161_;
	wire _0162_;
	wire _0163_;
	wire _0164_;
	wire _0165_;
	wire _0166_;
	wire _0167_;
	wire _0168_;
	wire _0169_;
	wire _0170_;
	wire _0171_;
	wire _0172_;
	wire _0173_;
	wire _0174_;
	wire _0175_;
	wire _0176_;
	wire _0177_;
	wire _0178_;
	wire _0179_;
	wire _0180_;
	wire _0181_;
	wire _0182_;
	wire _0183_;
	wire _0184_;
	wire _0185_;
	wire _0186_;
	wire _0187_;
	wire _0188_;
	wire _0189_;
	wire _0190_;
	wire _0191_;
	wire _0192_;
	wire _0193_;
	wire _0194_;
	wire _0195_;
	wire _0196_;
	wire _0197_;
	wire _0198_;
	wire _0199_;
	wire _0200_;
	wire _0201_;
	wire _0202_;
	wire _0203_;
	wire _0204_;
	wire _0205_;
	wire _0206_;
	wire _0207_;
	wire _0208_;
	wire _0209_;
	wire _0210_;
	wire _0211_;
	wire _0212_;
	wire _0213_;
	wire _0214_;
	wire _0215_;
	wire _0216_;
	wire _0217_;
	wire _0218_;
	wire _0219_;
	wire _0220_;
	wire _0221_;
	wire _0222_;
	wire _0223_;
	wire _0224_;
	wire _0225_;
	wire _0226_;
	wire _0227_;
	wire _0228_;
	wire _0229_;
	wire _0230_;
	wire _0231_;
	wire _0232_;
	wire _0233_;
	wire _0234_;
	wire _0235_;
	wire _0236_;
	wire _0237_;
	wire _0238_;
	wire _0239_;
	wire _0240_;
	wire _0241_;
	wire _0242_;
	wire _0243_;
	wire _0244_;
	wire _0245_;
	wire _0246_;
	wire _0247_;
	wire _0248_;
	wire _0249_;
	wire _0250_;
	wire _0251_;
	wire _0252_;
	wire _0253_;
	wire _0254_;
	wire _0255_;
	wire _0256_;
	wire _0257_;
	wire _0258_;
	wire _0259_;
	wire _0260_;
	wire _0261_;
	wire _0262_;
	wire _0263_;
	wire _0264_;
	wire _0265_;
	wire _0266_;
	wire _0267_;
	wire _0268_;
	wire _0269_;
	wire _0270_;
	wire _0271_;
	wire _0272_;
	wire _0273_;
	wire _0274_;
	wire _0275_;
	wire _0276_;
	wire _0277_;
	wire _0278_;
	wire _0279_;
	wire _0280_;
	wire _0281_;
	wire _0282_;
	wire _0283_;
	wire _0284_;
	wire _0285_;
	wire _0286_;
	wire _0287_;
	wire _0288_;
	wire _0289_;
	wire _0290_;
	wire _0291_;
	wire _0292_;
	wire _0293_;
	wire _0294_;
	wire _0295_;
	wire _0296_;
	wire _0297_;
	wire _0298_;
	wire _0299_;
	wire _0300_;
	wire _0301_;
	wire _0302_;
	wire _0303_;
	wire _0304_;
	wire _0305_;
	wire _0306_;
	wire _0307_;
	wire _0308_;
	wire _0309_;
	wire _0310_;
	wire _0311_;
	wire _0312_;
	wire _0313_;
	wire _0314_;
	wire _0315_;
	wire _0316_;
	wire _0317_;
	wire _0318_;
	wire _0319_;
	wire _0320_;
	wire _0321_;
	wire _0322_;
	wire _0323_;
	wire _0324_;
	wire _0325_;
	wire _0326_;
	wire _0327_;
	wire _0328_;
	wire _0329_;
	wire _0330_;
	wire _0331_;
	wire _0332_;
	wire _0333_;
	wire _0334_;
	wire _0335_;
	wire _0336_;
	wire _0337_;
	wire _0338_;
	wire _0339_;
	wire _0340_;
	wire _0341_;
	wire _0342_;
	wire _0343_;
	wire _0344_;
	wire _0345_;
	wire _0346_;
	wire _0347_;
	wire _0348_;
	wire _0349_;
	wire _0350_;
	wire _0351_;
	wire _0352_;
	wire _0353_;
	wire _0354_;
	wire _0355_;
	wire _0356_;
	wire _0357_;
	wire _0358_;
	wire _0359_;
	wire _0360_;
	wire _0361_;
	wire _0362_;
	wire _0363_;
	wire _0364_;
	wire _0365_;
	wire _0366_;
	wire _0367_;
	wire _0368_;
	wire _0369_;
	wire _0370_;
	wire _0371_;
	wire _0372_;
	wire _0373_;
	wire _0374_;
	wire _0375_;
	wire _0376_;
	wire _0377_;
	wire _0378_;
	wire _0379_;
	wire _0380_;
	wire _0381_;
	wire _0382_;
	wire _0383_;
	wire _0384_;
	wire _0385_;
	wire _0386_;
	wire _0387_;
	wire _0388_;
	wire _0389_;
	wire _0390_;
	wire _0391_;
	wire _0392_;
	wire _0393_;
	wire _0394_;
	wire _0395_;
	wire _0396_;
	wire _0397_;
	wire _0398_;
	wire _0399_;
	wire _0400_;
	wire _0401_;
	wire _0402_;
	wire _0403_;
	wire _0404_;
	wire _0405_;
	wire _0406_;
	wire _0407_;
	wire _0408_;
	wire _0409_;
	wire _0410_;
	wire _0411_;
	wire _0412_;
	wire _0413_;
	wire _0414_;
	wire _0415_;
	wire _0416_;
	wire _0417_;
	wire _0418_;
	wire _0419_;
	wire _0420_;
	wire _0421_;
	wire _0422_;
	wire _0423_;
	wire _0424_;
	wire _0425_;
	wire _0426_;
	wire _0427_;
	wire _0428_;
	wire _0429_;
	wire _0430_;
	wire _0431_;
	wire _0432_;
	wire _0433_;
	wire _0434_;
	wire _0435_;
	wire _0436_;
	wire _0437_;
	wire _0438_;
	wire _0439_;
	wire _0440_;
	wire _0441_;
	wire _0442_;
	wire _0443_;
	wire _0444_;
	wire _0445_;
	wire _0446_;
	wire _0447_;
	wire _0448_;
	wire _0449_;
	wire _0450_;
	wire _0451_;
	wire _0452_;
	wire _0453_;
	wire _0454_;
	wire _0455_;
	wire _0456_;
	wire _0457_;
	wire _0458_;
	wire _0459_;
	wire _0460_;
	wire _0461_;
	wire _0462_;
	wire _0463_;
	wire _0464_;
	wire _0465_;
	wire _0466_;
	wire _0467_;
	wire _0468_;
	wire _0469_;
	wire _0470_;
	wire _0471_;
	wire _0472_;
	wire _0473_;
	wire _0474_;
	wire _0475_;
	wire _0476_;
	wire _0477_;
	wire _0478_;
	wire _0479_;
	wire _0480_;
	wire _0481_;
	wire _0482_;
	wire _0483_;
	wire _0484_;
	wire _0485_;
	wire _0486_;
	wire _0487_;
	wire _0488_;
	wire _0489_;
	wire _0490_;
	wire _0491_;
	wire _0492_;
	wire _0493_;
	wire _0494_;
	wire _0495_;
	wire _0496_;
	wire _0497_;
	wire _0498_;
	wire _0499_;
	wire _0500_;
	wire _0501_;
	wire _0502_;
	wire _0503_;
	wire _0504_;
	wire _0505_;
	wire _0506_;
	wire _0507_;
	wire _0508_;
	wire _0509_;
	wire _0510_;
	wire _0511_;
	wire _0512_;
	wire _0513_;
	wire _0514_;
	wire _0515_;
	wire _0516_;
	wire _0517_;
	wire _0518_;
	wire _0519_;
	wire _0520_;
	wire _0521_;
	wire _0522_;
	wire _0523_;
	wire _0524_;
	wire _0525_;
	wire _0526_;
	wire _0527_;
	wire _0528_;
	wire _0529_;
	wire _0530_;
	wire _0531_;
	wire _0532_;
	wire _0533_;
	wire _0534_;
	wire _0535_;
	wire _0536_;
	wire _0537_;
	wire _0538_;
	wire _0539_;
	wire _0540_;
	wire _0541_;
	wire _0542_;
	wire _0543_;
	wire _0544_;
	wire _0545_;
	wire _0546_;
	wire _0547_;
	wire _0548_;
	wire _0549_;
	wire _0550_;
	wire _0551_;
	wire _0552_;
	wire _0553_;
	wire _0554_;
	wire _0555_;
	wire _0556_;
	wire _0557_;
	wire _0558_;
	wire _0559_;
	wire _0560_;
	wire _0561_;
	wire _0562_;
	wire _0563_;
	wire _0564_;
	wire _0565_;
	wire _0566_;
	wire _0567_;
	wire _0568_;
	wire _0569_;
	wire _0570_;
	wire _0571_;
	wire _0572_;
	wire _0573_;
	wire _0574_;
	wire _0575_;
	wire _0576_;
	wire _0577_;
	wire _0578_;
	wire _0579_;
	wire _0580_;
	wire _0581_;
	wire _0582_;
	wire _0583_;
	wire _0584_;
	wire _0585_;
	wire _0586_;
	wire _0587_;
	wire _0588_;
	wire _0589_;
	wire _0590_;
	wire _0591_;
	wire _0592_;
	wire _0593_;
	wire _0594_;
	wire _0595_;
	wire _0596_;
	wire _0597_;
	wire _0598_;
	wire _0599_;
	wire _0600_;
	wire _0601_;
	wire _0602_;
	wire _0603_;
	wire _0604_;
	wire _0605_;
	wire _0606_;
	wire _0607_;
	wire _0608_;
	wire _0609_;
	wire _0610_;
	wire _0611_;
	wire _0612_;
	wire _0613_;
	wire _0614_;
	wire _0615_;
	wire _0616_;
	wire _0617_;
	wire _0618_;
	wire _0619_;
	wire _0620_;
	wire _0621_;
	wire _0622_;
	wire _0623_;
	wire _0624_;
	wire _0625_;
	wire _0626_;
	wire _0627_;
	wire _0628_;
	wire _0629_;
	wire _0630_;
	wire _0631_;
	wire _0632_;
	wire _0633_;
	wire _0634_;
	wire _0635_;
	wire _0636_;
	wire _0637_;
	wire _0638_;
	wire _0639_;
	wire _0640_;
	wire _0641_;
	wire _0642_;
	wire _0643_;
	wire _0644_;
	wire _0645_;
	wire _0646_;
	wire _0647_;
	wire _0648_;
	wire _0649_;
	wire _0650_;
	wire _0651_;
	wire _0652_;
	wire _0653_;
	wire _0654_;
	wire _0655_;
	wire _0656_;
	wire _0657_;
	wire _0658_;
	wire _0659_;
	wire _0660_;
	wire _0661_;
	wire _0662_;
	wire _0663_;
	wire _0664_;
	wire _0665_;
	wire _0666_;
	wire _0667_;
	wire _0668_;
	wire _0669_;
	wire _0670_;
	wire _0671_;
	wire _0672_;
	wire _0673_;
	wire _0674_;
	wire _0675_;
	wire _0676_;
	wire _0677_;
	wire _0678_;
	wire _0679_;
	wire _0680_;
	wire _0681_;
	wire _0682_;
	wire _0683_;
	wire _0684_;
	wire _0685_;
	wire _0686_;
	wire _0687_;
	wire _0688_;
	wire _0689_;
	wire _0690_;
	wire _0691_;
	wire _0692_;
	wire _0693_;
	wire _0694_;
	wire _0695_;
	wire _0696_;
	wire _0697_;
	wire _0698_;
	wire _0699_;
	wire _0700_;
	wire _0701_;
	wire _0702_;
	wire _0703_;
	wire _0704_;
	wire _0705_;
	wire _0706_;
	wire _0707_;
	wire _0708_;
	wire _0709_;
	wire _0710_;
	wire _0711_;
	wire _0712_;
	wire _0713_;
	wire _0714_;
	wire _0715_;
	wire _0716_;
	wire _0717_;
	wire _0718_;
	wire _0719_;
	wire _0720_;
	wire _0721_;
	wire _0722_;
	wire _0723_;
	wire _0724_;
	wire _0725_;
	wire _0726_;
	wire _0727_;
	wire _0728_;
	wire _0729_;
	wire _0730_;
	wire _0731_;
	wire _0732_;
	wire _0733_;
	wire _0734_;
	wire _0735_;
	wire _0736_;
	wire _0737_;
	wire _0738_;
	wire _0739_;
	wire _0740_;
	wire _0741_;
	wire _0742_;
	wire _0743_;
	wire _0744_;
	wire _0745_;
	wire _0746_;
	wire _0747_;
	wire _0748_;
	wire _0749_;
	wire _0750_;
	wire _0751_;
	wire _0752_;
	wire _0753_;
	wire _0754_;
	wire _0755_;
	wire _0756_;
	wire _0757_;
	wire _0758_;
	wire _0759_;
	wire _0760_;
	wire _0761_;
	wire _0762_;
	wire _0763_;
	wire _0764_;
	wire _0765_;
	wire _0766_;
	wire _0767_;
	wire _0768_;
	wire _0769_;
	wire _0770_;
	wire _0771_;
	wire _0772_;
	wire _0773_;
	wire _0774_;
	wire _0775_;
	wire _0776_;
	wire _0777_;
	wire _0778_;
	wire _0779_;
	wire _0780_;
	wire _0781_;
	wire _0782_;
	wire _0783_;
	wire _0784_;
	wire _0785_;
	wire _0786_;
	wire _0787_;
	wire _0788_;
	wire _0789_;
	wire _0790_;
	wire _0791_;
	wire _0792_;
	wire _0793_;
	wire _0794_;
	wire _0795_;
	wire _0796_;
	wire _0797_;
	wire _0798_;
	wire _0799_;
	wire _0800_;
	wire _0801_;
	wire _0802_;
	wire _0803_;
	wire _0804_;
	wire _0805_;
	wire _0806_;
	wire _0807_;
	wire _0808_;
	wire [5:0] _0809_;
	input wire [13:0] io_in;
	output wire [13:0] io_out;
	wire [15:0] \mchip.addr ;
	reg [15:0] \mchip.addr_cache ;
	reg [7:0] \mchip.bf.acc ;
	wire [15:0] \mchip.bf.addr ;
	wire [2:0] \mchip.bf.bus_op ;
	wire \mchip.bf.clock ;
	reg [15:0] \mchip.bf.cursor ;
	reg [11:0] \mchip.bf.depth ;
	wire \mchip.bf.enable ;
	wire \mchip.bf.halted ;
	wire [7:0] \mchip.bf.next_acc ;
	wire [15:0] \mchip.bf.next_cursor ;
	wire [11:0] \mchip.bf.next_depth ;
	wire [15:0] \mchip.bf.next_pc ;
	reg [15:0] \mchip.bf.pc ;
	wire \mchip.bf.reset ;
	reg [5:0] \mchip.bf.state ;
	wire [13:0] \mchip.bf.ucode ;
	wire [7:0] \mchip.bf.val_in ;
	wire [7:0] \mchip.bf.val_out ;
	wire [7:0] \mchip.bus_in ;
	wire [2:0] \mchip.bus_op ;
	wire [7:0] \mchip.bus_out ;
	wire \mchip.clock ;
	wire \mchip.enable ;
	wire \mchip.halted ;
	wire [11:0] \mchip.io_in ;
	wire [11:0] \mchip.io_out ;
	wire [2:0] \mchip.next_state ;
	reg [2:0] \mchip.op_cache ;
	wire \mchip.op_done ;
	wire \mchip.reset ;
	reg [2:0] \mchip.state ;
	reg [7:0] \mchip.val_cache ;
	reg [7:0] \mchip.val_in ;
	wire [7:0] \mchip.val_out ;
	assign _0085_ = \mchip.state [0] | \mchip.state [1];
	assign _0086_ = _0085_ | \mchip.state [2];
	assign \mchip.bf.enable  = io_in[9] & ~_0086_;
	assign \mchip.bf.next_pc [0] = ~\mchip.bf.pc [0];
	assign \mchip.bf.next_cursor [0] = ~\mchip.bf.cursor [0];
	assign _0087_ = \mchip.bf.state [0] | ~\mchip.bf.state [1];
	assign _0088_ = \mchip.bf.state [3] | \mchip.bf.state [2];
	assign _0089_ = ~(_0088_ | _0087_);
	assign _0090_ = ~(\mchip.bf.state [5] | \mchip.bf.state [4]);
	assign \mchip.bf.halted  = _0090_ & _0089_;
	assign _0091_ = \mchip.bf.state [4] & ~\mchip.bf.state [5];
	assign _0092_ = \mchip.bf.state [2] | ~\mchip.bf.state [3];
	assign _0093_ = \mchip.bf.state [1] | ~\mchip.bf.state [0];
	assign _0094_ = _0093_ | _0092_;
	assign _0095_ = _0091_ & ~_0094_;
	assign _0096_ = _0092_ | _0087_;
	assign _0097_ = _0091_ & ~_0096_;
	assign _0098_ = _0097_ | _0095_;
	assign _0099_ = ~(\mchip.bf.state [0] & \mchip.bf.state [1]);
	assign _0100_ = _0099_ | _0092_;
	assign _0101_ = _0091_ & ~_0100_;
	assign _0102_ = ~(_0101_ | _0098_);
	assign _0103_ = \mchip.bf.state [0] | \mchip.bf.state [1];
	assign _0104_ = _0103_ | _0088_;
	assign _0105_ = _0090_ & ~_0104_;
	assign _0106_ = ~_0105_;
	assign _0107_ = \mchip.bf.state [3] | ~\mchip.bf.state [2];
	assign _0108_ = _0107_ | _0093_;
	assign _0109_ = _0090_ & ~_0108_;
	assign _0110_ = _0103_ | _0092_;
	assign _0111_ = _0090_ & ~_0110_;
	assign _0112_ = _0111_ | _0109_;
	assign _0113_ = _0090_ & ~_0094_;
	assign _0114_ = _0090_ & ~_0096_;
	assign _0115_ = _0114_ | _0113_;
	assign _0116_ = _0115_ | _0112_;
	assign _0117_ = ~(\mchip.bf.state [3] & \mchip.bf.state [2]);
	assign _0118_ = _0117_ | _0093_;
	assign _0119_ = _0090_ & ~_0118_;
	assign _0120_ = _0117_ | _0087_;
	assign _0121_ = _0090_ & ~_0120_;
	assign _0122_ = _0121_ | _0119_;
	assign _0123_ = _0117_ | _0099_;
	assign _0124_ = _0090_ & ~_0123_;
	assign _0125_ = _0107_ | _0099_;
	assign _0126_ = _0090_ & ~_0125_;
	assign _0127_ = _0126_ | _0124_;
	assign _0128_ = _0117_ | _0103_;
	assign _0129_ = _0090_ & ~_0128_;
	assign _0130_ = _0107_ | _0103_;
	assign _0131_ = _0090_ & ~_0130_;
	assign _0132_ = _0131_ | _0129_;
	assign _0133_ = _0132_ | _0127_;
	assign _0134_ = _0091_ & ~_0104_;
	assign _0135_ = _0134_ | _0133_;
	assign _0136_ = _0135_ | _0122_;
	assign _0137_ = _0136_ | _0116_;
	assign _0138_ = _0091_ & ~_0125_;
	assign _0139_ = _0090_ & ~_0100_;
	assign _0140_ = _0099_ | _0088_;
	assign _0141_ = _0090_ & ~_0140_;
	assign _0142_ = _0141_ | _0139_;
	assign _0143_ = _0093_ | _0088_;
	assign _0144_ = _0091_ & ~_0143_;
	assign _0145_ = _0107_ | _0087_;
	assign _0146_ = _0090_ & ~_0145_;
	assign _0147_ = _0146_ | _0144_;
	assign _0148_ = _0147_ | _0142_;
	assign _0149_ = _0148_ | _0138_;
	assign _0150_ = _0091_ & ~_0140_;
	assign _0151_ = _0150_ | _0149_;
	assign _0152_ = _0090_ & ~_0143_;
	assign _0153_ = _0091_ & _0089_;
	assign _0154_ = _0153_ | _0152_;
	assign _0155_ = _0091_ & ~_0110_;
	assign _0156_ = _0155_ | \mchip.bf.halted ;
	assign _0157_ = _0156_ | _0154_;
	assign _0158_ = _0157_ | _0098_;
	assign _0159_ = _0158_ | _0151_;
	assign _0160_ = _0091_ & ~_0118_;
	assign _0161_ = _0091_ & ~_0108_;
	assign _0162_ = _0161_ | _0160_;
	assign _0163_ = _0162_ | _0101_;
	assign _0164_ = _0091_ & ~_0120_;
	assign _0165_ = _0091_ & ~_0145_;
	assign _0166_ = _0165_ | _0164_;
	assign _0167_ = _0091_ & ~_0123_;
	assign _0168_ = \mchip.bf.state [4] | ~\mchip.bf.state [5];
	assign _0169_ = ~(_0168_ | _0104_);
	assign _0170_ = _0169_ | _0167_;
	assign _0171_ = _0170_ | _0166_;
	assign _0172_ = _0171_ | _0163_;
	assign _0173_ = _0172_ | _0159_;
	assign _0174_ = _0173_ | _0137_;
	assign _0175_ = _0106_ & ~_0174_;
	assign _0176_ = _0175_ | _0102_;
	assign _0177_ = _0170_ | _0150_;
	assign _0178_ = _0106_ & ~_0177_;
	assign _0179_ = ~(_0178_ | _0175_);
	assign _0180_ = _0179_ ^ _0176_;
	assign _0002_ = \mchip.bf.enable  & ~_0180_;
	assign _0181_ = _0175_ | ~_0114_;
	assign _0182_ = _0113_ & ~_0175_;
	assign _0183_ = _0182_ ^ _0181_;
	assign _0003_ = \mchip.bf.enable  & ~_0183_;
	assign _0184_ = \mchip.state [2] & ~_0085_;
	assign _0004_ = _0184_ & io_in[9];
	assign _0185_ = _0175_ | ~_0133_;
	assign _0001_ = \mchip.bf.enable  & ~_0185_;
	assign _0186_ = ~(_0166_ | _0162_);
	assign _0187_ = _0186_ | _0175_;
	assign _0188_ = _0158_ | _0149_;
	assign _0189_ = _0188_ | _0171_;
	assign _0190_ = _0189_ | _0137_;
	assign _0191_ = _0106_ & ~_0190_;
	assign _0192_ = ~(_0191_ | _0175_);
	assign _0193_ = _0187_ & ~_0192_;
	assign _0000_ = \mchip.bf.enable  & ~_0193_;
	assign _0194_ = _0134_ | _0119_;
	assign _0195_ = ~(_0194_ | _0112_);
	assign \mchip.bf.ucode [11] = ~(_0195_ | _0175_);
	assign _0196_ = _0150_ | _0101_;
	assign _0197_ = _0196_ | _0122_;
	assign _0198_ = _0106_ & ~_0197_;
	assign \mchip.bf.ucode [12] = ~(_0198_ | _0175_);
	assign _0199_ = _0134_ | _0122_;
	assign _0200_ = ~(_0199_ | _0112_);
	assign _0201_ = _0200_ & ~_0149_;
	assign \mchip.bf.ucode [13] = ~(_0201_ | _0175_);
	assign _0202_ = ~(_0186_ | _0175_);
	assign \mchip.bf.next_depth [0] = _0202_ & ~\mchip.bf.depth [0];
	assign _0203_ = ~\mchip.bf.depth [1];
	assign _0204_ = _0192_ & ~_0187_;
	assign _0205_ = _0204_ ^ _0203_;
	assign _0206_ = _0205_ ^ \mchip.bf.depth [0];
	assign \mchip.bf.next_depth [1] = _0202_ & ~_0206_;
	assign _0207_ = _0204_ & ~_0203_;
	assign _0208_ = \mchip.bf.depth [0] & ~_0205_;
	assign _0209_ = _0208_ | _0207_;
	assign _0210_ = ~\mchip.bf.depth [2];
	assign _0211_ = _0204_ ^ _0210_;
	assign _0212_ = _0211_ ^ _0209_;
	assign \mchip.bf.next_depth [2] = _0202_ & ~_0212_;
	assign _0213_ = _0204_ & ~_0210_;
	assign _0214_ = _0209_ & ~_0211_;
	assign _0215_ = _0214_ | _0213_;
	assign _0216_ = ~\mchip.bf.depth [3];
	assign _0217_ = _0204_ ^ _0216_;
	assign _0218_ = _0217_ ^ _0215_;
	assign \mchip.bf.next_depth [3] = _0202_ & ~_0218_;
	assign _0219_ = _0217_ | _0211_;
	assign _0220_ = _0209_ & ~_0219_;
	assign _0221_ = _0213_ & ~_0217_;
	assign _0222_ = _0204_ & ~_0216_;
	assign _0223_ = _0222_ | _0221_;
	assign _0224_ = _0223_ | _0220_;
	assign _0225_ = ~\mchip.bf.depth [4];
	assign _0226_ = _0204_ ^ _0225_;
	assign _0227_ = _0226_ ^ _0224_;
	assign \mchip.bf.next_depth [4] = _0202_ & ~_0227_;
	assign _0228_ = _0204_ & ~_0225_;
	assign _0229_ = _0224_ & ~_0226_;
	assign _0230_ = _0229_ | _0228_;
	assign _0231_ = ~\mchip.bf.depth [5];
	assign _0232_ = _0204_ ^ _0231_;
	assign _0233_ = _0232_ ^ _0230_;
	assign \mchip.bf.next_depth [5] = _0202_ & ~_0233_;
	assign _0234_ = _0232_ | _0226_;
	assign _0235_ = _0224_ & ~_0234_;
	assign _0236_ = _0228_ & ~_0232_;
	assign _0237_ = _0204_ & ~_0231_;
	assign _0238_ = _0237_ | _0236_;
	assign _0239_ = _0238_ | _0235_;
	assign _0240_ = ~\mchip.bf.depth [6];
	assign _0241_ = _0204_ ^ _0240_;
	assign _0242_ = _0241_ ^ _0239_;
	assign \mchip.bf.next_depth [6] = _0202_ & ~_0242_;
	assign _0243_ = _0204_ & ~_0240_;
	assign _0244_ = _0239_ & ~_0241_;
	assign _0245_ = _0244_ | _0243_;
	assign _0246_ = ~\mchip.bf.depth [7];
	assign _0247_ = _0204_ ^ _0246_;
	assign _0248_ = _0247_ ^ _0245_;
	assign \mchip.bf.next_depth [7] = _0202_ & ~_0248_;
	assign _0249_ = _0204_ & ~_0246_;
	assign _0250_ = _0243_ & ~_0247_;
	assign _0251_ = _0250_ | _0249_;
	assign _0252_ = _0247_ | _0241_;
	assign _0253_ = _0238_ & ~_0252_;
	assign _0254_ = _0253_ | _0251_;
	assign _0255_ = _0252_ | _0234_;
	assign _0256_ = _0224_ & ~_0255_;
	assign _0257_ = _0256_ | _0254_;
	assign _0258_ = ~\mchip.bf.depth [8];
	assign _0259_ = _0204_ ^ _0258_;
	assign _0260_ = _0259_ ^ _0257_;
	assign \mchip.bf.next_depth [8] = _0202_ & ~_0260_;
	assign _0261_ = _0204_ & ~_0258_;
	assign _0262_ = _0259_ | ~_0257_;
	assign _0263_ = _0262_ & ~_0261_;
	assign _0264_ = _0204_ ^ \mchip.bf.depth [9];
	assign _0265_ = _0264_ ^ _0263_;
	assign \mchip.bf.next_depth [9] = _0202_ & ~_0265_;
	assign _0266_ = ~(_0204_ & \mchip.bf.depth [9]);
	assign _0267_ = ~(_0264_ & _0261_);
	assign _0268_ = ~(_0267_ & _0266_);
	assign _0269_ = _0259_ | ~_0264_;
	assign _0270_ = _0257_ & ~_0269_;
	assign _0271_ = _0270_ | _0268_;
	assign _0272_ = ~\mchip.bf.depth [10];
	assign _0273_ = _0204_ ^ _0272_;
	assign _0274_ = _0273_ ^ _0271_;
	assign \mchip.bf.next_depth [10] = _0202_ & ~_0274_;
	assign _0275_ = _0271_ & ~_0273_;
	assign _0276_ = _0204_ & ~_0272_;
	assign _0277_ = _0276_ | _0275_;
	assign _0278_ = ~(_0204_ ^ \mchip.bf.depth [11]);
	assign _0279_ = _0278_ ^ _0277_;
	assign \mchip.bf.next_depth [11] = _0202_ & ~_0279_;
	assign _0280_ = _0091_ & ~_0128_;
	assign _0281_ = \mchip.val_in [7] | ~\mchip.val_in [6];
	assign _0282_ = \mchip.val_in [5] | ~\mchip.val_in [4];
	assign _0283_ = _0282_ | _0281_;
	assign _0284_ = \mchip.val_in [2] | ~\mchip.val_in [3];
	assign _0285_ = ~(\mchip.val_in [0] & \mchip.val_in [1]);
	assign _0286_ = _0285_ | _0284_;
	assign _0287_ = _0286_ | _0283_;
	assign _0288_ = ~(\mchip.bf.depth [1] | \mchip.bf.depth [0]);
	assign _0289_ = \mchip.bf.depth [3] | \mchip.bf.depth [2];
	assign _0290_ = _0288_ & ~_0289_;
	assign _0291_ = \mchip.bf.depth [7] | \mchip.bf.depth [6];
	assign _0292_ = \mchip.bf.depth [5] | \mchip.bf.depth [4];
	assign _0293_ = _0292_ | _0291_;
	assign _0294_ = _0290_ & ~_0293_;
	assign _0295_ = \mchip.bf.depth [11] | \mchip.bf.depth [10];
	assign _0296_ = \mchip.bf.depth [9] | \mchip.bf.depth [8];
	assign _0297_ = _0296_ | _0295_;
	assign _0298_ = _0294_ & ~_0297_;
	assign _0299_ = _0287_ | ~_0298_;
	assign _0300_ = \mchip.bf.enable  & ~io_in[13];
	assign _0301_ = ~_0300_;
	assign _0302_ = _0301_ | _0299_;
	assign _0303_ = _0280_ & ~_0302_;
	assign _0304_ = ~(\mchip.bf.enable  | io_in[13]);
	assign _0305_ = _0304_ & _0167_;
	assign _0306_ = _0305_ | _0303_;
	assign _0307_ = _0300_ & _0121_;
	assign _0308_ = _0304_ & _0124_;
	assign _0309_ = _0308_ | _0307_;
	assign _0310_ = _0309_ | _0306_;
	assign _0311_ = \mchip.val_in [1] | ~\mchip.val_in [0];
	assign _0312_ = ~(\mchip.val_in [3] & \mchip.val_in [2]);
	assign _0313_ = _0312_ | _0311_;
	assign _0314_ = _0313_ | _0283_;
	assign _0315_ = _0314_ | ~_0300_;
	assign _0316_ = _0152_ & ~_0315_;
	assign _0317_ = _0304_ & _0138_;
	assign _0318_ = _0317_ | _0316_;
	assign _0319_ = _0300_ & _0146_;
	assign _0320_ = _0304_ & _0126_;
	assign _0321_ = _0320_ | _0319_;
	assign _0322_ = _0321_ | _0318_;
	assign _0323_ = _0322_ | _0310_;
	assign _0324_ = ~(_0165_ | _0161_);
	assign _0325_ = _0324_ & _0300_;
	assign _0326_ = ~(_0164_ | _0097_);
	assign _0327_ = _0326_ & ~_0160_;
	assign _0328_ = _0325_ & ~_0327_;
	assign _0329_ = ~(\mchip.val_in [3] | \mchip.val_in [2]);
	assign _0330_ = \mchip.val_in [0] | \mchip.val_in [1];
	assign _0331_ = _0329_ & ~_0330_;
	assign _0332_ = \mchip.val_in [4] | \mchip.val_in [5];
	assign _0333_ = \mchip.val_in [6] | \mchip.val_in [7];
	assign _0334_ = _0333_ | _0332_;
	assign _0335_ = _0331_ & ~_0334_;
	assign _0336_ = _0287_ & ~_0335_;
	assign _0337_ = ~(_0336_ & _0300_);
	assign _0338_ = _0337_ | ~_0314_;
	assign _0339_ = _0280_ & ~_0338_;
	assign _0340_ = _0304_ & _0101_;
	assign _0341_ = _0340_ | _0339_;
	assign _0342_ = _0341_ | _0328_;
	assign _0343_ = \mchip.val_in [4] | ~\mchip.val_in [5];
	assign _0344_ = _0343_ | _0333_;
	assign _0345_ = \mchip.val_in [0] | ~\mchip.val_in [1];
	assign _0346_ = _0345_ | _0312_;
	assign _0347_ = ~(_0346_ | _0344_);
	assign _0348_ = ~(_0347_ & _0300_);
	assign _0349_ = _0152_ & ~_0348_;
	assign _0350_ = _0304_ & _0139_;
	assign _0351_ = _0350_ | _0349_;
	assign _0352_ = _0351_ | _0342_;
	assign _0353_ = _0300_ & ~_0324_;
	assign _0354_ = _0335_ & _0300_;
	assign _0355_ = _0354_ & _0153_;
	assign _0356_ = _0355_ | _0353_;
	assign _0357_ = _0091_ & ~_0130_;
	assign _0358_ = _0357_ & ~_0338_;
	assign _0359_ = _0304_ & _0150_;
	assign _0360_ = _0359_ | _0358_;
	assign _0361_ = _0360_ | _0356_;
	assign _0362_ = ~(_0344_ | _0286_);
	assign _0363_ = ~(_0362_ & _0300_);
	assign _0364_ = _0152_ & ~_0363_;
	assign _0365_ = _0304_ & _0141_;
	assign _0366_ = _0365_ | _0364_;
	assign _0367_ = _0366_ | _0361_;
	assign _0368_ = _0367_ | _0352_;
	assign _0369_ = ~(_0368_ | _0323_);
	assign _0370_ = _0280_ & ~_0315_;
	assign _0371_ = _0304_ & _0160_;
	assign _0372_ = _0371_ | _0370_;
	assign _0373_ = _0304_ & _0119_;
	assign _0374_ = _0300_ & _0129_;
	assign _0375_ = _0374_ | _0373_;
	assign _0376_ = _0375_ | _0372_;
	assign _0377_ = _0304_ & _0161_;
	assign _0378_ = _0287_ | ~_0300_;
	assign _0379_ = _0357_ & ~_0378_;
	assign _0380_ = _0379_ | _0377_;
	assign _0381_ = _0304_ & _0109_;
	assign _0382_ = _0300_ & _0131_;
	assign _0383_ = _0382_ | _0381_;
	assign _0384_ = _0383_ | _0380_;
	assign _0385_ = _0384_ | _0376_;
	assign _0386_ = _0304_ & _0095_;
	assign _0387_ = _0335_ | ~_0300_;
	assign _0388_ = _0155_ & ~_0387_;
	assign _0389_ = _0388_ | _0386_;
	assign _0390_ = _0304_ & _0113_;
	assign _0391_ = ~(\mchip.val_in [4] & \mchip.val_in [5]);
	assign _0392_ = _0391_ | _0333_;
	assign _0393_ = ~(_0392_ | _0346_);
	assign _0394_ = ~(_0393_ & _0300_);
	assign _0395_ = _0152_ & ~_0394_;
	assign _0396_ = _0395_ | _0390_;
	assign _0397_ = _0396_ | _0389_;
	assign _0398_ = _0304_ & _0144_;
	assign _0399_ = _0152_ & ~_0378_;
	assign _0400_ = _0399_ | _0398_;
	assign _0401_ = _0304_ & _0152_;
	assign _0402_ = _0300_ & ~_0106_;
	assign _0403_ = _0402_ | _0401_;
	assign _0404_ = _0403_ | _0400_;
	assign _0405_ = _0404_ | _0397_;
	assign _0406_ = _0405_ | _0385_;
	assign _0809_[0] = _0406_ | ~_0369_;
	assign _0407_ = _0304_ & _0164_;
	assign _0408_ = _0298_ | _0287_;
	assign _0409_ = _0408_ | _0301_;
	assign _0410_ = _0280_ & ~_0409_;
	assign _0411_ = _0410_ | _0407_;
	assign _0412_ = _0304_ & _0121_;
	assign _0413_ = _0330_ | _0312_;
	assign _0414_ = ~(_0413_ | _0344_);
	assign _0415_ = ~(_0414_ & _0300_);
	assign _0416_ = _0152_ & ~_0415_;
	assign _0417_ = _0416_ | _0412_;
	assign _0418_ = _0417_ | _0411_;
	assign _0419_ = _0304_ & _0165_;
	assign _0420_ = _0314_ | _0298_;
	assign _0421_ = _0420_ | _0301_;
	assign _0422_ = _0357_ & ~_0421_;
	assign _0423_ = _0422_ | _0419_;
	assign _0424_ = _0304_ & _0146_;
	assign _0425_ = ~(_0344_ | _0313_);
	assign _0426_ = ~(_0425_ & _0300_);
	assign _0427_ = _0152_ & ~_0426_;
	assign _0428_ = _0427_ | _0424_;
	assign _0429_ = _0428_ | _0423_;
	assign _0430_ = ~(_0429_ | _0418_);
	assign _0431_ = _0304_ & _0097_;
	assign _0432_ = _0300_ & _0095_;
	assign _0433_ = _0432_ | _0431_;
	assign _0434_ = ~(_0413_ | _0392_);
	assign _0435_ = ~(_0434_ & _0300_);
	assign _0436_ = _0152_ & ~_0435_;
	assign _0437_ = _0304_ & _0114_;
	assign _0438_ = _0437_ | _0436_;
	assign _0439_ = _0438_ | _0433_;
	assign _0440_ = _0304_ & _0153_;
	assign _0441_ = _0300_ & _0144_;
	assign _0442_ = _0441_ | _0440_;
	assign _0443_ = _0357_ | _0280_;
	assign _0444_ = ~(_0443_ | _0152_);
	assign _0445_ = _0354_ & ~_0444_;
	assign _0446_ = \mchip.bf.halted  & ~io_in[13];
	assign _0447_ = _0446_ | _0445_;
	assign _0448_ = _0447_ | _0442_;
	assign _0449_ = ~(_0448_ | _0439_);
	assign _0450_ = ~(_0449_ & _0430_);
	assign _0451_ = _0304_ & _0131_;
	assign _0452_ = _0300_ & _0141_;
	assign _0453_ = _0452_ | _0451_;
	assign _0454_ = _0300_ & _0150_;
	assign _0455_ = _0357_ & _0304_;
	assign _0456_ = _0455_ | _0454_;
	assign _0457_ = ~(_0456_ | _0453_);
	assign _0458_ = _0304_ & _0280_;
	assign _0459_ = _0300_ & _0101_;
	assign _0460_ = _0459_ | _0458_;
	assign _0461_ = _0300_ & _0139_;
	assign _0462_ = _0304_ & _0129_;
	assign _0463_ = _0462_ | _0461_;
	assign _0464_ = ~(_0463_ | _0460_);
	assign _0465_ = ~(_0464_ & _0457_);
	assign _0466_ = _0304_ & _0134_;
	assign _0467_ = _0300_ & _0124_;
	assign _0468_ = ~(_0467_ | _0466_);
	assign _0469_ = _0304_ & _0169_;
	assign _0470_ = _0300_ & _0167_;
	assign _0471_ = _0470_ | _0469_;
	assign _0472_ = _0471_ | ~_0468_;
	assign _0473_ = _0300_ & _0138_;
	assign _0474_ = _0304_ & _0155_;
	assign _0475_ = _0474_ | _0473_;
	assign _0476_ = _0304_ & _0111_;
	assign _0477_ = _0300_ & _0126_;
	assign _0478_ = _0477_ | _0476_;
	assign _0479_ = _0478_ | _0475_;
	assign _0480_ = _0479_ | _0472_;
	assign _0481_ = _0480_ | _0465_;
	assign _0482_ = _0481_ | _0450_;
	assign _0483_ = _0482_ | _0809_[0];
	assign _0484_ = _0369_ & ~_0450_;
	assign _0809_[1] = _0483_ & ~_0484_;
	assign _0485_ = _0430_ & ~_0465_;
	assign _0486_ = _0385_ | _0323_;
	assign _0487_ = _0485_ & ~_0486_;
	assign _0809_[2] = _0483_ & ~_0487_;
	assign _0488_ = _0464_ & ~_0479_;
	assign _0489_ = _0439_ | _0418_;
	assign _0490_ = _0488_ & ~_0489_;
	assign _0491_ = _0352_ | _0310_;
	assign _0492_ = _0397_ | _0376_;
	assign _0493_ = _0492_ | _0491_;
	assign _0494_ = _0490_ & ~_0493_;
	assign _0809_[3] = _0483_ & ~_0494_;
	assign _0495_ = _0468_ & ~_0475_;
	assign _0496_ = _0460_ | _0456_;
	assign _0497_ = _0495_ & ~_0496_;
	assign _0498_ = _0423_ | _0411_;
	assign _0499_ = _0442_ | _0433_;
	assign _0500_ = _0499_ | _0498_;
	assign _0501_ = _0497_ & ~_0500_;
	assign _0502_ = _0318_ | _0306_;
	assign _0503_ = _0361_ | _0342_;
	assign _0504_ = _0503_ | _0502_;
	assign _0505_ = _0380_ | _0372_;
	assign _0506_ = _0400_ | _0389_;
	assign _0507_ = _0506_ | _0505_;
	assign _0508_ = _0507_ | _0504_;
	assign _0509_ = _0501_ & ~_0508_;
	assign _0809_[4] = _0483_ & ~_0509_;
	assign _0809_[5] = _0483_ & _0471_;
	assign _0510_ = _0175_ | ~_0112_;
	assign _0511_ = ~_0510_;
	assign _0512_ = ~(_0194_ | _0111_);
	assign _0513_ = _0512_ | _0175_;
	assign _0514_ = _0510_ & ~_0513_;
	assign \mchip.val_out [0] = (\mchip.bf.acc [0] ? _0514_ : _0511_);
	assign _0515_ = ~(_0513_ & _0510_);
	assign _0516_ = ~\mchip.bf.acc [1];
	assign _0517_ = ~(_0513_ | _0510_);
	assign _0518_ = _0517_ ^ _0516_;
	assign _0519_ = _0518_ ^ \mchip.bf.acc [0];
	assign _0520_ = _0519_ | _0510_;
	assign _0521_ = _0514_ & ~_0516_;
	assign _0522_ = _0520_ & ~_0521_;
	assign \mchip.val_out [1] = _0515_ & ~_0522_;
	assign _0523_ = _0517_ & ~_0516_;
	assign _0524_ = \mchip.bf.acc [0] & ~_0518_;
	assign _0525_ = _0524_ | _0523_;
	assign _0526_ = ~\mchip.bf.acc [2];
	assign _0527_ = _0517_ ^ _0526_;
	assign _0528_ = _0527_ ^ _0525_;
	assign _0529_ = _0528_ | _0510_;
	assign _0530_ = _0514_ & ~_0526_;
	assign _0531_ = _0529_ & ~_0530_;
	assign \mchip.val_out [2] = _0515_ & ~_0531_;
	assign _0532_ = _0517_ & ~_0526_;
	assign _0533_ = _0525_ & ~_0527_;
	assign _0534_ = _0533_ | _0532_;
	assign _0535_ = ~\mchip.bf.acc [3];
	assign _0536_ = _0517_ ^ _0535_;
	assign _0537_ = _0536_ ^ _0534_;
	assign _0538_ = _0537_ | _0510_;
	assign _0539_ = _0514_ & ~_0535_;
	assign _0540_ = _0538_ & ~_0539_;
	assign \mchip.val_out [3] = _0515_ & ~_0540_;
	assign _0541_ = _0517_ & ~_0535_;
	assign _0542_ = _0532_ & ~_0536_;
	assign _0543_ = _0542_ | _0541_;
	assign _0544_ = _0536_ | _0527_;
	assign _0545_ = _0525_ & ~_0544_;
	assign _0546_ = _0545_ | _0543_;
	assign _0547_ = ~\mchip.bf.acc [4];
	assign _0548_ = _0517_ ^ _0547_;
	assign _0549_ = _0548_ ^ _0546_;
	assign _0550_ = _0549_ | _0510_;
	assign _0551_ = _0514_ & ~_0547_;
	assign _0552_ = _0550_ & ~_0551_;
	assign \mchip.val_out [4] = _0515_ & ~_0552_;
	assign _0553_ = _0517_ & ~_0547_;
	assign _0554_ = _0546_ & ~_0548_;
	assign _0555_ = _0554_ | _0553_;
	assign _0556_ = ~\mchip.bf.acc [5];
	assign _0557_ = _0517_ ^ _0556_;
	assign _0558_ = _0557_ ^ _0555_;
	assign _0559_ = _0558_ | _0510_;
	assign _0560_ = _0514_ & ~_0556_;
	assign _0561_ = _0559_ & ~_0560_;
	assign \mchip.val_out [5] = _0515_ & ~_0561_;
	assign _0562_ = _0517_ & ~_0556_;
	assign _0563_ = _0553_ & ~_0557_;
	assign _0564_ = _0563_ | _0562_;
	assign _0565_ = _0557_ | _0548_;
	assign _0566_ = _0546_ & ~_0565_;
	assign _0567_ = _0566_ | _0564_;
	assign _0568_ = ~\mchip.bf.acc [6];
	assign _0569_ = _0517_ ^ _0568_;
	assign _0570_ = _0569_ ^ _0567_;
	assign _0571_ = _0570_ | _0510_;
	assign _0572_ = _0514_ & ~_0568_;
	assign _0573_ = _0571_ & ~_0572_;
	assign \mchip.val_out [6] = _0515_ & ~_0573_;
	assign _0574_ = _0567_ & ~_0569_;
	assign _0575_ = _0517_ & ~_0568_;
	assign _0576_ = _0575_ | _0574_;
	assign _0577_ = ~(_0517_ ^ \mchip.bf.acc [7]);
	assign _0578_ = _0577_ ^ _0576_;
	assign _0579_ = _0578_ | _0510_;
	assign _0580_ = _0514_ & \mchip.bf.acc [7];
	assign _0581_ = _0579_ & ~_0580_;
	assign \mchip.val_out [7] = _0515_ & ~_0581_;
	assign _0582_ = ~(_0134_ | _0112_);
	assign _0583_ = _0582_ & ~_0149_;
	assign _0584_ = ~(_0583_ | _0175_);
	assign _0585_ = _0106_ & ~_0196_;
	assign _0586_ = ~(_0585_ | _0175_);
	assign _0587_ = _0584_ | ~_0586_;
	assign _0588_ = _0586_ | ~_0584_;
	assign _0589_ = ~(_0588_ & _0587_);
	assign _0590_ = _0587_ | \mchip.bf.next_pc [0];
	assign _0591_ = \mchip.bf.cursor [0] & ~_0588_;
	assign _0592_ = _0590_ & ~_0591_;
	assign \mchip.addr [0] = _0589_ & ~_0592_;
	assign _0593_ = ~\mchip.bf.cursor [1];
	assign _0594_ = _0588_ | _0593_;
	assign _0595_ = \mchip.bf.pc [1] & ~_0587_;
	assign _0596_ = _0594_ & ~_0595_;
	assign \mchip.addr [1] = _0589_ & ~_0596_;
	assign _0597_ = ~\mchip.bf.cursor [2];
	assign _0598_ = _0588_ | _0597_;
	assign _0599_ = \mchip.bf.pc [2] & ~_0587_;
	assign _0600_ = _0598_ & ~_0599_;
	assign \mchip.addr [2] = _0589_ & ~_0600_;
	assign _0601_ = ~\mchip.bf.cursor [3];
	assign _0602_ = _0588_ | _0601_;
	assign _0603_ = \mchip.bf.pc [3] & ~_0587_;
	assign _0604_ = _0602_ & ~_0603_;
	assign \mchip.addr [3] = _0589_ & ~_0604_;
	assign _0605_ = ~\mchip.bf.cursor [4];
	assign _0606_ = _0588_ | _0605_;
	assign _0607_ = \mchip.bf.pc [4] & ~_0587_;
	assign _0608_ = _0606_ & ~_0607_;
	assign \mchip.addr [4] = _0589_ & ~_0608_;
	assign _0609_ = ~\mchip.bf.cursor [5];
	assign _0610_ = _0588_ | _0609_;
	assign _0611_ = \mchip.bf.pc [5] & ~_0587_;
	assign _0612_ = _0610_ & ~_0611_;
	assign \mchip.addr [5] = _0589_ & ~_0612_;
	assign _0613_ = ~\mchip.bf.cursor [6];
	assign _0614_ = _0588_ | _0613_;
	assign _0615_ = \mchip.bf.pc [6] & ~_0587_;
	assign _0616_ = _0614_ & ~_0615_;
	assign \mchip.addr [6] = _0589_ & ~_0616_;
	assign _0617_ = ~\mchip.bf.cursor [7];
	assign _0618_ = _0588_ | _0617_;
	assign _0619_ = \mchip.bf.pc [7] & ~_0587_;
	assign _0620_ = _0618_ & ~_0619_;
	assign \mchip.addr [7] = _0589_ & ~_0620_;
	assign _0621_ = ~\mchip.bf.cursor [8];
	assign _0622_ = _0588_ | _0621_;
	assign _0623_ = \mchip.bf.pc [8] & ~_0587_;
	assign _0624_ = _0622_ & ~_0623_;
	assign \mchip.addr [8] = _0589_ & ~_0624_;
	assign _0625_ = ~\mchip.bf.cursor [9];
	assign _0626_ = _0588_ | _0625_;
	assign _0627_ = \mchip.bf.pc [9] & ~_0587_;
	assign _0628_ = _0626_ & ~_0627_;
	assign \mchip.addr [9] = _0589_ & ~_0628_;
	assign _0629_ = ~\mchip.bf.cursor [10];
	assign _0630_ = _0588_ | _0629_;
	assign _0631_ = \mchip.bf.pc [10] & ~_0587_;
	assign _0632_ = _0630_ & ~_0631_;
	assign \mchip.addr [10] = _0589_ & ~_0632_;
	assign _0633_ = ~\mchip.bf.cursor [11];
	assign _0634_ = _0588_ | _0633_;
	assign _0635_ = \mchip.bf.pc [11] & ~_0587_;
	assign _0636_ = _0634_ & ~_0635_;
	assign \mchip.addr [11] = _0589_ & ~_0636_;
	assign _0637_ = ~\mchip.bf.cursor [12];
	assign _0638_ = _0588_ | _0637_;
	assign _0639_ = \mchip.bf.pc [12] & ~_0587_;
	assign _0640_ = _0638_ & ~_0639_;
	assign \mchip.addr [12] = _0589_ & ~_0640_;
	assign _0641_ = ~\mchip.bf.cursor [13];
	assign _0642_ = _0588_ | _0641_;
	assign _0643_ = \mchip.bf.pc [13] & ~_0587_;
	assign _0644_ = _0642_ & ~_0643_;
	assign \mchip.addr [13] = _0589_ & ~_0644_;
	assign _0645_ = ~\mchip.bf.cursor [14];
	assign _0646_ = _0588_ | _0645_;
	assign _0647_ = \mchip.bf.pc [14] & ~_0587_;
	assign _0648_ = _0646_ & ~_0647_;
	assign \mchip.addr [14] = _0589_ & ~_0648_;
	assign _0649_ = _0588_ | ~\mchip.bf.cursor [15];
	assign _0650_ = \mchip.bf.pc [15] & ~_0587_;
	assign _0651_ = _0649_ & ~_0650_;
	assign \mchip.addr [15] = _0589_ & ~_0651_;
	assign _0652_ = \mchip.state [1] | ~\mchip.state [0];
	assign _0653_ = _0652_ | \mchip.state [2];
	assign _0654_ = \mchip.state [0] | ~\mchip.state [1];
	assign _0655_ = _0654_ | \mchip.state [2];
	assign _0656_ = ~(_0655_ & _0653_);
	assign _0657_ = ~(\mchip.state [0] & \mchip.state [1]);
	assign _0658_ = ~(_0657_ | \mchip.state [2]);
	assign _0659_ = _0658_ | _0184_;
	assign _0660_ = _0659_ | _0656_;
	assign _0661_ = _0653_ | ~\mchip.op_cache [0];
	assign _0662_ = \mchip.addr_cache [8] & ~_0655_;
	assign _0663_ = _0661_ & ~_0662_;
	assign _0664_ = _0658_ & \mchip.addr_cache [0];
	assign _0665_ = _0184_ & \mchip.val_cache [0];
	assign _0666_ = _0665_ | _0664_;
	assign _0667_ = _0663_ & ~_0666_;
	assign io_out[0] = _0660_ & ~_0667_;
	assign _0668_ = ~(_0184_ & \mchip.val_cache [1]);
	assign _0669_ = _0658_ & \mchip.addr_cache [1];
	assign _0670_ = _0668_ & ~_0669_;
	assign _0671_ = \mchip.op_cache [1] & ~_0653_;
	assign _0672_ = \mchip.addr_cache [9] & ~_0655_;
	assign _0673_ = _0672_ | _0671_;
	assign _0674_ = _0670_ & ~_0673_;
	assign io_out[1] = _0660_ & ~_0674_;
	assign _0675_ = ~(_0184_ & \mchip.val_cache [2]);
	assign _0676_ = _0658_ & \mchip.addr_cache [2];
	assign _0677_ = _0675_ & ~_0676_;
	assign _0678_ = \mchip.op_cache [2] & ~_0653_;
	assign _0679_ = \mchip.addr_cache [10] & ~_0655_;
	assign _0680_ = _0679_ | _0678_;
	assign _0681_ = _0677_ & ~_0680_;
	assign io_out[2] = _0660_ & ~_0681_;
	assign _0682_ = ~(_0184_ & \mchip.val_cache [3]);
	assign _0683_ = _0658_ & \mchip.addr_cache [3];
	assign _0684_ = _0682_ & ~_0683_;
	assign _0685_ = \mchip.addr_cache [11] & ~_0655_;
	assign _0686_ = _0684_ & ~_0685_;
	assign io_out[3] = _0660_ & ~_0686_;
	assign _0687_ = ~(_0184_ & \mchip.val_cache [4]);
	assign _0688_ = _0658_ & \mchip.addr_cache [4];
	assign _0689_ = _0687_ & ~_0688_;
	assign _0690_ = \mchip.addr_cache [12] & ~_0655_;
	assign _0691_ = _0689_ & ~_0690_;
	assign io_out[4] = _0660_ & ~_0691_;
	assign _0692_ = ~(_0184_ & \mchip.val_cache [5]);
	assign _0693_ = _0658_ & \mchip.addr_cache [5];
	assign _0694_ = _0692_ & ~_0693_;
	assign _0695_ = \mchip.addr_cache [13] & ~_0655_;
	assign _0696_ = _0694_ & ~_0695_;
	assign io_out[5] = _0660_ & ~_0696_;
	assign _0697_ = ~(_0184_ & \mchip.val_cache [6]);
	assign _0698_ = _0658_ & \mchip.addr_cache [6];
	assign _0699_ = _0697_ & ~_0698_;
	assign _0700_ = \mchip.addr_cache [14] & ~_0655_;
	assign _0701_ = _0699_ & ~_0700_;
	assign io_out[6] = _0660_ & ~_0701_;
	assign _0702_ = ~(_0184_ & \mchip.val_cache [7]);
	assign _0703_ = _0658_ & \mchip.addr_cache [7];
	assign _0704_ = _0702_ & ~_0703_;
	assign _0705_ = \mchip.addr_cache [15] & ~_0655_;
	assign _0706_ = _0704_ & ~_0705_;
	assign io_out[7] = _0660_ & ~_0706_;
	assign _0707_ = ~(\mchip.bf.ucode [12] | \mchip.bf.ucode [11]);
	assign _0708_ = _0707_ & ~\mchip.bf.ucode [13];
	assign _0709_ = ~(_0708_ | _0086_);
	assign _0710_ = _0709_ | ~_0655_;
	assign _0711_ = _0086_ & ~_0660_;
	assign \mchip.next_state [0] = _0710_ & ~_0711_;
	assign \mchip.next_state [1] = _0656_ & ~_0711_;
	assign _0712_ = _0184_ & ~io_in[8];
	assign _0713_ = _0712_ | _0658_;
	assign \mchip.next_state [2] = _0713_ & ~_0711_;
	assign _0714_ = ~\mchip.bf.pc [1];
	assign _0715_ = ~(_0179_ | _0176_);
	assign _0716_ = _0715_ ^ _0714_;
	assign \mchip.bf.next_pc [1] = _0716_ ^ \mchip.bf.next_pc [0];
	assign _0717_ = _0715_ & ~_0714_;
	assign _0718_ = \mchip.bf.pc [0] & ~_0716_;
	assign _0719_ = _0718_ | _0717_;
	assign _0720_ = ~\mchip.bf.pc [2];
	assign _0721_ = _0715_ ^ _0720_;
	assign \mchip.bf.next_pc [2] = ~(_0721_ ^ _0719_);
	assign _0722_ = _0715_ & ~_0720_;
	assign _0723_ = _0719_ & ~_0721_;
	assign _0724_ = ~(_0723_ | _0722_);
	assign _0725_ = ~\mchip.bf.pc [3];
	assign _0726_ = _0715_ ^ _0725_;
	assign \mchip.bf.next_pc [3] = _0726_ ^ _0724_;
	assign _0727_ = _0726_ | _0721_;
	assign _0728_ = _0719_ & ~_0727_;
	assign _0729_ = _0715_ & ~_0725_;
	assign _0730_ = _0722_ & ~_0726_;
	assign _0731_ = _0730_ | _0729_;
	assign _0732_ = _0731_ | _0728_;
	assign _0733_ = ~\mchip.bf.pc [4];
	assign _0734_ = _0715_ ^ _0733_;
	assign \mchip.bf.next_pc [4] = ~(_0734_ ^ _0732_);
	assign _0735_ = _0715_ & ~_0733_;
	assign _0736_ = _0732_ & ~_0734_;
	assign _0737_ = ~(_0736_ | _0735_);
	assign _0738_ = ~\mchip.bf.pc [5];
	assign _0739_ = _0715_ ^ _0738_;
	assign \mchip.bf.next_pc [5] = _0739_ ^ _0737_;
	assign _0740_ = _0739_ | _0734_;
	assign _0741_ = _0732_ & ~_0740_;
	assign _0742_ = _0715_ & ~_0738_;
	assign _0743_ = _0735_ & ~_0739_;
	assign _0744_ = _0743_ | _0742_;
	assign _0745_ = _0744_ | _0741_;
	assign _0746_ = ~\mchip.bf.pc [6];
	assign _0747_ = _0715_ ^ _0746_;
	assign \mchip.bf.next_pc [6] = ~(_0747_ ^ _0745_);
	assign _0748_ = _0715_ & ~_0746_;
	assign _0749_ = _0745_ & ~_0747_;
	assign _0750_ = ~(_0749_ | _0748_);
	assign _0751_ = ~\mchip.bf.pc [7];
	assign _0752_ = _0715_ ^ _0751_;
	assign \mchip.bf.next_pc [7] = _0752_ ^ _0750_;
	assign _0753_ = _0752_ | _0747_;
	assign _0754_ = _0753_ | _0740_;
	assign _0755_ = _0732_ & ~_0754_;
	assign _0756_ = _0744_ & ~_0753_;
	assign _0757_ = _0715_ & ~_0751_;
	assign _0758_ = _0748_ & ~_0752_;
	assign _0759_ = _0758_ | _0757_;
	assign _0760_ = _0759_ | _0756_;
	assign _0761_ = _0760_ | _0755_;
	assign _0762_ = ~\mchip.bf.pc [8];
	assign _0763_ = _0715_ ^ _0762_;
	assign \mchip.bf.next_pc [8] = ~(_0763_ ^ _0761_);
	assign _0764_ = _0715_ & ~_0762_;
	assign _0765_ = _0761_ & ~_0763_;
	assign _0766_ = ~(_0765_ | _0764_);
	assign _0767_ = ~\mchip.bf.pc [9];
	assign _0768_ = _0715_ ^ _0767_;
	assign \mchip.bf.next_pc [9] = _0768_ ^ _0766_;
	assign _0769_ = _0768_ | _0763_;
	assign _0770_ = _0761_ & ~_0769_;
	assign _0771_ = _0715_ & ~_0767_;
	assign _0772_ = _0764_ & ~_0768_;
	assign _0773_ = _0772_ | _0771_;
	assign _0774_ = _0773_ | _0770_;
	assign _0775_ = ~\mchip.bf.pc [10];
	assign _0776_ = _0715_ ^ _0775_;
	assign \mchip.bf.next_pc [10] = ~(_0776_ ^ _0774_);
	assign _0777_ = _0715_ & ~_0775_;
	assign _0778_ = _0774_ & ~_0776_;
	assign _0779_ = ~(_0778_ | _0777_);
	assign _0780_ = ~\mchip.bf.pc [11];
	assign _0781_ = _0715_ ^ _0780_;
	assign \mchip.bf.next_pc [11] = _0781_ ^ _0779_;
	assign _0782_ = _0715_ & ~_0780_;
	assign _0783_ = _0777_ & ~_0781_;
	assign _0784_ = _0783_ | _0782_;
	assign _0785_ = _0781_ | _0776_;
	assign _0786_ = _0773_ & ~_0785_;
	assign _0787_ = _0786_ | _0784_;
	assign _0788_ = _0785_ | _0769_;
	assign _0789_ = _0761_ & ~_0788_;
	assign _0790_ = _0789_ | _0787_;
	assign _0791_ = _0715_ ^ \mchip.bf.pc [12];
	assign \mchip.bf.next_pc [12] = _0791_ ^ _0790_;
	assign _0792_ = _0715_ & \mchip.bf.pc [12];
	assign _0793_ = _0791_ & _0790_;
	assign _0794_ = _0793_ | _0792_;
	assign _0795_ = _0715_ ^ \mchip.bf.pc [13];
	assign \mchip.bf.next_pc [13] = _0795_ ^ _0794_;
	assign _0796_ = ~(_0715_ & \mchip.bf.pc [13]);
	assign _0797_ = ~(_0795_ & _0792_);
	assign _0798_ = ~(_0797_ & _0796_);
	assign _0799_ = ~(_0795_ & _0791_);
	assign _0800_ = _0790_ & ~_0799_;
	assign _0801_ = _0800_ | _0798_;
	assign _0802_ = _0715_ ^ \mchip.bf.pc [14];
	assign \mchip.bf.next_pc [14] = _0802_ ^ _0801_;
	assign _0803_ = ~(_0715_ & \mchip.bf.pc [14]);
	assign _0804_ = ~(_0802_ & _0801_);
	assign _0805_ = ~(_0804_ & _0803_);
	assign _0806_ = _0715_ ^ \mchip.bf.pc [15];
	assign \mchip.bf.next_pc [15] = _0806_ ^ _0805_;
	assign _0807_ = ~(_0182_ | _0181_);
	assign _0808_ = _0807_ ^ _0593_;
	assign \mchip.bf.next_cursor [1] = _0808_ ^ \mchip.bf.next_cursor [0];
	assign _0005_ = _0807_ & ~_0593_;
	assign _0006_ = \mchip.bf.cursor [0] & ~_0808_;
	assign _0007_ = _0006_ | _0005_;
	assign _0008_ = _0807_ ^ _0597_;
	assign \mchip.bf.next_cursor [2] = ~(_0008_ ^ _0007_);
	assign _0009_ = _0807_ & ~_0597_;
	assign _0010_ = _0007_ & ~_0008_;
	assign _0011_ = ~(_0010_ | _0009_);
	assign _0012_ = _0807_ ^ _0601_;
	assign \mchip.bf.next_cursor [3] = _0012_ ^ _0011_;
	assign _0013_ = _0012_ | _0008_;
	assign _0014_ = _0007_ & ~_0013_;
	assign _0015_ = _0807_ & ~_0601_;
	assign _0016_ = _0009_ & ~_0012_;
	assign _0017_ = _0016_ | _0015_;
	assign _0018_ = _0017_ | _0014_;
	assign _0019_ = _0807_ ^ _0605_;
	assign \mchip.bf.next_cursor [4] = ~(_0019_ ^ _0018_);
	assign _0020_ = _0807_ & ~_0605_;
	assign _0021_ = _0018_ & ~_0019_;
	assign _0022_ = ~(_0021_ | _0020_);
	assign _0023_ = _0807_ ^ _0609_;
	assign \mchip.bf.next_cursor [5] = _0023_ ^ _0022_;
	assign _0024_ = _0023_ | _0019_;
	assign _0025_ = _0018_ & ~_0024_;
	assign _0026_ = _0807_ & ~_0609_;
	assign _0027_ = _0020_ & ~_0023_;
	assign _0028_ = _0027_ | _0026_;
	assign _0029_ = _0028_ | _0025_;
	assign _0030_ = _0807_ ^ _0613_;
	assign \mchip.bf.next_cursor [6] = ~(_0030_ ^ _0029_);
	assign _0031_ = _0807_ & ~_0613_;
	assign _0032_ = _0029_ & ~_0030_;
	assign _0033_ = ~(_0032_ | _0031_);
	assign _0034_ = _0807_ ^ _0617_;
	assign \mchip.bf.next_cursor [7] = _0034_ ^ _0033_;
	assign _0035_ = _0034_ | _0030_;
	assign _0036_ = _0035_ | _0024_;
	assign _0037_ = _0018_ & ~_0036_;
	assign _0038_ = _0028_ & ~_0035_;
	assign _0039_ = _0807_ & ~_0617_;
	assign _0040_ = _0031_ & ~_0034_;
	assign _0041_ = _0040_ | _0039_;
	assign _0042_ = _0041_ | _0038_;
	assign _0043_ = _0042_ | _0037_;
	assign _0044_ = _0807_ ^ _0621_;
	assign \mchip.bf.next_cursor [8] = ~(_0044_ ^ _0043_);
	assign _0045_ = _0807_ & ~_0621_;
	assign _0046_ = _0043_ & ~_0044_;
	assign _0047_ = ~(_0046_ | _0045_);
	assign _0048_ = _0807_ ^ _0625_;
	assign \mchip.bf.next_cursor [9] = _0048_ ^ _0047_;
	assign _0049_ = _0048_ | _0044_;
	assign _0050_ = _0043_ & ~_0049_;
	assign _0051_ = _0807_ & ~_0625_;
	assign _0052_ = _0045_ & ~_0048_;
	assign _0053_ = _0052_ | _0051_;
	assign _0054_ = _0053_ | _0050_;
	assign _0055_ = _0807_ ^ _0629_;
	assign \mchip.bf.next_cursor [10] = ~(_0055_ ^ _0054_);
	assign _0056_ = _0807_ & ~_0629_;
	assign _0057_ = _0054_ & ~_0055_;
	assign _0058_ = ~(_0057_ | _0056_);
	assign _0059_ = _0807_ ^ _0633_;
	assign \mchip.bf.next_cursor [11] = _0059_ ^ _0058_;
	assign _0060_ = _0807_ & ~_0633_;
	assign _0061_ = _0056_ & ~_0059_;
	assign _0062_ = _0061_ | _0060_;
	assign _0063_ = _0059_ | _0055_;
	assign _0064_ = _0053_ & ~_0063_;
	assign _0065_ = _0064_ | _0062_;
	assign _0066_ = _0063_ | _0049_;
	assign _0067_ = _0043_ & ~_0066_;
	assign _0068_ = _0067_ | _0065_;
	assign _0069_ = _0807_ ^ \mchip.bf.cursor [12];
	assign \mchip.bf.next_cursor [12] = _0069_ ^ _0068_;
	assign _0070_ = _0807_ & ~_0637_;
	assign _0071_ = _0069_ & _0068_;
	assign _0072_ = _0071_ | _0070_;
	assign _0073_ = _0807_ ^ \mchip.bf.cursor [13];
	assign \mchip.bf.next_cursor [13] = _0073_ ^ _0072_;
	assign _0074_ = _0807_ & ~_0641_;
	assign _0075_ = _0073_ & _0070_;
	assign _0076_ = _0075_ | _0074_;
	assign _0077_ = ~(_0073_ & _0069_);
	assign _0078_ = _0068_ & ~_0077_;
	assign _0079_ = _0078_ | _0076_;
	assign _0080_ = _0807_ ^ \mchip.bf.cursor [14];
	assign \mchip.bf.next_cursor [14] = _0080_ ^ _0079_;
	assign _0081_ = _0807_ & ~_0645_;
	assign _0082_ = _0080_ & _0079_;
	assign _0083_ = _0082_ | _0081_;
	assign _0084_ = _0807_ ^ \mchip.bf.cursor [15];
	assign \mchip.bf.next_cursor [15] = _0084_ ^ _0083_;
	always @(posedge io_in[12]) \mchip.bf.state [0] <= _0809_[0];
	always @(posedge io_in[12]) \mchip.bf.state [1] <= _0809_[1];
	always @(posedge io_in[12]) \mchip.bf.state [2] <= _0809_[2];
	always @(posedge io_in[12]) \mchip.bf.state [3] <= _0809_[3];
	always @(posedge io_in[12]) \mchip.bf.state [4] <= _0809_[4];
	always @(posedge io_in[12]) \mchip.bf.state [5] <= _0809_[5];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.bf.cursor [0] <= 1'h0;
		else if (_0003_)
			\mchip.bf.cursor [0] <= \mchip.bf.next_cursor [0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.bf.cursor [1] <= 1'h0;
		else if (_0003_)
			\mchip.bf.cursor [1] <= \mchip.bf.next_cursor [1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.bf.cursor [2] <= 1'h0;
		else if (_0003_)
			\mchip.bf.cursor [2] <= \mchip.bf.next_cursor [2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.bf.cursor [3] <= 1'h0;
		else if (_0003_)
			\mchip.bf.cursor [3] <= \mchip.bf.next_cursor [3];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.bf.cursor [4] <= 1'h0;
		else if (_0003_)
			\mchip.bf.cursor [4] <= \mchip.bf.next_cursor [4];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.bf.cursor [5] <= 1'h0;
		else if (_0003_)
			\mchip.bf.cursor [5] <= \mchip.bf.next_cursor [5];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.bf.cursor [6] <= 1'h0;
		else if (_0003_)
			\mchip.bf.cursor [6] <= \mchip.bf.next_cursor [6];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.bf.cursor [7] <= 1'h0;
		else if (_0003_)
			\mchip.bf.cursor [7] <= \mchip.bf.next_cursor [7];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.bf.cursor [8] <= 1'h0;
		else if (_0003_)
			\mchip.bf.cursor [8] <= \mchip.bf.next_cursor [8];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.bf.cursor [9] <= 1'h0;
		else if (_0003_)
			\mchip.bf.cursor [9] <= \mchip.bf.next_cursor [9];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.bf.cursor [10] <= 1'h0;
		else if (_0003_)
			\mchip.bf.cursor [10] <= \mchip.bf.next_cursor [10];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.bf.cursor [11] <= 1'h0;
		else if (_0003_)
			\mchip.bf.cursor [11] <= \mchip.bf.next_cursor [11];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.bf.cursor [12] <= 1'h0;
		else if (_0003_)
			\mchip.bf.cursor [12] <= \mchip.bf.next_cursor [12];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.bf.cursor [13] <= 1'h0;
		else if (_0003_)
			\mchip.bf.cursor [13] <= \mchip.bf.next_cursor [13];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.bf.cursor [14] <= 1'h0;
		else if (_0003_)
			\mchip.bf.cursor [14] <= \mchip.bf.next_cursor [14];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.bf.cursor [15] <= 1'h0;
		else if (_0003_)
			\mchip.bf.cursor [15] <= \mchip.bf.next_cursor [15];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.bf.pc [0] <= 1'h0;
		else if (_0002_)
			\mchip.bf.pc [0] <= \mchip.bf.next_pc [0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.bf.pc [1] <= 1'h0;
		else if (_0002_)
			\mchip.bf.pc [1] <= \mchip.bf.next_pc [1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.bf.pc [2] <= 1'h0;
		else if (_0002_)
			\mchip.bf.pc [2] <= \mchip.bf.next_pc [2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.bf.pc [3] <= 1'h0;
		else if (_0002_)
			\mchip.bf.pc [3] <= \mchip.bf.next_pc [3];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.bf.pc [4] <= 1'h0;
		else if (_0002_)
			\mchip.bf.pc [4] <= \mchip.bf.next_pc [4];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.bf.pc [5] <= 1'h0;
		else if (_0002_)
			\mchip.bf.pc [5] <= \mchip.bf.next_pc [5];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.bf.pc [6] <= 1'h0;
		else if (_0002_)
			\mchip.bf.pc [6] <= \mchip.bf.next_pc [6];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.bf.pc [7] <= 1'h0;
		else if (_0002_)
			\mchip.bf.pc [7] <= \mchip.bf.next_pc [7];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.bf.pc [8] <= 1'h0;
		else if (_0002_)
			\mchip.bf.pc [8] <= \mchip.bf.next_pc [8];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.bf.pc [9] <= 1'h0;
		else if (_0002_)
			\mchip.bf.pc [9] <= \mchip.bf.next_pc [9];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.bf.pc [10] <= 1'h0;
		else if (_0002_)
			\mchip.bf.pc [10] <= \mchip.bf.next_pc [10];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.bf.pc [11] <= 1'h0;
		else if (_0002_)
			\mchip.bf.pc [11] <= \mchip.bf.next_pc [11];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.bf.pc [12] <= 1'h0;
		else if (_0002_)
			\mchip.bf.pc [12] <= \mchip.bf.next_pc [12];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.bf.pc [13] <= 1'h0;
		else if (_0002_)
			\mchip.bf.pc [13] <= \mchip.bf.next_pc [13];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.bf.pc [14] <= 1'h0;
		else if (_0002_)
			\mchip.bf.pc [14] <= \mchip.bf.next_pc [14];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.bf.pc [15] <= 1'h0;
		else if (_0002_)
			\mchip.bf.pc [15] <= \mchip.bf.next_pc [15];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.bf.acc [0] <= 1'h0;
		else if (_0001_)
			\mchip.bf.acc [0] <= \mchip.val_in [0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.bf.acc [1] <= 1'h0;
		else if (_0001_)
			\mchip.bf.acc [1] <= \mchip.val_in [1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.bf.acc [2] <= 1'h0;
		else if (_0001_)
			\mchip.bf.acc [2] <= \mchip.val_in [2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.bf.acc [3] <= 1'h0;
		else if (_0001_)
			\mchip.bf.acc [3] <= \mchip.val_in [3];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.bf.acc [4] <= 1'h0;
		else if (_0001_)
			\mchip.bf.acc [4] <= \mchip.val_in [4];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.bf.acc [5] <= 1'h0;
		else if (_0001_)
			\mchip.bf.acc [5] <= \mchip.val_in [5];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.bf.acc [6] <= 1'h0;
		else if (_0001_)
			\mchip.bf.acc [6] <= \mchip.val_in [6];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.bf.acc [7] <= 1'h0;
		else if (_0001_)
			\mchip.bf.acc [7] <= \mchip.val_in [7];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.bf.depth [0] <= 1'h0;
		else if (_0000_)
			\mchip.bf.depth [0] <= \mchip.bf.next_depth [0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.bf.depth [1] <= 1'h0;
		else if (_0000_)
			\mchip.bf.depth [1] <= \mchip.bf.next_depth [1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.bf.depth [2] <= 1'h0;
		else if (_0000_)
			\mchip.bf.depth [2] <= \mchip.bf.next_depth [2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.bf.depth [3] <= 1'h0;
		else if (_0000_)
			\mchip.bf.depth [3] <= \mchip.bf.next_depth [3];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.bf.depth [4] <= 1'h0;
		else if (_0000_)
			\mchip.bf.depth [4] <= \mchip.bf.next_depth [4];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.bf.depth [5] <= 1'h0;
		else if (_0000_)
			\mchip.bf.depth [5] <= \mchip.bf.next_depth [5];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.bf.depth [6] <= 1'h0;
		else if (_0000_)
			\mchip.bf.depth [6] <= \mchip.bf.next_depth [6];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.bf.depth [7] <= 1'h0;
		else if (_0000_)
			\mchip.bf.depth [7] <= \mchip.bf.next_depth [7];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.bf.depth [8] <= 1'h0;
		else if (_0000_)
			\mchip.bf.depth [8] <= \mchip.bf.next_depth [8];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.bf.depth [9] <= 1'h0;
		else if (_0000_)
			\mchip.bf.depth [9] <= \mchip.bf.next_depth [9];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.bf.depth [10] <= 1'h0;
		else if (_0000_)
			\mchip.bf.depth [10] <= \mchip.bf.next_depth [10];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.bf.depth [11] <= 1'h0;
		else if (_0000_)
			\mchip.bf.depth [11] <= \mchip.bf.next_depth [11];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.val_cache [0] <= 1'h0;
		else if (\mchip.bf.enable )
			\mchip.val_cache [0] <= \mchip.val_out [0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.val_cache [1] <= 1'h0;
		else if (\mchip.bf.enable )
			\mchip.val_cache [1] <= \mchip.val_out [1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.val_cache [2] <= 1'h0;
		else if (\mchip.bf.enable )
			\mchip.val_cache [2] <= \mchip.val_out [2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.val_cache [3] <= 1'h0;
		else if (\mchip.bf.enable )
			\mchip.val_cache [3] <= \mchip.val_out [3];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.val_cache [4] <= 1'h0;
		else if (\mchip.bf.enable )
			\mchip.val_cache [4] <= \mchip.val_out [4];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.val_cache [5] <= 1'h0;
		else if (\mchip.bf.enable )
			\mchip.val_cache [5] <= \mchip.val_out [5];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.val_cache [6] <= 1'h0;
		else if (\mchip.bf.enable )
			\mchip.val_cache [6] <= \mchip.val_out [6];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.val_cache [7] <= 1'h0;
		else if (\mchip.bf.enable )
			\mchip.val_cache [7] <= \mchip.val_out [7];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.addr_cache [0] <= 1'h0;
		else if (\mchip.bf.enable )
			\mchip.addr_cache [0] <= \mchip.addr [0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.addr_cache [1] <= 1'h0;
		else if (\mchip.bf.enable )
			\mchip.addr_cache [1] <= \mchip.addr [1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.addr_cache [2] <= 1'h0;
		else if (\mchip.bf.enable )
			\mchip.addr_cache [2] <= \mchip.addr [2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.addr_cache [3] <= 1'h0;
		else if (\mchip.bf.enable )
			\mchip.addr_cache [3] <= \mchip.addr [3];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.addr_cache [4] <= 1'h0;
		else if (\mchip.bf.enable )
			\mchip.addr_cache [4] <= \mchip.addr [4];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.addr_cache [5] <= 1'h0;
		else if (\mchip.bf.enable )
			\mchip.addr_cache [5] <= \mchip.addr [5];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.addr_cache [6] <= 1'h0;
		else if (\mchip.bf.enable )
			\mchip.addr_cache [6] <= \mchip.addr [6];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.addr_cache [7] <= 1'h0;
		else if (\mchip.bf.enable )
			\mchip.addr_cache [7] <= \mchip.addr [7];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.addr_cache [8] <= 1'h0;
		else if (\mchip.bf.enable )
			\mchip.addr_cache [8] <= \mchip.addr [8];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.addr_cache [9] <= 1'h0;
		else if (\mchip.bf.enable )
			\mchip.addr_cache [9] <= \mchip.addr [9];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.addr_cache [10] <= 1'h0;
		else if (\mchip.bf.enable )
			\mchip.addr_cache [10] <= \mchip.addr [10];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.addr_cache [11] <= 1'h0;
		else if (\mchip.bf.enable )
			\mchip.addr_cache [11] <= \mchip.addr [11];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.addr_cache [12] <= 1'h0;
		else if (\mchip.bf.enable )
			\mchip.addr_cache [12] <= \mchip.addr [12];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.addr_cache [13] <= 1'h0;
		else if (\mchip.bf.enable )
			\mchip.addr_cache [13] <= \mchip.addr [13];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.addr_cache [14] <= 1'h0;
		else if (\mchip.bf.enable )
			\mchip.addr_cache [14] <= \mchip.addr [14];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.addr_cache [15] <= 1'h0;
		else if (\mchip.bf.enable )
			\mchip.addr_cache [15] <= \mchip.addr [15];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.op_cache [0] <= 1'h0;
		else if (\mchip.bf.enable )
			\mchip.op_cache [0] <= \mchip.bf.ucode [11];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.op_cache [1] <= 1'h0;
		else if (\mchip.bf.enable )
			\mchip.op_cache [1] <= \mchip.bf.ucode [12];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.op_cache [2] <= 1'h0;
		else if (\mchip.bf.enable )
			\mchip.op_cache [2] <= \mchip.bf.ucode [13];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.state [0] <= 1'h0;
		else if (io_in[9])
			\mchip.state [0] <= \mchip.next_state [0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.state [1] <= 1'h0;
		else if (io_in[9])
			\mchip.state [1] <= \mchip.next_state [1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.state [2] <= 1'h0;
		else if (io_in[9])
			\mchip.state [2] <= \mchip.next_state [2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.val_in [0] <= 1'h0;
		else if (_0004_)
			\mchip.val_in [0] <= io_in[0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.val_in [1] <= 1'h0;
		else if (_0004_)
			\mchip.val_in [1] <= io_in[1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.val_in [2] <= 1'h0;
		else if (_0004_)
			\mchip.val_in [2] <= io_in[2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.val_in [3] <= 1'h0;
		else if (_0004_)
			\mchip.val_in [3] <= io_in[3];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.val_in [4] <= 1'h0;
		else if (_0004_)
			\mchip.val_in [4] <= io_in[4];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.val_in [5] <= 1'h0;
		else if (_0004_)
			\mchip.val_in [5] <= io_in[5];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.val_in [6] <= 1'h0;
		else if (_0004_)
			\mchip.val_in [6] <= io_in[6];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.val_in [7] <= 1'h0;
		else if (_0004_)
			\mchip.val_in [7] <= io_in[7];
	assign io_out[13:8] = {2'h0, \mchip.bf.halted , \mchip.state };
	assign \mchip.bf.addr  = \mchip.addr ;
	assign \mchip.bf.bus_op  = \mchip.bf.ucode [13:11];
	assign \mchip.bf.clock  = io_in[12];
	assign \mchip.bf.next_acc  = \mchip.val_in ;
	assign \mchip.bf.reset  = io_in[13];
	assign \mchip.bf.ucode [10:0] = 11'h000;
	assign \mchip.bf.val_in  = \mchip.val_in ;
	assign \mchip.bf.val_out  = \mchip.val_out ;
	assign \mchip.bus_in  = io_in[7:0];
	assign \mchip.bus_op  = \mchip.bf.ucode [13:11];
	assign \mchip.bus_out  = io_out[7:0];
	assign \mchip.clock  = io_in[12];
	assign \mchip.enable  = io_in[9];
	assign \mchip.halted  = \mchip.bf.halted ;
	assign \mchip.io_in  = io_in[11:0];
	assign \mchip.io_out  = {\mchip.bf.halted , \mchip.state , io_out[7:0]};
	assign \mchip.op_done  = io_in[8];
	assign \mchip.reset  = io_in[13];
endmodule
module d12_oball_i2c (
	io_in,
	io_out
);
	wire _0000_;
	wire _0001_;
	wire _0002_;
	wire _0003_;
	wire _0004_;
	wire _0005_;
	wire _0006_;
	wire _0007_;
	wire _0008_;
	wire _0009_;
	wire _0010_;
	wire _0011_;
	wire _0012_;
	wire _0013_;
	wire _0014_;
	wire _0015_;
	wire _0016_;
	wire _0017_;
	wire _0018_;
	wire _0019_;
	wire _0020_;
	wire _0021_;
	wire _0022_;
	wire _0023_;
	wire _0024_;
	wire _0025_;
	wire _0026_;
	wire _0027_;
	wire _0028_;
	wire _0029_;
	wire _0030_;
	wire _0031_;
	wire _0032_;
	wire _0033_;
	wire _0034_;
	wire _0035_;
	wire _0036_;
	wire _0037_;
	wire _0038_;
	wire _0039_;
	wire _0040_;
	wire _0041_;
	wire _0042_;
	wire _0043_;
	wire _0044_;
	wire _0045_;
	wire _0046_;
	wire _0047_;
	wire _0048_;
	wire _0049_;
	wire _0050_;
	wire _0051_;
	wire _0052_;
	wire _0053_;
	wire _0054_;
	wire _0055_;
	wire _0056_;
	wire _0057_;
	wire _0058_;
	wire _0059_;
	wire _0060_;
	wire _0061_;
	wire _0062_;
	wire _0063_;
	wire _0064_;
	wire _0065_;
	wire _0066_;
	wire _0067_;
	wire _0068_;
	wire _0069_;
	wire _0070_;
	wire _0071_;
	wire _0072_;
	wire _0073_;
	wire _0074_;
	wire _0075_;
	wire _0076_;
	wire _0077_;
	wire _0078_;
	wire _0079_;
	wire _0080_;
	wire _0081_;
	wire _0082_;
	wire _0083_;
	wire _0084_;
	wire _0085_;
	wire _0086_;
	wire _0087_;
	wire _0088_;
	wire _0089_;
	wire _0090_;
	wire _0091_;
	wire _0092_;
	wire _0093_;
	wire _0094_;
	wire _0095_;
	wire _0096_;
	wire _0097_;
	wire _0098_;
	wire _0099_;
	wire _0100_;
	wire _0101_;
	wire _0102_;
	wire _0103_;
	wire _0104_;
	wire _0105_;
	wire _0106_;
	wire _0107_;
	wire _0108_;
	wire _0109_;
	wire _0110_;
	wire _0111_;
	wire _0112_;
	wire _0113_;
	wire _0114_;
	wire _0115_;
	wire _0116_;
	wire _0117_;
	wire _0118_;
	wire _0119_;
	wire _0120_;
	reg _0121_;
	reg _0122_;
	reg _0123_;
	reg _0124_;
	reg _0125_;
	reg _0126_;
	reg _0127_;
	reg _0128_;
	reg _0129_;
	reg _0130_;
	reg _0131_;
	reg _0132_;
	reg _0133_;
	reg _0134_;
	reg _0135_;
	reg _0136_;
	reg _0137_;
	reg _0138_;
	reg _0139_;
	reg _0140_;
	reg _0141_;
	reg _0142_;
	reg _0143_;
	reg _0144_;
	reg _0145_;
	reg _0146_;
	reg _0147_;
	reg _0148_;
	reg _0149_;
	reg _0150_;
	reg _0151_;
	reg _0152_;
	reg _0153_;
	reg _0154_;
	reg _0155_;
	reg _0156_;
	reg _0157_;
	reg _0158_;
	reg _0159_;
	reg _0160_;
	reg _0161_;
	reg _0162_;
	reg _0163_;
	reg _0164_;
	reg _0165_;
	reg _0166_;
	reg _0167_;
	reg _0168_;
	reg _0169_;
	reg _0170_;
	reg _0171_;
	reg _0172_;
	reg _0173_;
	reg _0174_;
	reg _0175_;
	reg _0176_;
	reg _0177_;
	reg _0178_;
	reg _0179_;
	reg _0180_;
	reg _0181_;
	reg _0182_;
	reg _0183_;
	reg _0184_;
	reg _0185_;
	reg _0186_;
	reg _0187_;
	reg _0188_;
	reg _0189_;
	reg _0190_;
	reg _0191_;
	reg _0192_;
	reg _0193_;
	reg _0194_;
	reg _0195_;
	reg _0196_;
	reg _0197_;
	reg _0198_;
	reg _0199_;
	reg _0200_;
	reg _0201_;
	reg _0202_;
	reg _0203_;
	reg _0204_;
	reg _0205_;
	reg _0206_;
	reg _0207_;
	reg _0208_;
	reg _0209_;
	reg _0210_;
	reg _0211_;
	reg _0212_;
	reg _0213_;
	reg _0214_;
	reg _0215_;
	reg _0216_;
	reg _0217_;
	reg _0218_;
	reg _0219_;
	reg _0220_;
	reg _0221_;
	reg _0222_;
	reg _0223_;
	reg _0224_;
	reg _0225_;
	reg _0226_;
	reg _0227_;
	reg _0228_;
	reg _0229_;
	reg _0230_;
	reg _0231_;
	reg _0232_;
	reg _0233_;
	reg _0234_;
	reg _0235_;
	reg _0236_;
	reg _0237_;
	reg _0238_;
	reg _0239_;
	reg _0240_;
	reg _0241_;
	reg _0242_;
	reg _0243_;
	reg _0244_;
	reg _0245_;
	reg _0246_;
	reg _0247_;
	reg _0248_;
	reg _0249_;
	reg _0250_;
	reg _0251_;
	reg _0252_;
	reg _0253_;
	reg _0254_;
	reg _0255_;
	reg _0256_;
	reg _0257_;
	reg _0258_;
	reg _0259_;
	reg _0260_;
	reg _0261_;
	reg _0262_;
	reg _0263_;
	reg _0264_;
	reg _0265_;
	reg _0266_;
	reg _0267_;
	reg _0268_;
	reg _0269_;
	reg _0270_;
	reg _0271_;
	reg _0272_;
	reg _0273_;
	reg _0274_;
	reg _0275_;
	reg _0276_;
	reg _0277_;
	reg _0278_;
	reg _0279_;
	reg _0280_;
	reg _0281_;
	reg _0282_;
	reg _0283_;
	reg _0284_;
	reg _0285_;
	reg _0286_;
	reg _0287_;
	reg _0288_;
	reg _0289_;
	reg _0290_;
	reg _0291_;
	reg _0292_;
	reg _0293_;
	reg _0294_;
	reg _0295_;
	reg _0296_;
	reg _0297_;
	reg _0298_;
	reg _0299_;
	reg _0300_;
	reg _0301_;
	reg _0302_;
	reg _0303_;
	reg _0304_;
	reg _0305_;
	reg _0306_;
	reg _0307_;
	reg _0308_;
	reg _0309_;
	reg _0310_;
	reg _0311_;
	reg _0312_;
	reg _0313_;
	reg _0314_;
	reg _0315_;
	reg _0316_;
	reg _0317_;
	reg _0318_;
	reg _0319_;
	reg _0320_;
	reg _0321_;
	reg _0322_;
	reg _0323_;
	reg _0324_;
	reg _0325_;
	reg _0326_;
	reg _0327_;
	reg _0328_;
	reg _0329_;
	reg _0330_;
	reg _0331_;
	reg _0332_;
	reg _0333_;
	reg _0334_;
	reg _0335_;
	reg _0336_;
	reg _0337_;
	reg _0338_;
	reg _0339_;
	reg _0340_;
	reg _0341_;
	reg _0342_;
	reg _0343_;
	reg _0344_;
	reg _0345_;
	reg _0346_;
	reg _0347_;
	reg _0348_;
	reg _0349_;
	reg _0350_;
	reg _0351_;
	reg _0352_;
	reg _0353_;
	reg _0354_;
	reg _0355_;
	reg _0356_;
	reg _0357_;
	reg _0358_;
	reg _0359_;
	reg _0360_;
	reg _0361_;
	reg _0362_;
	reg _0363_;
	reg _0364_;
	reg _0365_;
	reg _0366_;
	reg _0367_;
	reg _0368_;
	reg _0369_;
	reg _0370_;
	reg _0371_;
	reg _0372_;
	reg _0373_;
	reg _0374_;
	reg _0375_;
	reg _0376_;
	reg _0377_;
	reg _0378_;
	reg _0379_;
	reg _0380_;
	reg _0381_;
	reg _0382_;
	reg _0383_;
	reg _0384_;
	reg _0385_;
	reg _0386_;
	reg _0387_;
	reg _0388_;
	reg _0389_;
	reg _0390_;
	reg _0391_;
	reg _0392_;
	reg _0393_;
	reg _0394_;
	reg _0395_;
	reg _0396_;
	reg _0397_;
	reg _0398_;
	reg _0399_;
	reg _0400_;
	reg _0401_;
	reg _0402_;
	reg _0403_;
	reg _0404_;
	wire _0405_;
	wire _0406_;
	wire _0407_;
	wire _0408_;
	wire _0409_;
	wire _0410_;
	wire _0411_;
	wire _0412_;
	wire _0413_;
	wire _0414_;
	wire _0415_;
	wire _0416_;
	wire _0417_;
	wire _0418_;
	wire _0419_;
	wire _0420_;
	wire _0421_;
	wire _0422_;
	wire _0423_;
	wire _0424_;
	wire _0425_;
	wire _0426_;
	wire _0427_;
	wire _0428_;
	wire _0429_;
	wire _0430_;
	wire _0431_;
	wire _0432_;
	wire _0433_;
	wire _0434_;
	wire _0435_;
	wire _0436_;
	wire _0437_;
	wire _0438_;
	wire _0439_;
	wire _0440_;
	wire _0441_;
	wire _0442_;
	wire _0443_;
	wire _0444_;
	wire _0445_;
	wire _0446_;
	wire _0447_;
	wire _0448_;
	wire _0449_;
	wire _0450_;
	wire _0451_;
	wire _0452_;
	wire _0453_;
	wire _0454_;
	wire _0455_;
	wire _0456_;
	wire _0457_;
	wire _0458_;
	wire _0459_;
	wire _0460_;
	wire _0461_;
	wire _0462_;
	wire _0463_;
	wire _0464_;
	wire _0465_;
	wire _0466_;
	wire _0467_;
	wire _0468_;
	wire _0469_;
	wire _0470_;
	wire _0471_;
	wire _0472_;
	wire _0473_;
	wire _0474_;
	wire _0475_;
	wire _0476_;
	wire _0477_;
	wire _0478_;
	wire _0479_;
	wire _0480_;
	wire _0481_;
	wire _0482_;
	wire _0483_;
	wire _0484_;
	wire _0485_;
	wire _0486_;
	wire _0487_;
	wire _0488_;
	wire _0489_;
	wire _0490_;
	wire _0491_;
	wire _0492_;
	wire _0493_;
	wire _0494_;
	wire _0495_;
	wire _0496_;
	wire _0497_;
	wire _0498_;
	wire _0499_;
	wire _0500_;
	wire _0501_;
	wire _0502_;
	wire _0503_;
	wire _0504_;
	wire _0505_;
	wire _0506_;
	wire _0507_;
	wire _0508_;
	wire _0509_;
	wire _0510_;
	wire _0511_;
	wire _0512_;
	wire _0513_;
	wire _0514_;
	wire _0515_;
	wire _0516_;
	wire _0517_;
	wire _0518_;
	wire _0519_;
	wire _0520_;
	wire _0521_;
	wire _0522_;
	wire _0523_;
	wire _0524_;
	wire _0525_;
	wire _0526_;
	wire _0527_;
	wire _0528_;
	wire _0529_;
	wire _0530_;
	wire _0531_;
	wire _0532_;
	wire _0533_;
	wire _0534_;
	wire _0535_;
	wire _0536_;
	wire _0537_;
	wire _0538_;
	wire _0539_;
	wire _0540_;
	wire _0541_;
	wire _0542_;
	wire _0543_;
	wire _0544_;
	wire _0545_;
	wire _0546_;
	wire _0547_;
	wire _0548_;
	wire _0549_;
	wire _0550_;
	wire _0551_;
	wire _0552_;
	wire _0553_;
	wire _0554_;
	wire _0555_;
	wire _0556_;
	wire _0557_;
	wire _0558_;
	wire _0559_;
	wire _0560_;
	wire _0561_;
	wire _0562_;
	wire _0563_;
	wire _0564_;
	wire _0565_;
	wire _0566_;
	wire _0567_;
	wire _0568_;
	wire _0569_;
	wire _0570_;
	wire _0571_;
	wire _0572_;
	wire _0573_;
	wire _0574_;
	wire _0575_;
	wire _0576_;
	wire _0577_;
	wire _0578_;
	wire _0579_;
	wire _0580_;
	wire _0581_;
	wire _0582_;
	wire _0583_;
	wire _0584_;
	wire _0585_;
	wire _0586_;
	wire _0587_;
	wire _0588_;
	wire _0589_;
	wire _0590_;
	wire _0591_;
	wire _0592_;
	wire _0593_;
	wire _0594_;
	wire _0595_;
	wire _0596_;
	wire _0597_;
	wire _0598_;
	wire _0599_;
	wire _0600_;
	wire _0601_;
	wire _0602_;
	wire _0603_;
	wire _0604_;
	wire _0605_;
	wire _0606_;
	wire _0607_;
	wire _0608_;
	wire _0609_;
	wire _0610_;
	wire _0611_;
	wire _0612_;
	wire _0613_;
	wire _0614_;
	wire _0615_;
	wire _0616_;
	wire _0617_;
	wire _0618_;
	wire _0619_;
	wire _0620_;
	wire _0621_;
	wire _0622_;
	wire _0623_;
	wire _0624_;
	wire _0625_;
	wire _0626_;
	wire _0627_;
	wire _0628_;
	wire _0629_;
	wire _0630_;
	wire _0631_;
	wire _0632_;
	wire _0633_;
	wire _0634_;
	wire _0635_;
	wire _0636_;
	wire _0637_;
	wire _0638_;
	wire _0639_;
	wire _0640_;
	wire _0641_;
	wire _0642_;
	wire _0643_;
	wire _0644_;
	wire _0645_;
	wire _0646_;
	wire _0647_;
	wire _0648_;
	wire _0649_;
	wire _0650_;
	wire _0651_;
	wire _0652_;
	wire _0653_;
	wire _0654_;
	wire _0655_;
	wire _0656_;
	wire _0657_;
	wire _0658_;
	wire _0659_;
	wire _0660_;
	wire _0661_;
	wire _0662_;
	wire _0663_;
	wire _0664_;
	wire _0665_;
	wire _0666_;
	wire _0667_;
	wire _0668_;
	wire _0669_;
	wire _0670_;
	wire _0671_;
	wire _0672_;
	wire _0673_;
	wire _0674_;
	wire _0675_;
	wire _0676_;
	wire _0677_;
	wire _0678_;
	wire _0679_;
	wire _0680_;
	wire _0681_;
	wire _0682_;
	wire _0683_;
	wire _0684_;
	wire _0685_;
	wire _0686_;
	wire _0687_;
	wire _0688_;
	wire _0689_;
	wire _0690_;
	wire _0691_;
	wire _0692_;
	wire _0693_;
	wire _0694_;
	wire _0695_;
	wire _0696_;
	wire _0697_;
	wire _0698_;
	wire _0699_;
	wire _0700_;
	wire _0701_;
	wire _0702_;
	wire _0703_;
	wire _0704_;
	wire _0705_;
	wire _0706_;
	wire _0707_;
	wire _0708_;
	wire _0709_;
	wire _0710_;
	wire _0711_;
	wire _0712_;
	wire _0713_;
	wire _0714_;
	wire _0715_;
	wire _0716_;
	wire _0717_;
	wire _0718_;
	wire _0719_;
	wire _0720_;
	wire _0721_;
	wire _0722_;
	wire _0723_;
	wire _0724_;
	wire _0725_;
	wire _0726_;
	wire _0727_;
	wire _0728_;
	wire _0729_;
	wire _0730_;
	wire _0731_;
	wire _0732_;
	wire _0733_;
	wire _0734_;
	wire _0735_;
	wire _0736_;
	wire _0737_;
	wire _0738_;
	wire _0739_;
	wire _0740_;
	wire _0741_;
	wire _0742_;
	wire _0743_;
	wire _0744_;
	wire _0745_;
	wire _0746_;
	wire _0747_;
	wire _0748_;
	wire _0749_;
	wire _0750_;
	wire _0751_;
	wire _0752_;
	wire _0753_;
	wire _0754_;
	wire _0755_;
	wire _0756_;
	wire _0757_;
	wire _0758_;
	wire _0759_;
	wire _0760_;
	wire _0761_;
	wire _0762_;
	wire _0763_;
	wire _0764_;
	wire _0765_;
	wire _0766_;
	wire _0767_;
	wire _0768_;
	wire _0769_;
	wire _0770_;
	wire _0771_;
	wire _0772_;
	wire _0773_;
	wire _0774_;
	wire _0775_;
	wire _0776_;
	wire _0777_;
	wire _0778_;
	wire _0779_;
	wire _0780_;
	wire _0781_;
	wire _0782_;
	wire _0783_;
	wire _0784_;
	wire _0785_;
	wire _0786_;
	wire _0787_;
	wire _0788_;
	wire _0789_;
	wire _0790_;
	wire _0791_;
	wire _0792_;
	wire _0793_;
	wire _0794_;
	wire _0795_;
	wire _0796_;
	wire _0797_;
	wire _0798_;
	wire _0799_;
	wire _0800_;
	wire _0801_;
	wire _0802_;
	wire _0803_;
	wire _0804_;
	wire _0805_;
	wire _0806_;
	wire _0807_;
	wire _0808_;
	wire _0809_;
	wire _0810_;
	wire _0811_;
	wire _0812_;
	wire _0813_;
	wire _0814_;
	wire _0815_;
	wire _0816_;
	wire _0817_;
	wire _0818_;
	wire _0819_;
	wire _0820_;
	wire _0821_;
	wire _0822_;
	wire _0823_;
	wire _0824_;
	wire _0825_;
	wire _0826_;
	wire _0827_;
	wire _0828_;
	wire _0829_;
	wire _0830_;
	wire _0831_;
	wire _0832_;
	wire _0833_;
	wire _0834_;
	wire _0835_;
	wire _0836_;
	wire _0837_;
	wire _0838_;
	wire _0839_;
	wire _0840_;
	wire _0841_;
	wire _0842_;
	wire _0843_;
	wire _0844_;
	wire _0845_;
	wire _0846_;
	wire _0847_;
	wire _0848_;
	wire _0849_;
	wire _0850_;
	wire _0851_;
	wire _0852_;
	wire _0853_;
	wire _0854_;
	wire _0855_;
	wire _0856_;
	wire _0857_;
	wire _0858_;
	wire _0859_;
	wire _0860_;
	wire _0861_;
	wire _0862_;
	wire _0863_;
	wire _0864_;
	wire _0865_;
	wire _0866_;
	wire _0867_;
	wire _0868_;
	wire _0869_;
	wire _0870_;
	wire _0871_;
	wire _0872_;
	wire _0873_;
	wire _0874_;
	wire _0875_;
	wire _0876_;
	wire _0877_;
	wire _0878_;
	wire _0879_;
	wire _0880_;
	wire _0881_;
	wire _0882_;
	wire _0883_;
	wire _0884_;
	wire _0885_;
	wire _0886_;
	wire _0887_;
	wire _0888_;
	wire _0889_;
	wire _0890_;
	wire _0891_;
	wire _0892_;
	wire _0893_;
	wire _0894_;
	wire _0895_;
	wire _0896_;
	wire _0897_;
	wire _0898_;
	wire _0899_;
	wire _0900_;
	wire _0901_;
	wire _0902_;
	wire _0903_;
	wire _0904_;
	wire _0905_;
	wire _0906_;
	wire _0907_;
	wire _0908_;
	wire _0909_;
	wire _0910_;
	wire _0911_;
	wire _0912_;
	wire _0913_;
	wire _0914_;
	wire _0915_;
	wire _0916_;
	wire _0917_;
	wire _0918_;
	wire _0919_;
	wire _0920_;
	wire _0921_;
	wire _0922_;
	wire _0923_;
	wire _0924_;
	wire _0925_;
	wire _0926_;
	wire _0927_;
	wire _0928_;
	wire _0929_;
	wire _0930_;
	wire _0931_;
	wire _0932_;
	wire _0933_;
	wire _0934_;
	wire _0935_;
	wire _0936_;
	wire _0937_;
	wire _0938_;
	wire _0939_;
	wire _0940_;
	wire _0941_;
	wire _0942_;
	wire _0943_;
	wire _0944_;
	wire _0945_;
	wire _0946_;
	wire _0947_;
	wire _0948_;
	wire _0949_;
	wire _0950_;
	wire _0951_;
	wire _0952_;
	wire _0953_;
	wire _0954_;
	wire _0955_;
	wire _0956_;
	wire _0957_;
	wire _0958_;
	wire _0959_;
	wire _0960_;
	wire _0961_;
	wire _0962_;
	wire _0963_;
	wire _0964_;
	wire _0965_;
	wire _0966_;
	wire _0967_;
	wire _0968_;
	wire _0969_;
	wire _0970_;
	wire _0971_;
	wire _0972_;
	wire _0973_;
	wire _0974_;
	wire _0975_;
	wire _0976_;
	wire _0977_;
	wire _0978_;
	wire _0979_;
	wire _0980_;
	wire _0981_;
	wire _0982_;
	wire _0983_;
	wire _0984_;
	wire _0985_;
	wire _0986_;
	wire _0987_;
	wire _0988_;
	wire _0989_;
	wire _0990_;
	wire _0991_;
	wire _0992_;
	wire _0993_;
	wire _0994_;
	wire _0995_;
	wire _0996_;
	wire _0997_;
	wire _0998_;
	wire _0999_;
	wire _1000_;
	wire _1001_;
	wire _1002_;
	wire _1003_;
	wire _1004_;
	wire _1005_;
	wire _1006_;
	wire _1007_;
	wire _1008_;
	wire _1009_;
	wire _1010_;
	wire _1011_;
	wire _1012_;
	wire _1013_;
	wire _1014_;
	wire _1015_;
	wire _1016_;
	wire _1017_;
	wire _1018_;
	wire _1019_;
	wire _1020_;
	wire _1021_;
	wire _1022_;
	wire _1023_;
	wire _1024_;
	wire _1025_;
	wire _1026_;
	wire _1027_;
	wire _1028_;
	wire _1029_;
	wire _1030_;
	wire _1031_;
	wire _1032_;
	wire _1033_;
	wire _1034_;
	wire _1035_;
	wire _1036_;
	wire _1037_;
	wire _1038_;
	wire _1039_;
	wire _1040_;
	wire _1041_;
	wire _1042_;
	wire _1043_;
	wire _1044_;
	wire _1045_;
	wire _1046_;
	wire _1047_;
	wire _1048_;
	wire _1049_;
	wire _1050_;
	wire _1051_;
	wire _1052_;
	wire _1053_;
	wire _1054_;
	wire _1055_;
	wire _1056_;
	wire _1057_;
	wire _1058_;
	wire _1059_;
	wire _1060_;
	wire _1061_;
	wire _1062_;
	wire _1063_;
	wire _1064_;
	wire _1065_;
	wire _1066_;
	wire _1067_;
	wire _1068_;
	wire _1069_;
	wire _1070_;
	wire _1071_;
	wire _1072_;
	wire _1073_;
	wire _1074_;
	wire _1075_;
	wire _1076_;
	wire _1077_;
	wire _1078_;
	wire _1079_;
	wire _1080_;
	wire _1081_;
	wire _1082_;
	wire _1083_;
	wire _1084_;
	wire _1085_;
	wire _1086_;
	wire _1087_;
	wire _1088_;
	wire _1089_;
	wire _1090_;
	wire _1091_;
	wire _1092_;
	wire _1093_;
	wire _1094_;
	wire _1095_;
	wire _1096_;
	wire _1097_;
	wire _1098_;
	wire _1099_;
	wire _1100_;
	wire _1101_;
	wire _1102_;
	wire _1103_;
	wire _1104_;
	wire _1105_;
	wire _1106_;
	wire _1107_;
	wire _1108_;
	wire _1109_;
	wire _1110_;
	wire _1111_;
	wire _1112_;
	wire _1113_;
	wire _1114_;
	wire _1115_;
	wire _1116_;
	wire _1117_;
	wire _1118_;
	wire _1119_;
	wire _1120_;
	wire _1121_;
	wire _1122_;
	wire _1123_;
	wire _1124_;
	wire _1125_;
	wire _1126_;
	wire _1127_;
	wire _1128_;
	wire _1129_;
	wire _1130_;
	wire _1131_;
	wire _1132_;
	wire _1133_;
	wire _1134_;
	wire _1135_;
	wire _1136_;
	wire _1137_;
	wire _1138_;
	wire _1139_;
	wire _1140_;
	wire _1141_;
	wire _1142_;
	wire _1143_;
	wire _1144_;
	wire _1145_;
	wire _1146_;
	wire _1147_;
	wire _1148_;
	wire _1149_;
	wire _1150_;
	wire _1151_;
	wire _1152_;
	wire _1153_;
	wire _1154_;
	wire _1155_;
	wire _1156_;
	wire _1157_;
	wire _1158_;
	wire _1159_;
	wire _1160_;
	wire _1161_;
	wire _1162_;
	wire _1163_;
	wire _1164_;
	wire _1165_;
	wire _1166_;
	wire _1167_;
	wire _1168_;
	wire _1169_;
	wire _1170_;
	wire _1171_;
	wire _1172_;
	wire _1173_;
	wire _1174_;
	wire _1175_;
	wire _1176_;
	wire _1177_;
	wire _1178_;
	wire _1179_;
	wire _1180_;
	wire _1181_;
	wire _1182_;
	wire _1183_;
	wire _1184_;
	wire _1185_;
	wire _1186_;
	wire _1187_;
	wire _1188_;
	wire _1189_;
	wire _1190_;
	wire _1191_;
	wire _1192_;
	wire _1193_;
	wire _1194_;
	wire _1195_;
	wire _1196_;
	wire _1197_;
	wire _1198_;
	wire _1199_;
	wire _1200_;
	wire _1201_;
	wire _1202_;
	wire _1203_;
	wire _1204_;
	wire _1205_;
	wire _1206_;
	wire _1207_;
	wire _1208_;
	wire _1209_;
	wire _1210_;
	wire _1211_;
	wire _1212_;
	wire _1213_;
	wire _1214_;
	wire _1215_;
	wire _1216_;
	wire _1217_;
	wire _1218_;
	wire _1219_;
	wire _1220_;
	wire _1221_;
	wire _1222_;
	wire _1223_;
	wire _1224_;
	wire _1225_;
	wire _1226_;
	wire _1227_;
	wire _1228_;
	wire _1229_;
	wire _1230_;
	wire _1231_;
	wire _1232_;
	wire _1233_;
	wire _1234_;
	wire _1235_;
	wire _1236_;
	wire _1237_;
	wire _1238_;
	wire _1239_;
	wire _1240_;
	wire _1241_;
	wire _1242_;
	wire _1243_;
	wire _1244_;
	wire _1245_;
	wire _1246_;
	wire _1247_;
	wire _1248_;
	wire _1249_;
	wire _1250_;
	wire _1251_;
	wire _1252_;
	wire _1253_;
	wire _1254_;
	wire _1255_;
	wire _1256_;
	wire _1257_;
	wire _1258_;
	wire _1259_;
	wire _1260_;
	wire _1261_;
	wire _1262_;
	wire _1263_;
	wire _1264_;
	wire _1265_;
	wire _1266_;
	wire _1267_;
	wire _1268_;
	wire _1269_;
	wire _1270_;
	wire _1271_;
	wire _1272_;
	wire _1273_;
	wire _1274_;
	wire _1275_;
	wire _1276_;
	wire _1277_;
	wire _1278_;
	wire _1279_;
	wire _1280_;
	wire _1281_;
	wire _1282_;
	wire _1283_;
	wire _1284_;
	wire _1285_;
	wire _1286_;
	wire _1287_;
	wire _1288_;
	wire _1289_;
	wire _1290_;
	wire _1291_;
	wire _1292_;
	wire _1293_;
	wire _1294_;
	wire _1295_;
	wire _1296_;
	wire _1297_;
	wire _1298_;
	wire _1299_;
	wire _1300_;
	wire _1301_;
	wire _1302_;
	wire _1303_;
	wire _1304_;
	wire _1305_;
	wire _1306_;
	wire _1307_;
	wire _1308_;
	wire _1309_;
	wire _1310_;
	wire _1311_;
	wire _1312_;
	wire _1313_;
	wire _1314_;
	wire _1315_;
	wire _1316_;
	wire _1317_;
	wire _1318_;
	wire _1319_;
	wire _1320_;
	wire _1321_;
	wire _1322_;
	wire _1323_;
	wire _1324_;
	wire _1325_;
	wire _1326_;
	wire _1327_;
	wire _1328_;
	wire _1329_;
	wire _1330_;
	wire _1331_;
	wire _1332_;
	wire _1333_;
	wire _1334_;
	wire _1335_;
	wire _1336_;
	wire _1337_;
	wire _1338_;
	wire _1339_;
	wire _1340_;
	wire _1341_;
	wire _1342_;
	wire _1343_;
	wire _1344_;
	wire _1345_;
	wire _1346_;
	wire _1347_;
	wire _1348_;
	wire _1349_;
	wire _1350_;
	wire _1351_;
	wire _1352_;
	wire _1353_;
	wire _1354_;
	wire _1355_;
	wire _1356_;
	wire _1357_;
	wire _1358_;
	wire _1359_;
	wire _1360_;
	wire _1361_;
	wire _1362_;
	wire _1363_;
	wire _1364_;
	wire _1365_;
	wire _1366_;
	wire _1367_;
	wire _1368_;
	wire _1369_;
	wire _1370_;
	wire _1371_;
	wire _1372_;
	wire _1373_;
	wire _1374_;
	wire _1375_;
	wire _1376_;
	wire _1377_;
	wire _1378_;
	wire _1379_;
	wire _1380_;
	wire _1381_;
	wire _1382_;
	wire _1383_;
	wire _1384_;
	wire _1385_;
	wire _1386_;
	wire _1387_;
	wire _1388_;
	wire _1389_;
	wire _1390_;
	wire _1391_;
	wire _1392_;
	wire _1393_;
	wire _1394_;
	wire _1395_;
	wire _1396_;
	wire _1397_;
	wire _1398_;
	wire _1399_;
	wire _1400_;
	wire _1401_;
	wire _1402_;
	wire _1403_;
	wire _1404_;
	wire _1405_;
	wire _1406_;
	wire _1407_;
	wire _1408_;
	wire _1409_;
	wire _1410_;
	wire _1411_;
	wire _1412_;
	wire _1413_;
	wire _1414_;
	wire _1415_;
	wire _1416_;
	wire _1417_;
	wire _1418_;
	wire _1419_;
	wire _1420_;
	wire _1421_;
	wire _1422_;
	wire _1423_;
	wire _1424_;
	wire _1425_;
	wire _1426_;
	wire _1427_;
	wire _1428_;
	wire _1429_;
	wire _1430_;
	wire _1431_;
	wire _1432_;
	wire _1433_;
	wire _1434_;
	wire _1435_;
	wire _1436_;
	wire _1437_;
	wire _1438_;
	wire _1439_;
	wire _1440_;
	wire _1441_;
	wire _1442_;
	wire _1443_;
	wire _1444_;
	wire _1445_;
	wire _1446_;
	wire _1447_;
	wire _1448_;
	wire _1449_;
	wire _1450_;
	wire _1451_;
	wire _1452_;
	wire _1453_;
	wire _1454_;
	wire _1455_;
	wire _1456_;
	wire _1457_;
	wire _1458_;
	wire _1459_;
	wire _1460_;
	wire _1461_;
	wire _1462_;
	wire _1463_;
	wire _1464_;
	wire _1465_;
	wire _1466_;
	wire _1467_;
	wire _1468_;
	wire _1469_;
	wire _1470_;
	wire _1471_;
	wire _1472_;
	wire _1473_;
	wire _1474_;
	wire _1475_;
	wire _1476_;
	wire _1477_;
	wire _1478_;
	wire _1479_;
	wire _1480_;
	wire _1481_;
	wire _1482_;
	wire _1483_;
	wire _1484_;
	wire _1485_;
	wire _1486_;
	wire _1487_;
	wire _1488_;
	wire _1489_;
	wire _1490_;
	wire _1491_;
	wire _1492_;
	wire _1493_;
	wire _1494_;
	wire _1495_;
	wire _1496_;
	wire _1497_;
	wire _1498_;
	wire _1499_;
	wire _1500_;
	wire _1501_;
	wire _1502_;
	wire _1503_;
	wire _1504_;
	wire _1505_;
	wire _1506_;
	wire _1507_;
	wire _1508_;
	wire _1509_;
	wire _1510_;
	wire _1511_;
	wire _1512_;
	wire _1513_;
	wire _1514_;
	wire _1515_;
	wire _1516_;
	wire _1517_;
	wire _1518_;
	wire _1519_;
	wire _1520_;
	wire _1521_;
	wire _1522_;
	wire _1523_;
	wire _1524_;
	wire _1525_;
	wire _1526_;
	wire _1527_;
	wire _1528_;
	wire _1529_;
	wire _1530_;
	wire _1531_;
	wire _1532_;
	wire _1533_;
	wire _1534_;
	wire _1535_;
	wire _1536_;
	wire _1537_;
	wire _1538_;
	wire _1539_;
	wire _1540_;
	wire _1541_;
	wire _1542_;
	wire _1543_;
	wire _1544_;
	wire _1545_;
	wire _1546_;
	wire _1547_;
	wire _1548_;
	wire _1549_;
	wire _1550_;
	wire _1551_;
	wire _1552_;
	wire _1553_;
	wire _1554_;
	wire _1555_;
	wire _1556_;
	wire _1557_;
	wire _1558_;
	wire _1559_;
	wire _1560_;
	wire _1561_;
	wire _1562_;
	wire _1563_;
	wire _1564_;
	wire _1565_;
	wire _1566_;
	wire _1567_;
	wire _1568_;
	wire _1569_;
	wire _1570_;
	wire _1571_;
	wire _1572_;
	wire _1573_;
	wire _1574_;
	wire _1575_;
	wire _1576_;
	wire _1577_;
	wire _1578_;
	wire _1579_;
	wire _1580_;
	wire _1581_;
	wire _1582_;
	wire _1583_;
	wire _1584_;
	wire _1585_;
	wire _1586_;
	wire _1587_;
	wire _1588_;
	wire _1589_;
	wire _1590_;
	wire _1591_;
	wire _1592_;
	wire _1593_;
	wire _1594_;
	wire _1595_;
	wire _1596_;
	wire _1597_;
	wire _1598_;
	wire _1599_;
	wire _1600_;
	wire _1601_;
	wire _1602_;
	wire _1603_;
	wire _1604_;
	wire _1605_;
	wire _1606_;
	wire _1607_;
	wire _1608_;
	wire _1609_;
	wire _1610_;
	wire _1611_;
	wire _1612_;
	wire _1613_;
	wire _1614_;
	wire _1615_;
	wire _1616_;
	wire _1617_;
	wire _1618_;
	wire _1619_;
	wire _1620_;
	wire _1621_;
	wire _1622_;
	wire _1623_;
	wire _1624_;
	wire _1625_;
	wire _1626_;
	wire _1627_;
	wire _1628_;
	wire _1629_;
	wire _1630_;
	wire _1631_;
	wire _1632_;
	wire _1633_;
	wire _1634_;
	wire _1635_;
	wire _1636_;
	wire _1637_;
	wire _1638_;
	wire _1639_;
	wire _1640_;
	wire _1641_;
	wire _1642_;
	wire _1643_;
	wire _1644_;
	wire _1645_;
	wire _1646_;
	wire _1647_;
	wire _1648_;
	wire _1649_;
	wire _1650_;
	wire _1651_;
	wire _1652_;
	wire _1653_;
	wire _1654_;
	wire _1655_;
	wire _1656_;
	wire _1657_;
	wire _1658_;
	wire _1659_;
	wire _1660_;
	wire _1661_;
	wire _1662_;
	wire _1663_;
	wire _1664_;
	wire _1665_;
	wire _1666_;
	wire _1667_;
	wire _1668_;
	wire _1669_;
	wire _1670_;
	wire _1671_;
	wire _1672_;
	wire _1673_;
	wire _1674_;
	wire _1675_;
	wire _1676_;
	wire _1677_;
	wire _1678_;
	wire _1679_;
	wire _1680_;
	wire _1681_;
	wire _1682_;
	wire _1683_;
	wire _1684_;
	wire _1685_;
	wire _1686_;
	wire _1687_;
	wire _1688_;
	wire _1689_;
	wire _1690_;
	wire _1691_;
	wire _1692_;
	wire _1693_;
	wire _1694_;
	wire _1695_;
	wire _1696_;
	wire _1697_;
	wire _1698_;
	wire _1699_;
	wire _1700_;
	wire _1701_;
	wire _1702_;
	wire _1703_;
	wire _1704_;
	wire _1705_;
	wire _1706_;
	wire _1707_;
	wire _1708_;
	wire _1709_;
	wire _1710_;
	wire _1711_;
	wire _1712_;
	wire _1713_;
	wire _1714_;
	wire _1715_;
	wire _1716_;
	wire _1717_;
	wire _1718_;
	wire _1719_;
	wire _1720_;
	wire _1721_;
	wire _1722_;
	wire _1723_;
	wire _1724_;
	wire _1725_;
	wire _1726_;
	wire _1727_;
	wire _1728_;
	wire _1729_;
	wire _1730_;
	wire _1731_;
	wire _1732_;
	wire _1733_;
	wire _1734_;
	wire _1735_;
	wire _1736_;
	wire _1737_;
	wire _1738_;
	wire _1739_;
	wire _1740_;
	wire _1741_;
	wire _1742_;
	wire _1743_;
	wire _1744_;
	wire _1745_;
	wire _1746_;
	wire _1747_;
	wire _1748_;
	wire _1749_;
	wire _1750_;
	wire _1751_;
	wire _1752_;
	wire _1753_;
	wire _1754_;
	wire _1755_;
	wire _1756_;
	wire _1757_;
	wire _1758_;
	wire _1759_;
	wire _1760_;
	wire _1761_;
	wire _1762_;
	wire _1763_;
	wire _1764_;
	wire _1765_;
	wire _1766_;
	wire _1767_;
	wire _1768_;
	wire _1769_;
	wire _1770_;
	wire _1771_;
	wire _1772_;
	wire _1773_;
	wire _1774_;
	wire _1775_;
	wire _1776_;
	wire _1777_;
	wire _1778_;
	wire _1779_;
	wire _1780_;
	wire _1781_;
	wire _1782_;
	wire _1783_;
	wire _1784_;
	wire _1785_;
	wire _1786_;
	wire _1787_;
	wire _1788_;
	wire _1789_;
	wire _1790_;
	wire _1791_;
	wire _1792_;
	wire _1793_;
	wire _1794_;
	wire _1795_;
	wire _1796_;
	wire _1797_;
	wire _1798_;
	wire _1799_;
	wire _1800_;
	wire _1801_;
	wire _1802_;
	wire _1803_;
	wire _1804_;
	wire _1805_;
	wire _1806_;
	wire _1807_;
	wire _1808_;
	wire _1809_;
	wire _1810_;
	wire _1811_;
	wire _1812_;
	wire _1813_;
	wire _1814_;
	wire _1815_;
	wire _1816_;
	wire _1817_;
	wire _1818_;
	wire _1819_;
	wire _1820_;
	wire _1821_;
	wire _1822_;
	wire _1823_;
	wire _1824_;
	wire _1825_;
	wire _1826_;
	wire _1827_;
	wire _1828_;
	wire _1829_;
	wire _1830_;
	wire _1831_;
	wire _1832_;
	wire _1833_;
	wire _1834_;
	wire _1835_;
	wire _1836_;
	wire _1837_;
	wire _1838_;
	wire _1839_;
	wire _1840_;
	wire _1841_;
	wire _1842_;
	wire _1843_;
	wire _1844_;
	wire _1845_;
	wire _1846_;
	wire _1847_;
	wire _1848_;
	wire _1849_;
	wire _1850_;
	wire _1851_;
	wire _1852_;
	wire _1853_;
	wire _1854_;
	wire _1855_;
	wire _1856_;
	wire _1857_;
	wire _1858_;
	wire _1859_;
	wire _1860_;
	wire _1861_;
	wire _1862_;
	wire _1863_;
	wire _1864_;
	wire _1865_;
	wire _1866_;
	wire _1867_;
	wire _1868_;
	wire _1869_;
	wire _1870_;
	wire _1871_;
	wire _1872_;
	wire _1873_;
	wire _1874_;
	wire _1875_;
	wire _1876_;
	wire _1877_;
	wire _1878_;
	wire _1879_;
	wire _1880_;
	wire _1881_;
	wire _1882_;
	wire _1883_;
	wire _1884_;
	wire _1885_;
	wire _1886_;
	wire _1887_;
	wire _1888_;
	wire [3:0] _1889_;
	wire [3:0] _1890_;
	input wire [13:0] io_in;
	output wire [13:0] io_out;
	wire \mchip.M1.ACK ;
	wire [6:0] \mchip.M1.ADDR.addr ;
	wire [1:0] \mchip.M1.ADDR.addr_sel ;
	wire [6:0] \mchip.M1.ADDR.data_in ;
	wire \mchip.M1.COUNT.clear ;
	wire \mchip.M1.COUNT.clock ;
	wire [3:0] \mchip.M1.COUNT.count ;
	wire \mchip.M1.COUNT.en ;
	wire \mchip.M1.IN_REG.SCL_posedge ;
	wire \mchip.M1.IN_REG.SDA ;
	wire [7:0] \mchip.M1.IN_REG.SHIFT.Q ;
	wire \mchip.M1.IN_REG.SHIFT.clock ;
	wire \mchip.M1.IN_REG.SHIFT.en ;
	wire \mchip.M1.IN_REG.SHIFT.reset ;
	wire \mchip.M1.IN_REG.SHIFT.serial ;
	wire \mchip.M1.IN_REG.clock ;
	wire [7:0] \mchip.M1.IN_REG.data_in ;
	wire \mchip.M1.IN_REG.reset ;
	wire \mchip.M1.M.ACK ;
	wire \mchip.M1.M.SCL_negedge ;
	wire \mchip.M1.M.clear_counter ;
	wire \mchip.M1.M.clock ;
	wire [11:0] \mchip.M1.M.currState ;
	wire [7:0] \mchip.M1.M.data_in ;
	wire \mchip.M1.M.out_en ;
	wire \mchip.M1.M.read_write ;
	wire \mchip.M1.M.reg_sel_en ;
	wire \mchip.M1.M.reset ;
	wire \mchip.M1.MEM.SCL_negedge ;
	wire \mchip.M1.MEM.clock ;
	wire [2:0] \mchip.M1.MEM.count ;
	wire [7:0] \mchip.M1.MEM.data_in ;
	reg [2:0] \mchip.M1.MEM.index ;
	wire [31:0] \mchip.M1.MEM.j ;
	wire [7:0] \mchip.M1.MEM.parallel_in ;
	reg [7:0] \mchip.M1.MEM.parallel_in_temp ;
	wire [7:0] \mchip.M1.MEM.reg_out ;
	reg [7:0] \mchip.M1.MEM.registers[0] ;
	wire [7:0] \mchip.M1.MEM.registers[1] ;
	wire [191:0] \mchip.M1.MEM.registers_packed ;
	wire \mchip.M1.MEM.reset ;
	wire \mchip.M1.OUT.out_en ;
	reg \mchip.M1.READ_ACK.ACK ;
	wire \mchip.M1.READ_ACK.SCL_posedge ;
	wire \mchip.M1.READ_ACK.SDA ;
	wire \mchip.M1.READ_ACK.clock ;
	wire \mchip.M1.REG.SCL_negedge ;
	wire \mchip.M1.REG.clock ;
	wire \mchip.M1.REG.en ;
	wire \mchip.M1.REG.reset ;
	wire [4:0] \mchip.M1.REG.sel_in ;
	wire \mchip.M1.S1.EDGE.clock ;
	reg \mchip.M1.S1.EDGE.prev ;
	wire \mchip.M1.S1.EDGE.sig ;
	reg \mchip.M1.S1.EDGE.sig_negedge ;
	wire \mchip.M1.S1.EDGE.sig_out ;
	reg \mchip.M1.S1.EDGE.sig_posedge ;
	wire \mchip.M1.S1.async ;
	wire \mchip.M1.S1.clock ;
	wire \mchip.M1.S1.m1.D ;
	reg \mchip.M1.S1.m1.Q ;
	wire \mchip.M1.S1.m1.clock ;
	wire \mchip.M1.S1.sig_negedge ;
	wire \mchip.M1.S1.sig_posedge ;
	wire \mchip.M1.S1.sync ;
	wire \mchip.M1.S1.temp ;
	wire \mchip.M1.S2.EDGE.clock ;
	reg \mchip.M1.S2.EDGE.prev ;
	wire \mchip.M1.S2.EDGE.sig ;
	reg \mchip.M1.S2.EDGE.sig_negedge ;
	wire \mchip.M1.S2.EDGE.sig_out ;
	reg \mchip.M1.S2.EDGE.sig_posedge ;
	wire \mchip.M1.S2.async ;
	wire \mchip.M1.S2.clock ;
	wire \mchip.M1.S2.m1.D ;
	reg \mchip.M1.S2.m1.Q ;
	wire \mchip.M1.S2.m1.clock ;
	wire \mchip.M1.S2.sig_negedge ;
	wire \mchip.M1.S2.sig_posedge ;
	wire \mchip.M1.S2.sync ;
	wire \mchip.M1.S2.temp ;
	wire \mchip.M1.SCL_in ;
	wire \mchip.M1.SCL_negedge ;
	wire \mchip.M1.SCL_posedge ;
	wire \mchip.M1.SCL_sync ;
	wire \mchip.M1.SDA_in ;
	wire \mchip.M1.SDA_negedge ;
	wire \mchip.M1.SDA_posedge ;
	wire \mchip.M1.SDA_sync ;
	wire \mchip.M1.START.SCL ;
	wire \mchip.M1.START.SDA_negedge ;
	wire \mchip.M1.START.clear_start ;
	wire \mchip.M1.START.clock ;
	wire \mchip.M1.STOP.SCL ;
	wire \mchip.M1.STOP.SDA_posedge ;
	wire \mchip.M1.STOP.clear_stop ;
	wire \mchip.M1.STOP.clock ;
	wire [1:0] \mchip.M1.addr_sel ;
	wire \mchip.M1.clear_counter ;
	wire \mchip.M1.clock ;
	wire [3:0] \mchip.M1.count ;
	wire [7:0] \mchip.M1.data_in ;
	wire \mchip.M1.out_en ;
	wire [7:0] \mchip.M1.parallel_in ;
	wire [7:0] \mchip.M1.reg_out ;
	wire \mchip.M1.reg_sel_en ;
	wire [191:0] \mchip.M1.registers_packed ;
	wire \mchip.M1.reset ;
	wire \mchip.M2.PWM1 ;
	wire \mchip.M2.PWM2 ;
	wire \mchip.M2.PWM_DRIVER.P1.PWM_out ;
	wire \mchip.M2.PWM_DRIVER.P1.clock ;
	wire \mchip.M2.PWM_DRIVER.P1.reset ;
	wire \mchip.M2.PWM_DRIVER.P2.PWM_out ;
	wire \mchip.M2.PWM_DRIVER.P2.clock ;
	wire \mchip.M2.PWM_DRIVER.P2.reset ;
	wire \mchip.M2.PWM_DRIVER.PWM1 ;
	wire \mchip.M2.PWM_DRIVER.PWM2 ;
	wire \mchip.M2.PWM_DRIVER.clock ;
	wire [191:0] \mchip.M2.PWM_DRIVER.registers_packed ;
	wire \mchip.M2.PWM_DRIVER.reset ;
	wire \mchip.M2.UART_DRIVER.clock ;
	wire [7:0] \mchip.M2.UART_DRIVER.data ;
	wire [15:0] \mchip.M2.UART_DRIVER.frame ;
	wire \mchip.M2.UART_DRIVER.reset ;
	wire \mchip.M2.UART_DRIVER.tx ;
	wire \mchip.M2.clock ;
	wire [10:0] \mchip.M2.data_out ;
	wire [7:0] \mchip.M2.reg_out ;
	wire [191:0] \mchip.M2.registers_packed ;
	wire \mchip.M2.reset ;
	wire \mchip.M2.tx ;
	wire \mchip.SCL_in ;
	wire \mchip.SDA_in ;
	wire \mchip.SDA_out ;
	wire \mchip.clock ;
	wire [10:0] \mchip.data_out ;
	wire [11:0] \mchip.io_in ;
	wire [11:0] \mchip.io_out ;
	wire [7:0] \mchip.reg_out ;
	wire [191:0] \mchip.registers_packed ;
	wire \mchip.reset ;
	assign _1404_ = _0131_ & ~io_in[13];
	assign _1405_ = _0127_ & ~io_in[13];
	assign _1406_ = _0130_ & ~io_in[13];
	assign _1407_ = _1406_ | _1405_;
	assign \mchip.M1.START.clear_start  = _1407_ | io_in[13];
	assign _1408_ = _0192_ & ~\mchip.M1.START.clear_start ;
	assign _1409_ = _1408_ & _1404_;
	assign _1410_ = _0126_ & ~io_in[13];
	assign _1411_ = _0125_ & ~io_in[13];
	assign _1412_ = _1411_ | _1410_;
	assign _1413_ = _0124_ & ~io_in[13];
	assign _1414_ = _0123_ & ~io_in[13];
	assign _1415_ = _1414_ | _1413_;
	assign _1416_ = _1415_ | _1412_;
	assign _1417_ = _0128_ & ~io_in[13];
	assign _1418_ = _1417_ | _1416_;
	assign _1419_ = _1418_ | _1409_;
	assign _1420_ = ~(_1418_ | _1404_);
	assign \mchip.M1.COUNT.clear  = _1419_ & ~_1420_;
	assign \mchip.M1.COUNT.count [0] = _0193_ & ~\mchip.M1.COUNT.clear ;
	assign _1889_[0] = ~\mchip.M1.COUNT.count [0];
	assign \mchip.M1.COUNT.count [1] = _0194_ & ~\mchip.M1.COUNT.clear ;
	assign \mchip.M1.COUNT.count [2] = _0195_ & ~\mchip.M1.COUNT.clear ;
	assign _1421_ = \mchip.M1.COUNT.clear  | ~_0196_;
	assign _1422_ = _1421_ | \mchip.M1.COUNT.count [2];
	assign _1423_ = \mchip.M1.COUNT.count [1] | \mchip.M1.COUNT.count [0];
	assign _1424_ = _1423_ | _1422_;
	assign _1425_ = _1424_ | ~_1404_;
	assign _1426_ = \mchip.M1.S1.EDGE.sig_negedge  & ~_1425_;
	assign _1427_ = io_in[13] | ~_0191_;
	assign _1428_ = _0187_ & ~io_in[13];
	assign _1429_ = _0188_ & ~io_in[13];
	assign _1430_ = _1429_ | _1428_;
	assign _1431_ = _0190_ & ~io_in[13];
	assign _1432_ = _0189_ & ~io_in[13];
	assign _1433_ = _1432_ | _1431_;
	assign _1434_ = _1433_ | _1430_;
	assign _1435_ = _1427_ & ~_1434_;
	assign _1436_ = _1426_ & ~_1435_;
	assign _1437_ = _1428_ | ~_1429_;
	assign _1438_ = _1437_ | _1433_;
	assign _1439_ = ~(_1438_ | _1427_);
	assign _0016_ = _1439_ & _1436_;
	assign _1440_ = _0328_ & ~io_in[13];
	assign _1441_ = _0182_ & ~io_in[13];
	assign _1442_ = _1440_ | ~_1441_;
	assign _1443_ = _1441_ ^ _1440_;
	assign _1444_ = _0327_ & ~io_in[13];
	assign _1445_ = _0181_ & ~io_in[13];
	assign _1446_ = _1445_ & ~_1444_;
	assign _1447_ = _1446_ & ~_1443_;
	assign _1448_ = _1442_ & ~_1447_;
	assign _1449_ = _0326_ & ~io_in[13];
	assign _1450_ = _0180_ & ~io_in[13];
	assign _1451_ = _1450_ & ~_1449_;
	assign _1452_ = _0179_ & ~io_in[13];
	assign _1453_ = _0325_ & ~io_in[13];
	assign _1454_ = _1452_ | ~_1453_;
	assign _1455_ = _1450_ ^ _1449_;
	assign _1456_ = _1454_ & ~_1455_;
	assign _1457_ = _1456_ | _1451_;
	assign _1458_ = _1445_ ^ _1444_;
	assign _1459_ = _1458_ | _1443_;
	assign _1460_ = _1457_ & ~_1459_;
	assign _1461_ = _1448_ & ~_1460_;
	assign _1462_ = _0183_ & ~io_in[13];
	assign _1463_ = _0329_ & ~io_in[13];
	assign _1464_ = _1463_ ^ _1462_;
	assign _1465_ = _0184_ & ~io_in[13];
	assign _1466_ = _0330_ & ~io_in[13];
	assign _1467_ = _1466_ ^ _1465_;
	assign _1468_ = _1467_ | _1464_;
	assign _1469_ = _0186_ & ~io_in[13];
	assign _1470_ = _0332_ & ~io_in[13];
	assign _1471_ = ~(_1470_ ^ _1469_);
	assign _1472_ = _0185_ & ~io_in[13];
	assign _1473_ = _0331_ & ~io_in[13];
	assign _1474_ = _1473_ ^ _1472_;
	assign _1475_ = _1474_ | ~_1471_;
	assign _1476_ = _1475_ | _1468_;
	assign _1477_ = _1476_ | _1461_;
	assign _1478_ = _1466_ | ~_1465_;
	assign _1479_ = _1462_ & ~_1463_;
	assign _1480_ = _1479_ & ~_1467_;
	assign _1481_ = _1478_ & ~_1480_;
	assign _1482_ = ~(_1481_ | _1475_);
	assign _1483_ = _1473_ | ~_1472_;
	assign _1484_ = _1471_ & ~_1483_;
	assign _1485_ = _1469_ & ~_1470_;
	assign _1486_ = _1485_ | _1484_;
	assign _1487_ = _1486_ | _1482_;
	assign _1488_ = _1477_ & ~_1487_;
	assign _1489_ = _1453_ ^ _1452_;
	assign _1490_ = _1489_ | _1455_;
	assign _1491_ = _1490_ | _1459_;
	assign _1492_ = ~(_1491_ | _1476_);
	assign _0118_ = _1488_ & ~_1492_;
	assign _1493_ = _0177_ & ~io_in[13];
	assign _1494_ = _0292_ & ~io_in[13];
	assign _1495_ = ~(_1494_ ^ _1493_);
	assign _1496_ = _0176_ & ~io_in[13];
	assign _1497_ = _0291_ & ~io_in[13];
	assign _1498_ = _1497_ ^ _1496_;
	assign _1499_ = _1495_ & ~_1498_;
	assign _1500_ = _0174_ & ~io_in[13];
	assign _1501_ = _0289_ & ~io_in[13];
	assign _1502_ = _1501_ ^ _1500_;
	assign _1503_ = _0175_ & ~io_in[13];
	assign _1504_ = _0290_ & ~io_in[13];
	assign _1505_ = _1504_ ^ _1503_;
	assign _1506_ = _1505_ | _1502_;
	assign _1507_ = _1499_ & ~_1506_;
	assign _1508_ = _0288_ & ~io_in[13];
	assign _1509_ = _0173_ & ~io_in[13];
	assign _1510_ = _1508_ | ~_1509_;
	assign _1511_ = ~(_1509_ ^ _1508_);
	assign _1512_ = _0287_ & ~io_in[13];
	assign _1513_ = _0172_ & ~io_in[13];
	assign _1514_ = _1512_ | ~_1513_;
	assign _1515_ = _1511_ & ~_1514_;
	assign _1516_ = _1510_ & ~_1515_;
	assign _1517_ = _1513_ ^ _1512_;
	assign _1518_ = _1511_ & ~_1517_;
	assign _1519_ = _0286_ & ~io_in[13];
	assign _1520_ = _0171_ & ~io_in[13];
	assign _1521_ = _1519_ | ~_1520_;
	assign _1522_ = _0170_ & ~io_in[13];
	assign _1523_ = _0285_ & ~io_in[13];
	assign _1524_ = _1522_ | ~_1523_;
	assign _1525_ = _1520_ ^ _1519_;
	assign _1526_ = _1524_ & ~_1525_;
	assign _1527_ = _1521_ & ~_1526_;
	assign _1528_ = _1518_ & ~_1527_;
	assign _1529_ = _1516_ & ~_1528_;
	assign _1530_ = _1529_ | ~_1507_;
	assign _1531_ = _1504_ | ~_1503_;
	assign _1532_ = _1500_ & ~_1501_;
	assign _1533_ = _1532_ & ~_1505_;
	assign _1534_ = _1531_ & ~_1533_;
	assign _1535_ = _1499_ & ~_1534_;
	assign _1536_ = _1497_ | ~_1496_;
	assign _1537_ = _1495_ & ~_1536_;
	assign _1538_ = _1493_ & ~_1494_;
	assign _1539_ = _1538_ | _1537_;
	assign _1540_ = _1539_ | _1535_;
	assign _1541_ = _1530_ & ~_1540_;
	assign _1542_ = _1523_ ^ _1522_;
	assign _1543_ = ~(_1542_ | _1525_);
	assign _1544_ = ~(_1543_ & _1518_);
	assign _1545_ = _1507_ & ~_1544_;
	assign _0119_ = _1541_ & ~_1545_;
	assign \mchip.M1.M.read_write  = _0373_ & ~io_in[13];
	assign _1546_ = _0129_ & ~io_in[13];
	assign _1547_ = ~\mchip.M1.S1.EDGE.sig_negedge ;
	assign _1548_ = _1547_ & ~_1408_;
	assign \mchip.M1.STOP.clear_stop  = _0127_ | io_in[13];
	assign _1549_ = _0178_ & ~\mchip.M1.STOP.clear_stop ;
	assign _1550_ = _1548_ & ~_1549_;
	assign _1551_ = _1550_ & _1546_;
	assign _1552_ = _1549_ | \mchip.M1.M.read_write ;
	assign _1553_ = _1408_ | _1547_;
	assign _1554_ = _1553_ | _1552_;
	assign _1555_ = _1414_ & ~_1554_;
	assign _1556_ = _1549_ | ~_1424_;
	assign _1557_ = _1556_ | _1553_;
	assign _1558_ = _1546_ & ~_1557_;
	assign _1559_ = _1558_ | _1555_;
	assign _0008_ = _1559_ | _1551_;
	assign _1560_ = ~(_1429_ & _1428_);
	assign _1561_ = _1560_ | _1433_;
	assign _1562_ = ~(_1561_ | _1427_);
	assign _0015_ = _1562_ & _1436_;
	assign _1563_ = _1550_ & _1417_;
	assign _1564_ = _1549_ | _1424_;
	assign _1565_ = _1564_ | _1553_;
	assign _1566_ = _1404_ & ~_1565_;
	assign _0007_ = _1566_ | _1563_;
	assign _1567_ = _1431_ | ~_1432_;
	assign _1568_ = _1567_ | _1430_;
	assign _1569_ = ~(_1568_ | _1427_);
	assign _0014_ = _1569_ & _1436_;
	assign \mchip.M1.IN_REG.SHIFT.Q [1] = _0374_ & ~io_in[13];
	assign \mchip.M1.IN_REG.SHIFT.Q [2] = _0375_ & ~io_in[13];
	assign \mchip.M1.IN_REG.SHIFT.Q [4] = _0377_ & ~io_in[13];
	assign \mchip.M1.IN_REG.SHIFT.Q [3] = _0376_ & ~io_in[13];
	assign \mchip.M1.IN_REG.SHIFT.Q [5] = _0378_ & ~io_in[13];
	assign \mchip.M1.IN_REG.SHIFT.Q [6] = _0379_ & ~io_in[13];
	assign \mchip.M1.IN_REG.SHIFT.Q [7] = _0380_ & ~io_in[13];
	assign _1570_ = io_in[3] | ~io_in[2];
	assign _1571_ = io_in[2] & io_in[3];
	assign _1572_ = _1570_ & ~_1571_;
	assign _1573_ = ~(_1572_ ^ \mchip.M1.IN_REG.SHIFT.Q [1]);
	assign _1574_ = io_in[3] & ~io_in[2];
	assign _1575_ = _1574_ | _1571_;
	assign _1576_ = ~(io_in[2] | io_in[3]);
	assign _1577_ = _1575_ & ~_1576_;
	assign _1578_ = _1577_ ^ \mchip.M1.IN_REG.SHIFT.Q [2];
	assign _1579_ = ~(_1578_ | _1573_);
	assign _1580_ = \mchip.M1.IN_REG.SHIFT.Q [3] | \mchip.M1.IN_REG.SHIFT.Q [4];
	assign _1581_ = _1579_ & ~_1580_;
	assign _1582_ = \mchip.M1.IN_REG.SHIFT.Q [5] | ~\mchip.M1.IN_REG.SHIFT.Q [6];
	assign _1583_ = _1582_ | \mchip.M1.IN_REG.SHIFT.Q [7];
	assign _1584_ = _1581_ & ~_1583_;
	assign _1585_ = _1584_ | _1549_;
	assign _1586_ = _1585_ | _1553_;
	assign _1587_ = _1586_ | _1424_;
	assign _1588_ = _1406_ & ~_1587_;
	assign _1589_ = ~(_1549_ | _1408_);
	assign _1590_ = ~(_0121_ | io_in[13]);
	assign _1591_ = _1589_ & ~_1590_;
	assign _1592_ = _1591_ | _1549_;
	assign _0006_ = _1592_ | _1588_;
	assign _1593_ = _1550_ & _1410_;
	assign _1594_ = _1546_ & ~_1565_;
	assign _0005_ = _1594_ | _1593_;
	assign _1595_ = _0136_ & ~io_in[13];
	assign _1596_ = io_in[13] | ~_0137_;
	assign _1597_ = _1595_ & ~_1596_;
	assign _1598_ = _0135_ & ~io_in[13];
	assign _1599_ = _0134_ & ~io_in[13];
	assign _1600_ = ~(_1599_ | _1598_);
	assign _1601_ = _1600_ | ~_1597_;
	assign _1602_ = _0133_ & ~io_in[13];
	assign _1603_ = _0132_ & ~io_in[13];
	assign _1604_ = _1603_ & _1602_;
	assign _1605_ = ~(_1604_ & _1600_);
	assign _1606_ = _1597_ & ~_1605_;
	assign _0120_ = _1601_ & ~_1606_;
	assign _1607_ = _1429_ | ~_1428_;
	assign _1608_ = _1607_ | _1433_;
	assign _1609_ = ~(_1608_ | _1427_);
	assign _0017_ = _1609_ & _1436_;
	assign _1610_ = _1410_ & ~_1547_;
	assign _1611_ = ~(_1417_ | _1411_);
	assign _1612_ = \mchip.M1.S1.EDGE.sig_negedge  & ~_1611_;
	assign _1613_ = _1431_ & ~_1427_;
	assign _1614_ = ~_1432_;
	assign _1615_ = _1431_ | _1427_;
	assign _1616_ = _1615_ | _1560_;
	assign _1617_ = ~(_1616_ | _1614_);
	assign _0010_ = _1612_ | _1610_;
	assign \mchip.M2.UART_DRIVER.tx  = _0389_ & ~io_in[13];
	assign _1618_ = _0391_ & ~io_in[13];
	assign _1619_ = _0390_ & ~io_in[13];
	assign _1620_ = ~(_1619_ | _1618_);
	assign _1621_ = _0393_ & ~io_in[13];
	assign _1622_ = _0392_ & ~io_in[13];
	assign _1623_ = _1622_ | _1621_;
	assign _1624_ = _1620_ & ~_1623_;
	assign _1625_ = _0395_ & ~io_in[13];
	assign _1626_ = _0394_ & ~io_in[13];
	assign _1627_ = _1626_ | _1625_;
	assign _1628_ = _0397_ & ~io_in[13];
	assign _1629_ = _0396_ & ~io_in[13];
	assign _1630_ = _1629_ | _1628_;
	assign _1631_ = _1630_ | _1627_;
	assign _1632_ = _1624_ & ~_1631_;
	assign _1633_ = _0399_ | io_in[13];
	assign _1634_ = _0398_ | io_in[13];
	assign _1635_ = _1634_ | _1633_;
	assign _1636_ = _0401_ | io_in[13];
	assign _1637_ = _0400_ | io_in[13];
	assign _1638_ = _1637_ | _1636_;
	assign _1639_ = _1638_ | _1635_;
	assign _1640_ = _1632_ & ~_1639_;
	assign _1641_ = _0403_ | io_in[13];
	assign _1642_ = _0402_ | io_in[13];
	assign _1643_ = _1642_ | _1641_;
	assign _1644_ = _1640_ & ~_1643_;
	assign _1645_ = _0404_ | io_in[13];
	assign _1646_ = _1644_ & ~_1645_;
	assign _1647_ = \mchip.M2.UART_DRIVER.tx  & ~_1619_;
	assign _1648_ = _1622_ | _1618_;
	assign _1649_ = _1647_ & ~_1648_;
	assign _1650_ = _1629_ | _1625_;
	assign _1651_ = _1626_ | _1621_;
	assign _1652_ = _1651_ | _1650_;
	assign _1653_ = _1649_ & ~_1652_;
	assign _1654_ = _1645_ | _1641_;
	assign _1655_ = _1642_ | _1636_;
	assign _1656_ = _1655_ | _1654_;
	assign _1657_ = _1637_ | _1633_;
	assign _1658_ = _1634_ | _1628_;
	assign _1659_ = _1658_ | _1657_;
	assign _1660_ = _1659_ | _1656_;
	assign _1661_ = _1653_ & ~_1660_;
	assign _1662_ = ~(_1661_ | _1646_);
	assign _0035_ = ~_1662_;
	assign _1663_ = \mchip.M1.S1.EDGE.sig_negedge  & ~_1436_;
	assign _0034_ = _1663_ & ~io_in[13];
	assign _1664_ = _1427_ & ~_1608_;
	assign _0033_ = _1664_ & _1436_;
	assign _1665_ = _1427_ & ~_1438_;
	assign _0032_ = _1665_ & _1436_;
	assign _1666_ = _1427_ & ~_1561_;
	assign _0031_ = _1666_ & _1436_;
	assign _1667_ = _1427_ & ~_1568_;
	assign _0030_ = _1667_ & _1436_;
	assign _1668_ = _1607_ | _1567_;
	assign _1669_ = _1427_ & ~_1668_;
	assign _0029_ = _1669_ & _1436_;
	assign _1670_ = _1567_ | _1437_;
	assign _1671_ = _1670_ | ~_1427_;
	assign _0028_ = _1436_ & ~_1671_;
	assign _1672_ = _1549_ | ~\mchip.M1.READ_ACK.ACK ;
	assign _1673_ = _1672_ | _1553_;
	assign _1674_ = _1411_ & ~_1673_;
	assign _1675_ = io_in[13] | ~_0122_;
	assign _1676_ = ~(_1675_ | _1557_);
	assign _1677_ = _1676_ | _1674_;
	assign _1678_ = _1549_ | ~\mchip.M1.M.read_write ;
	assign _1679_ = _1678_ | _1553_;
	assign _1680_ = _1414_ & ~_1679_;
	assign _1681_ = _1550_ & ~_1675_;
	assign _1682_ = _1681_ | _1680_;
	assign _0002_ = _1682_ | _1677_;
	assign _1683_ = _1567_ | _1560_;
	assign _1684_ = _1427_ & ~_1683_;
	assign _0027_ = _1684_ & _1436_;
	assign _1685_ = _1432_ | ~_1431_;
	assign _1686_ = _1685_ | _1430_;
	assign _1687_ = _1427_ & ~_1686_;
	assign _0026_ = _1687_ & _1436_;
	assign _1688_ = _1550_ & _1406_;
	assign _1689_ = _1406_ & ~_1557_;
	assign _1690_ = _1408_ & ~_1549_;
	assign _1691_ = _1690_ | _1689_;
	assign _0009_ = _1691_ | _1688_;
	assign _1692_ = ~(_1413_ | _1405_);
	assign _1693_ = _1549_ | ~_1692_;
	assign _1694_ = ~(_1693_ | _1553_);
	assign _1695_ = ~(_1417_ | _1410_);
	assign _1696_ = _1694_ & ~_1695_;
	assign _1697_ = _1404_ & ~_1557_;
	assign _1698_ = _1550_ & _1404_;
	assign _1699_ = _1698_ | _1697_;
	assign _0001_ = _1699_ | _1696_;
	assign _1700_ = ~(_1434_ | _1427_);
	assign _0018_ = _1700_ & _1436_;
	assign _1701_ = ~(_1668_ | _1427_);
	assign _0013_ = _1701_ & _1436_;
	assign _1702_ = ~(_1432_ & _1431_);
	assign _1703_ = _1702_ | _1560_;
	assign _1704_ = _1427_ & ~_1703_;
	assign _0019_ = _1704_ & _1436_;
	assign _1705_ = _1702_ | _1437_;
	assign _1706_ = _1427_ & ~_1705_;
	assign _0020_ = _1706_ & _1436_;
	assign _1707_ = _1702_ | _1607_;
	assign _1708_ = _1427_ & ~_1707_;
	assign _0021_ = _1708_ & _1436_;
	assign _1709_ = _1702_ | _1430_;
	assign _1710_ = _1427_ & ~_1709_;
	assign _0022_ = _1710_ & _1436_;
	assign _1711_ = _1685_ | _1560_;
	assign _1712_ = _1711_ | ~_1427_;
	assign _0023_ = _1436_ & ~_1712_;
	assign _1713_ = _1685_ | _1437_;
	assign _1714_ = _1427_ & ~_1713_;
	assign _0024_ = _1714_ & _1436_;
	assign _1715_ = _1685_ | _1607_;
	assign _1716_ = _1427_ & ~_1715_;
	assign _0025_ = _1716_ & _1436_;
	assign _1717_ = _1550_ & _1411_;
	assign _1718_ = ~(_1675_ | _1565_);
	assign _0004_ = _1718_ | _1717_;
	assign _1719_ = ~(_1670_ | _1427_);
	assign _0012_ = _1719_ & _1436_;
	assign _1720_ = _1614_ | ~_1436_;
	assign _0011_ = ~(_1720_ | _1616_);
	assign _1721_ = _1549_ | ~_1584_;
	assign _1722_ = _1721_ | _1553_;
	assign _1723_ = _1722_ | _1424_;
	assign _1724_ = _1406_ & ~_1723_;
	assign _1725_ = _1550_ & _1414_;
	assign _0003_ = _1725_ | _1724_;
	assign _1726_ = _0316_ & ~io_in[13];
	assign _1727_ = _0153_ & ~io_in[13];
	assign _1728_ = _1726_ | ~_1727_;
	assign _1729_ = ~(_1727_ ^ _1726_);
	assign _1730_ = _0315_ & ~io_in[13];
	assign _1731_ = _0152_ & ~io_in[13];
	assign _1732_ = _1730_ | ~_1731_;
	assign _1733_ = _1729_ & ~_1732_;
	assign _1734_ = _1728_ & ~_1733_;
	assign _1735_ = _1731_ ^ _1730_;
	assign _1736_ = _1729_ & ~_1735_;
	assign _1737_ = _0314_ & ~io_in[13];
	assign _1738_ = _0151_ & ~io_in[13];
	assign _1739_ = _1737_ | ~_1738_;
	assign _1740_ = _0150_ & ~io_in[13];
	assign _1741_ = _0313_ & ~io_in[13];
	assign _1742_ = _1740_ & ~_1741_;
	assign _1743_ = _1738_ ^ _1737_;
	assign _1744_ = _1742_ & ~_1743_;
	assign _1745_ = _1739_ & ~_1744_;
	assign _1746_ = _1736_ & ~_1745_;
	assign _1747_ = _1734_ & ~_1746_;
	assign _1748_ = _1741_ ^ _1740_;
	assign _1749_ = _1748_ | _1743_;
	assign _1750_ = _1736_ & ~_1749_;
	assign _1751_ = _0312_ & ~io_in[13];
	assign _1752_ = _0149_ & ~io_in[13];
	assign _1753_ = _1751_ | ~_1752_;
	assign _1754_ = ~(_1752_ ^ _1751_);
	assign _1755_ = _0311_ & ~io_in[13];
	assign _1756_ = _0148_ & ~io_in[13];
	assign _1757_ = _1755_ | ~_1756_;
	assign _1758_ = _1754_ & ~_1757_;
	assign _1759_ = _1753_ & ~_1758_;
	assign _1760_ = _1756_ ^ _1755_;
	assign _1761_ = _1754_ & ~_1760_;
	assign _1762_ = _0310_ & ~io_in[13];
	assign _1763_ = _0147_ & ~io_in[13];
	assign _1764_ = _1762_ | ~_1763_;
	assign _1765_ = _0146_ & ~io_in[13];
	assign _1766_ = _0309_ & ~io_in[13];
	assign _1767_ = _1765_ & ~_1766_;
	assign _1768_ = _1763_ ^ _1762_;
	assign _1769_ = _1767_ & ~_1768_;
	assign _1770_ = _1764_ & ~_1769_;
	assign _1771_ = _1761_ & ~_1770_;
	assign _1772_ = _1759_ & ~_1771_;
	assign _1773_ = _1750_ & ~_1772_;
	assign _1774_ = _1747_ & ~_1773_;
	assign _1775_ = _1766_ ^ _1765_;
	assign _1776_ = ~(_1775_ | _1768_);
	assign _1777_ = ~(_1776_ & _1761_);
	assign _1778_ = _1750_ & ~_1777_;
	assign _1779_ = _0324_ & ~io_in[13];
	assign _1780_ = _0145_ & ~io_in[13];
	assign _1781_ = _1779_ | ~_1780_;
	assign _1782_ = ~(_1780_ ^ _1779_);
	assign _1783_ = _0323_ & ~io_in[13];
	assign _1784_ = _0144_ & ~io_in[13];
	assign _1785_ = _1783_ | ~_1784_;
	assign _1786_ = _1782_ & ~_1785_;
	assign _1787_ = _1781_ & ~_1786_;
	assign _1788_ = _1784_ ^ _1783_;
	assign _1789_ = _1782_ & ~_1788_;
	assign _1790_ = _0322_ & ~io_in[13];
	assign _1791_ = _0143_ & ~io_in[13];
	assign _1792_ = _1790_ | ~_1791_;
	assign _1793_ = _0142_ & ~io_in[13];
	assign _1794_ = _0321_ & ~io_in[13];
	assign _1795_ = _1793_ & ~_1794_;
	assign _1796_ = _1791_ ^ _1790_;
	assign _1797_ = _1795_ & ~_1796_;
	assign _1798_ = _1792_ & ~_1797_;
	assign _1799_ = _1789_ & ~_1798_;
	assign _1800_ = _1787_ & ~_1799_;
	assign _1801_ = _1794_ ^ _1793_;
	assign _1802_ = _1801_ | _1796_;
	assign _1803_ = _1789_ & ~_1802_;
	assign _1804_ = _0320_ & ~io_in[13];
	assign _1805_ = _0141_ & ~io_in[13];
	assign _1806_ = _1804_ | ~_1805_;
	assign _1807_ = ~(_1805_ ^ _1804_);
	assign _1808_ = _0319_ & ~io_in[13];
	assign _1809_ = _0140_ & ~io_in[13];
	assign _1810_ = _1808_ | ~_1809_;
	assign _1811_ = _1807_ & ~_1810_;
	assign _1812_ = _1806_ & ~_1811_;
	assign _1813_ = _1809_ ^ _1808_;
	assign _1814_ = _1807_ & ~_1813_;
	assign _1815_ = _0318_ & ~io_in[13];
	assign _1816_ = _0139_ & ~io_in[13];
	assign _1817_ = _1815_ | ~_1816_;
	assign _1818_ = ~(_1816_ ^ _1815_);
	assign _1819_ = _0317_ & ~io_in[13];
	assign _1820_ = ~(_0138_ | io_in[13]);
	assign _1821_ = _1820_ & _1819_;
	assign _1822_ = _1818_ & ~_1821_;
	assign _1823_ = _1817_ & ~_1822_;
	assign _1824_ = _1814_ & ~_1823_;
	assign _1825_ = _1812_ & ~_1824_;
	assign _1826_ = _1803_ & ~_1825_;
	assign _1827_ = _1800_ & ~_1826_;
	assign _1828_ = _1778_ & ~_1827_;
	assign _1829_ = _1774_ & ~_1828_;
	assign _1830_ = ~(_1523_ | _1519_);
	assign _1831_ = _1512_ | _1508_;
	assign _1832_ = _1830_ & ~_1831_;
	assign _1833_ = _1497_ | _1494_;
	assign _1834_ = _1504_ | _1501_;
	assign _1835_ = _1834_ | _1833_;
	assign _1836_ = _1832_ & ~_1835_;
	assign \mchip.M2.PWM2  = _1829_ & ~_1836_;
	assign _1837_ = _0356_ & ~io_in[13];
	assign _1838_ = _0169_ & ~io_in[13];
	assign _1839_ = _1837_ | ~_1838_;
	assign _1840_ = ~(_1838_ ^ _1837_);
	assign _1841_ = _0355_ & ~io_in[13];
	assign _1842_ = _0168_ & ~io_in[13];
	assign _1843_ = _1841_ | ~_1842_;
	assign _1844_ = _1840_ & ~_1843_;
	assign _1845_ = _1839_ & ~_1844_;
	assign _1846_ = _1842_ ^ _1841_;
	assign _1847_ = _1840_ & ~_1846_;
	assign _1848_ = _0354_ & ~io_in[13];
	assign _1849_ = _0167_ & ~io_in[13];
	assign _1850_ = _1848_ | ~_1849_;
	assign _1851_ = _0166_ & ~io_in[13];
	assign _1852_ = _0353_ & ~io_in[13];
	assign _1853_ = _1851_ & ~_1852_;
	assign _1854_ = _1849_ ^ _1848_;
	assign _1855_ = _1853_ & ~_1854_;
	assign _1856_ = _1850_ & ~_1855_;
	assign _1857_ = _1847_ & ~_1856_;
	assign _1858_ = _1845_ & ~_1857_;
	assign _1859_ = _1852_ ^ _1851_;
	assign _1860_ = _1859_ | _1854_;
	assign _1861_ = _1847_ & ~_1860_;
	assign _1862_ = _0352_ & ~io_in[13];
	assign _1863_ = _0165_ & ~io_in[13];
	assign _1864_ = _1862_ | ~_1863_;
	assign _1865_ = ~(_1863_ ^ _1862_);
	assign _1866_ = _0351_ & ~io_in[13];
	assign _1867_ = _0164_ & ~io_in[13];
	assign _1868_ = _1866_ | ~_1867_;
	assign _1869_ = _1865_ & ~_1868_;
	assign _1870_ = _1864_ & ~_1869_;
	assign _1871_ = _1867_ ^ _1866_;
	assign _1872_ = _1865_ & ~_1871_;
	assign _1873_ = _0350_ & ~io_in[13];
	assign _1874_ = _0163_ & ~io_in[13];
	assign _1875_ = _1873_ | ~_1874_;
	assign _1876_ = _0162_ & ~io_in[13];
	assign _1877_ = _0349_ & ~io_in[13];
	assign _1878_ = _1876_ & ~_1877_;
	assign _1879_ = _1874_ ^ _1873_;
	assign _1880_ = _1878_ & ~_1879_;
	assign _1881_ = _1875_ & ~_1880_;
	assign _1882_ = _1872_ & ~_1881_;
	assign _1883_ = _1870_ & ~_1882_;
	assign _1884_ = _1861_ & ~_1883_;
	assign _1885_ = _1858_ & ~_1884_;
	assign _1886_ = _1877_ ^ _1876_;
	assign _1887_ = ~(_1886_ | _1879_);
	assign _1888_ = ~(_1887_ & _1872_);
	assign _0405_ = _1861_ & ~_1888_;
	assign _0406_ = _0364_ & ~io_in[13];
	assign _0407_ = _0161_ & ~io_in[13];
	assign _0408_ = _0406_ | ~_0407_;
	assign _0409_ = ~(_0407_ ^ _0406_);
	assign _0410_ = _0363_ & ~io_in[13];
	assign _0411_ = _0160_ & ~io_in[13];
	assign _0412_ = _0410_ | ~_0411_;
	assign _0413_ = _0409_ & ~_0412_;
	assign _0414_ = _0408_ & ~_0413_;
	assign _0415_ = _0411_ ^ _0410_;
	assign _0416_ = _0409_ & ~_0415_;
	assign _0417_ = _0362_ & ~io_in[13];
	assign _0418_ = _0159_ & ~io_in[13];
	assign _0419_ = _0417_ | ~_0418_;
	assign _0420_ = _0158_ & ~io_in[13];
	assign _0421_ = _0361_ & ~io_in[13];
	assign _0422_ = _0420_ & ~_0421_;
	assign _0423_ = _0418_ ^ _0417_;
	assign _0424_ = _0422_ & ~_0423_;
	assign _0425_ = _0419_ & ~_0424_;
	assign _0426_ = _0416_ & ~_0425_;
	assign _0427_ = _0414_ & ~_0426_;
	assign _0428_ = _0421_ ^ _0420_;
	assign _0429_ = _0428_ | _0423_;
	assign _0430_ = _0416_ & ~_0429_;
	assign _0431_ = _0360_ & ~io_in[13];
	assign _0432_ = _0157_ & ~io_in[13];
	assign _0433_ = _0431_ | ~_0432_;
	assign _0434_ = ~(_0432_ ^ _0431_);
	assign _0435_ = _0359_ & ~io_in[13];
	assign _0436_ = _0156_ & ~io_in[13];
	assign _0437_ = _0435_ | ~_0436_;
	assign _0438_ = _0434_ & ~_0437_;
	assign _0439_ = _0433_ & ~_0438_;
	assign _0440_ = _0436_ ^ _0435_;
	assign _0441_ = _0434_ & ~_0440_;
	assign _0442_ = _0358_ & ~io_in[13];
	assign _0443_ = _0155_ & ~io_in[13];
	assign _0444_ = _0442_ | ~_0443_;
	assign _0445_ = ~(_0443_ ^ _0442_);
	assign _0446_ = _0357_ & ~io_in[13];
	assign _0447_ = ~(_0154_ | io_in[13]);
	assign _0448_ = _0447_ & _0446_;
	assign _0449_ = _0445_ & ~_0448_;
	assign _0450_ = _0444_ & ~_0449_;
	assign _0451_ = _0441_ & ~_0450_;
	assign _0452_ = _0439_ & ~_0451_;
	assign _0453_ = _0430_ & ~_0452_;
	assign _0454_ = _0427_ & ~_0453_;
	assign _0455_ = _0405_ & ~_0454_;
	assign _0456_ = _1885_ & ~_0455_;
	assign _0457_ = ~(_1453_ | _1449_);
	assign _0458_ = _1444_ | _1440_;
	assign _0459_ = _0457_ & ~_0458_;
	assign _0460_ = _1473_ | _1470_;
	assign _0461_ = _1466_ | _1463_;
	assign _0462_ = _0461_ | _0460_;
	assign _0463_ = _0459_ & ~_0462_;
	assign \mchip.M2.PWM1  = _0456_ & ~_0463_;
	assign _0097_ = _0120_ & ~_1603_;
	assign _0464_ = ~(_1603_ ^ _1602_);
	assign _0098_ = _0120_ & ~_0464_;
	assign _0465_ = ~_1599_;
	assign _0466_ = _1604_ ^ _0465_;
	assign _0099_ = _0120_ & ~_0466_;
	assign _0467_ = ~(_1604_ & _1599_);
	assign _0468_ = _0467_ ^ _1598_;
	assign _0100_ = _0120_ & ~_0468_;
	assign _0469_ = ~_1595_;
	assign _0470_ = ~(_1599_ & _1598_);
	assign _0471_ = _1604_ & ~_0470_;
	assign _0472_ = _0471_ ^ _0469_;
	assign _0101_ = _0120_ & ~_0472_;
	assign _0473_ = _0471_ & ~_0469_;
	assign _0474_ = _0473_ ^ _1596_;
	assign _0102_ = _0120_ & ~_0474_;
	assign _0103_ = _1662_ & _1619_;
	assign io_out[4] = _0365_ & ~io_in[13];
	assign _0109_ = (_1662_ ? _1618_ : io_out[4]);
	assign io_out[5] = _0366_ & ~io_in[13];
	assign _0110_ = (_1662_ ? _1622_ : io_out[5]);
	assign io_out[6] = _0367_ & ~io_in[13];
	assign _0111_ = (_1662_ ? _1621_ : io_out[6]);
	assign io_out[7] = _0368_ & ~io_in[13];
	assign _0112_ = (_1662_ ? _1626_ : io_out[7]);
	assign io_out[8] = _0369_ & ~io_in[13];
	assign _0113_ = (_1662_ ? _1625_ : io_out[8]);
	assign io_out[9] = _0370_ & ~io_in[13];
	assign _0114_ = (_1662_ ? _1629_ : io_out[9]);
	assign io_out[10] = _0371_ & ~io_in[13];
	assign _0115_ = (_1662_ ? _1628_ : io_out[10]);
	assign io_out[11] = _0372_ & ~io_in[13];
	assign _0116_ = (_1662_ ? _1634_ : io_out[11]);
	assign _0117_ = _1633_ | ~_1662_;
	assign _0104_ = _1637_ | ~_1662_;
	assign _0105_ = _1636_ | ~_1662_;
	assign _0106_ = _1642_ | ~_1662_;
	assign _0107_ = _1641_ | ~_1662_;
	assign _0108_ = _1645_ | ~_1662_;
	assign _0073_ = ~(_0119_ & _1522_);
	assign _0475_ = ~(_1522_ ^ _1520_);
	assign _0074_ = _0119_ & ~_0475_;
	assign _0476_ = ~_1513_;
	assign _0477_ = _1522_ & _1520_;
	assign _0478_ = _0477_ ^ _0476_;
	assign _0075_ = _0119_ & ~_0478_;
	assign _0479_ = ~(_0477_ & _1513_);
	assign _0480_ = _0479_ ^ _1509_;
	assign _0076_ = _0119_ & ~_0480_;
	assign _0481_ = ~_1500_;
	assign _0482_ = ~(_1513_ & _1509_);
	assign _0483_ = _0477_ & ~_0482_;
	assign _0484_ = _0483_ ^ _0481_;
	assign _0077_ = _0119_ & ~_0484_;
	assign _0485_ = ~(_0483_ & _1500_);
	assign _0486_ = _0485_ ^ _1503_;
	assign _0078_ = _0119_ & ~_0486_;
	assign _0487_ = ~(_1503_ & _1500_);
	assign _0488_ = _0483_ & ~_0487_;
	assign _0489_ = ~(_0488_ ^ _1496_);
	assign _0079_ = _0119_ & ~_0489_;
	assign _0490_ = ~(_0488_ & _1496_);
	assign _0491_ = _0490_ ^ _1493_;
	assign _0080_ = _0119_ & ~_0491_;
	assign _0492_ = io_in[13] | ~_0308_;
	assign _0493_ = _0307_ & ~io_in[13];
	assign _0494_ = _0492_ & ~_0493_;
	assign _0495_ = _0306_ & ~io_in[13];
	assign _0496_ = _0305_ & ~io_in[13];
	assign _0497_ = _0496_ | _0495_;
	assign _0498_ = _0494_ & ~_0497_;
	assign _0499_ = io_in[13] | ~_0304_;
	assign _0500_ = _0303_ & ~io_in[13];
	assign _0501_ = _0499_ & ~_0500_;
	assign _0502_ = _0301_ & ~io_in[13];
	assign _0503_ = _0302_ & ~io_in[13];
	assign _0504_ = _0503_ | _0502_;
	assign _0505_ = _0501_ & ~_0504_;
	assign _0506_ = _0498_ & ~_0505_;
	assign _0507_ = _0498_ & ~_0506_;
	assign _0508_ = _0293_ & ~io_in[13];
	assign _0509_ = _0508_ ^ _0507_;
	assign _0510_ = _0509_ ^ _1765_;
	assign _0511_ = ~_1763_;
	assign _0512_ = _0507_ & ~_0508_;
	assign _0513_ = _0294_ & ~io_in[13];
	assign _0514_ = _0513_ ^ _0512_;
	assign _0515_ = _0514_ ^ _0511_;
	assign _0516_ = _0515_ & ~_0510_;
	assign _0517_ = ~_1752_;
	assign _0518_ = _0506_ | ~_0498_;
	assign _0519_ = _0513_ | _0508_;
	assign _0520_ = _0519_ | _0518_;
	assign _0521_ = _0295_ & ~io_in[13];
	assign _0522_ = _0521_ | _0520_;
	assign _0523_ = _0296_ & ~io_in[13];
	assign _0524_ = ~(_0523_ ^ _0522_);
	assign _0525_ = _0524_ ^ _0517_;
	assign _0526_ = ~_1756_;
	assign _0527_ = _0521_ ^ _0520_;
	assign _0528_ = _0527_ ^ _0526_;
	assign _0529_ = _0528_ | ~_0525_;
	assign _0530_ = _0516_ & ~_0529_;
	assign _0531_ = ~_1727_;
	assign _0532_ = _0298_ & ~io_in[13];
	assign _0533_ = _0297_ & ~io_in[13];
	assign _0534_ = ~(_0533_ | _0532_);
	assign _0535_ = _0523_ | _0521_;
	assign _0536_ = _0535_ | _0519_;
	assign _0537_ = _0518_ & ~_0536_;
	assign _0538_ = _0537_ | _0536_;
	assign _0539_ = _0538_ | ~_0534_;
	assign _0540_ = _0299_ & ~io_in[13];
	assign _0541_ = _0540_ | _0539_;
	assign _0542_ = _0300_ & ~io_in[13];
	assign _0543_ = ~_0542_;
	assign _0544_ = _0543_ ^ _0541_;
	assign _0545_ = _0544_ ^ _0531_;
	assign _0546_ = ~_1731_;
	assign _0547_ = _0540_ ^ _0539_;
	assign _0548_ = _0547_ ^ _0546_;
	assign _0549_ = _0545_ & ~_0548_;
	assign _0550_ = ~_1740_;
	assign _0551_ = _0538_ ^ _0533_;
	assign _0552_ = _0551_ ^ _0550_;
	assign _0553_ = ~_0533_;
	assign _0554_ = _0553_ & ~_0538_;
	assign _0555_ = _0554_ ^ _0532_;
	assign _0556_ = _0555_ ^ _1738_;
	assign _0557_ = _0556_ | _0552_;
	assign _0558_ = _0557_ | ~_0549_;
	assign _0559_ = _0530_ & ~_0558_;
	assign _0560_ = _0505_ ^ _0496_;
	assign _0561_ = _0560_ ^ _1793_;
	assign _0562_ = ~_1791_;
	assign _0563_ = _0505_ & ~_0496_;
	assign _0564_ = _0563_ ^ _0495_;
	assign _0565_ = _0564_ ^ _0562_;
	assign _0566_ = _0565_ & ~_0561_;
	assign _0567_ = ~_1780_;
	assign _0568_ = _0505_ & ~_0497_;
	assign _0569_ = _0568_ & ~_0493_;
	assign _0570_ = ~(_0569_ ^ _0492_);
	assign _0571_ = _0570_ ^ _0567_;
	assign _0572_ = ~_1784_;
	assign _0573_ = ~_0493_;
	assign _0574_ = _0568_ ^ _0573_;
	assign _0575_ = _0574_ ^ _0572_;
	assign _0576_ = _0575_ | ~_0571_;
	assign _0577_ = _0566_ & ~_0576_;
	assign _0578_ = ~_1809_;
	assign _0579_ = ~(_0504_ ^ _0500_);
	assign _0580_ = _0579_ ^ _0578_;
	assign _0581_ = _0504_ | _0500_;
	assign _0582_ = _0581_ ^ _0499_;
	assign _0583_ = _0582_ ^ _1805_;
	assign _0584_ = _0580_ & ~_0583_;
	assign _0585_ = ~_1816_;
	assign _0586_ = ~(_0503_ ^ _0502_);
	assign _0587_ = _0586_ ^ _0585_;
	assign _0588_ = ~(_0502_ ^ _1820_);
	assign _0589_ = _0588_ & _0587_;
	assign _0590_ = _0589_ & _0584_;
	assign _0591_ = ~(_0590_ & _0577_);
	assign _0592_ = _0591_ | ~_0559_;
	assign _0593_ = _0570_ | _0567_;
	assign _0594_ = ~(_0574_ & _1784_);
	assign _0595_ = _0571_ & ~_0594_;
	assign _0596_ = _0593_ & ~_0595_;
	assign _0597_ = _0564_ | _0562_;
	assign _0598_ = ~_1793_;
	assign _0599_ = _0560_ | _0598_;
	assign _0600_ = _0565_ & ~_0599_;
	assign _0601_ = _0597_ & ~_0600_;
	assign _0602_ = ~(_0601_ | _0576_);
	assign _0603_ = _0596_ & ~_0602_;
	assign _0604_ = ~_1805_;
	assign _0605_ = _0582_ | _0604_;
	assign _0606_ = _1809_ & ~_0579_;
	assign _0607_ = _0606_ & ~_0583_;
	assign _0608_ = _0605_ & ~_0607_;
	assign _0609_ = _0586_ | _0585_;
	assign _0610_ = _1820_ & ~_0502_;
	assign _0611_ = _0587_ & ~_0610_;
	assign _0612_ = _0609_ & ~_0611_;
	assign _0613_ = _0584_ & ~_0612_;
	assign _0614_ = _0608_ & ~_0613_;
	assign _0615_ = _0577_ & ~_0614_;
	assign _0616_ = _0603_ & ~_0615_;
	assign _0617_ = _0559_ & ~_0616_;
	assign _0618_ = _0524_ | _0517_;
	assign _0619_ = ~(_0527_ & _1756_);
	assign _0620_ = _0525_ & ~_0619_;
	assign _0621_ = _0618_ & ~_0620_;
	assign _0622_ = _0514_ | _0511_;
	assign _0623_ = ~_1765_;
	assign _0624_ = _0509_ | _0623_;
	assign _0625_ = _0515_ & ~_0624_;
	assign _0626_ = _0622_ & ~_0625_;
	assign _0627_ = ~(_0626_ | _0529_);
	assign _0628_ = _0621_ & ~_0627_;
	assign _0629_ = ~(_0628_ | _0558_);
	assign _0630_ = ~_1738_;
	assign _0631_ = _0555_ | _0630_;
	assign _0632_ = _0551_ & ~_0550_;
	assign _0633_ = _0632_ & ~_0556_;
	assign _0634_ = _0631_ & ~_0633_;
	assign _0635_ = _0549_ & ~_0634_;
	assign _0636_ = ~(_0547_ & _1731_);
	assign _0637_ = _0545_ & ~_0636_;
	assign _0638_ = _1727_ & ~_0544_;
	assign _0639_ = _0638_ | _0637_;
	assign _0640_ = _0639_ | _0635_;
	assign _0641_ = _0640_ | _0629_;
	assign _0642_ = _0641_ | _0617_;
	assign _0643_ = _0592_ & ~_0642_;
	assign _0081_ = _0643_ & _1820_;
	assign _0644_ = _1820_ ^ _1816_;
	assign _0088_ = _0643_ & ~_0644_;
	assign _0645_ = _1816_ & ~_1820_;
	assign _0646_ = _0645_ ^ _0578_;
	assign _0089_ = _0643_ & ~_0646_;
	assign _0647_ = _0645_ & ~_0578_;
	assign _0648_ = _0647_ ^ _0604_;
	assign _0090_ = _0643_ & ~_0648_;
	assign _0649_ = ~(_1809_ & _1805_);
	assign _0650_ = _0645_ & ~_0649_;
	assign _0651_ = _0650_ ^ _0598_;
	assign _0091_ = _0643_ & ~_0651_;
	assign _0652_ = _0650_ & ~_0598_;
	assign _0653_ = _0652_ ^ _0562_;
	assign _0092_ = _0643_ & ~_0653_;
	assign _0654_ = ~(_1793_ & _1791_);
	assign _0655_ = _0650_ & ~_0654_;
	assign _0656_ = _0655_ ^ _0572_;
	assign _0093_ = _0643_ & ~_0656_;
	assign _0657_ = _0655_ & ~_0572_;
	assign _0658_ = _0657_ ^ _0567_;
	assign _0094_ = _0643_ & ~_0658_;
	assign _0659_ = ~(_1784_ & _1780_);
	assign _0660_ = _0659_ | _0654_;
	assign _0661_ = _0650_ & ~_0660_;
	assign _0662_ = _0661_ ^ _0623_;
	assign _0095_ = _0643_ & ~_0662_;
	assign _0663_ = _0661_ & ~_0623_;
	assign _0664_ = _0663_ ^ _0511_;
	assign _0096_ = _0643_ & ~_0664_;
	assign _0665_ = ~(_1765_ & _1763_);
	assign _0666_ = _0661_ & ~_0665_;
	assign _0667_ = _0666_ ^ _0526_;
	assign _0082_ = _0643_ & ~_0667_;
	assign _0668_ = _0666_ & ~_0526_;
	assign _0669_ = _0668_ ^ _0517_;
	assign _0083_ = _0643_ & ~_0669_;
	assign _0670_ = ~(_1756_ & _1752_);
	assign _0671_ = _0670_ | _0665_;
	assign _0672_ = _0661_ & ~_0671_;
	assign _0673_ = _0672_ ^ _0550_;
	assign _0084_ = _0643_ & ~_0673_;
	assign _0674_ = _0672_ & ~_0550_;
	assign _0675_ = _0674_ ^ _0630_;
	assign _0085_ = _0643_ & ~_0675_;
	assign _0676_ = ~(_1740_ & _1738_);
	assign _0677_ = _0672_ & ~_0676_;
	assign _0678_ = _0677_ ^ _0546_;
	assign _0086_ = _0643_ & ~_0678_;
	assign _0679_ = _0677_ & ~_0546_;
	assign _0680_ = _0679_ ^ _0531_;
	assign _0087_ = _0643_ & ~_0680_;
	assign _0049_ = ~(_0118_ & _1452_);
	assign _0681_ = ~(_1452_ ^ _1450_);
	assign _0050_ = _0118_ & ~_0681_;
	assign _0682_ = ~_1445_;
	assign _0683_ = _1452_ & _1450_;
	assign _0684_ = _0683_ ^ _0682_;
	assign _0051_ = _0118_ & ~_0684_;
	assign _0685_ = ~(_0683_ & _1445_);
	assign _0686_ = _0685_ ^ _1441_;
	assign _0052_ = _0118_ & ~_0686_;
	assign _0687_ = ~_1462_;
	assign _0688_ = ~(_1445_ & _1441_);
	assign _0689_ = _0683_ & ~_0688_;
	assign _0690_ = _0689_ ^ _0687_;
	assign _0053_ = _0118_ & ~_0690_;
	assign _0691_ = ~(_0689_ & _1462_);
	assign _0692_ = _0691_ ^ _1465_;
	assign _0054_ = _0118_ & ~_0692_;
	assign _0693_ = ~(_1465_ & _1462_);
	assign _0694_ = _0689_ & ~_0693_;
	assign _0695_ = ~(_0694_ ^ _1472_);
	assign _0055_ = _0118_ & ~_0695_;
	assign _0696_ = ~(_0694_ & _1472_);
	assign _0697_ = _0696_ ^ _1469_;
	assign _0056_ = _0118_ & ~_0697_;
	assign _0698_ = io_in[13] | ~_0341_;
	assign _0699_ = ~(_0698_ ^ _0447_);
	assign _0700_ = _0342_ & ~io_in[13];
	assign _0701_ = _0700_ ^ _0698_;
	assign _0702_ = _0701_ ^ _0443_;
	assign _0703_ = _0702_ | _0699_;
	assign _0704_ = ~_0432_;
	assign _0705_ = _0698_ & ~_0700_;
	assign _0706_ = _0343_ & ~io_in[13];
	assign _0707_ = _0705_ & ~_0706_;
	assign _0708_ = _0344_ & ~io_in[13];
	assign _0709_ = _0708_ ^ _0707_;
	assign _0710_ = _0709_ ^ _0704_;
	assign _0711_ = _0706_ ^ _0705_;
	assign _0712_ = _0711_ ^ _0436_;
	assign _0713_ = _0712_ | ~_0710_;
	assign _0714_ = _0713_ | _0703_;
	assign _0715_ = ~_0407_;
	assign _0716_ = _0346_ & ~io_in[13];
	assign _0717_ = _0345_ & ~io_in[13];
	assign _0718_ = _0717_ | _0716_;
	assign _0719_ = _0708_ | _0706_;
	assign _0720_ = _0719_ | ~_0705_;
	assign _0721_ = _0720_ | _0718_;
	assign _0722_ = _0347_ & ~io_in[13];
	assign _0723_ = _0722_ | _0721_;
	assign _0724_ = _0348_ & ~io_in[13];
	assign _0725_ = ~_0724_;
	assign _0726_ = _0725_ ^ _0723_;
	assign _0727_ = _0726_ ^ _0715_;
	assign _0728_ = ~_0411_;
	assign _0729_ = _0722_ ^ _0721_;
	assign _0730_ = _0729_ ^ _0728_;
	assign _0731_ = _0727_ & ~_0730_;
	assign _0732_ = ~_0420_;
	assign _0733_ = ~_0717_;
	assign _0734_ = _0720_ ^ _0733_;
	assign _0735_ = _0734_ ^ _0732_;
	assign _0736_ = ~_0418_;
	assign _0737_ = _0733_ & ~_0720_;
	assign _0738_ = _0737_ ^ _0716_;
	assign _0739_ = _0738_ ^ _0736_;
	assign _0740_ = ~(_0739_ & _0735_);
	assign _0741_ = _0740_ | ~_0731_;
	assign _0742_ = _0741_ | _0714_;
	assign _0743_ = ~_1838_;
	assign _0744_ = _0338_ & ~io_in[13];
	assign _0745_ = _0337_ & ~io_in[13];
	assign _0746_ = ~(_0745_ | _0744_);
	assign _0747_ = io_in[13] | ~_0336_;
	assign _0748_ = _0335_ & ~io_in[13];
	assign _0749_ = _0747_ & ~_0748_;
	assign _0750_ = _0334_ & ~io_in[13];
	assign _0751_ = _0333_ & ~io_in[13];
	assign _0752_ = _0751_ | _0750_;
	assign _0753_ = _0752_ | ~_0749_;
	assign _0754_ = _0749_ & ~_0752_;
	assign _0755_ = _0724_ | _0722_;
	assign _0756_ = ~(_0755_ | _0718_);
	assign _0757_ = _0755_ | _0718_;
	assign _0758_ = _0720_ & ~_0757_;
	assign _0759_ = _0756_ & ~_0758_;
	assign _0760_ = _0754_ & ~_0759_;
	assign _0761_ = _0760_ | _0753_;
	assign _0762_ = _0761_ | ~_0746_;
	assign _0763_ = _0339_ & ~io_in[13];
	assign _0764_ = _0763_ | _0762_;
	assign _0765_ = _0340_ & ~io_in[13];
	assign _0766_ = ~_0765_;
	assign _0767_ = _0766_ ^ _0764_;
	assign _0768_ = _0767_ ^ _0743_;
	assign _0769_ = ~_1842_;
	assign _0770_ = _0763_ ^ _0762_;
	assign _0771_ = _0770_ ^ _0769_;
	assign _0772_ = _0768_ & ~_0771_;
	assign _0773_ = ~_1851_;
	assign _0774_ = _0761_ ^ _0745_;
	assign _0775_ = _0774_ ^ _0773_;
	assign _0776_ = ~_0745_;
	assign _0777_ = _0776_ & ~_0761_;
	assign _0778_ = _0777_ ^ _0744_;
	assign _0779_ = _0778_ ^ _1849_;
	assign _0780_ = _0779_ | _0775_;
	assign _0781_ = _0772_ & ~_0780_;
	assign _0782_ = _0759_ ^ _0751_;
	assign _0783_ = _0782_ ^ _1876_;
	assign _0784_ = ~_1874_;
	assign _0785_ = _0759_ & ~_0751_;
	assign _0786_ = _0785_ ^ _0750_;
	assign _0787_ = _0786_ ^ _0784_;
	assign _0788_ = _0787_ & ~_0783_;
	assign _0789_ = ~_1863_;
	assign _0790_ = _0759_ & ~_0752_;
	assign _0791_ = _0790_ & ~_0748_;
	assign _0792_ = ~(_0791_ ^ _0747_);
	assign _0793_ = _0792_ ^ _0789_;
	assign _0794_ = ~_1867_;
	assign _0795_ = ~_0748_;
	assign _0796_ = _0790_ ^ _0795_;
	assign _0797_ = _0796_ ^ _0794_;
	assign _0798_ = _0793_ & ~_0797_;
	assign _0799_ = ~(_0798_ & _0788_);
	assign _0800_ = _0799_ | ~_0781_;
	assign _0801_ = _0800_ | _0742_;
	assign _0802_ = _0726_ | _0715_;
	assign _0803_ = ~(_0729_ & _0411_);
	assign _0804_ = _0727_ & ~_0803_;
	assign _0805_ = _0802_ & ~_0804_;
	assign _0806_ = _0738_ | _0736_;
	assign _0807_ = _0734_ | _0732_;
	assign _0808_ = _0739_ & ~_0807_;
	assign _0809_ = _0806_ & ~_0808_;
	assign _0810_ = _0731_ & ~_0809_;
	assign _0811_ = _0805_ & ~_0810_;
	assign _0812_ = _0709_ | _0704_;
	assign _0813_ = ~_0436_;
	assign _0814_ = _0711_ | _0813_;
	assign _0815_ = _0710_ & ~_0814_;
	assign _0816_ = _0812_ & ~_0815_;
	assign _0817_ = _0701_ | ~_0443_;
	assign _0818_ = ~(_0698_ & _0447_);
	assign _0819_ = _0818_ & ~_0702_;
	assign _0820_ = _0817_ & ~_0819_;
	assign _0821_ = ~(_0820_ | _0713_);
	assign _0822_ = _0816_ & ~_0821_;
	assign _0823_ = ~(_0822_ | _0741_);
	assign _0824_ = _0811_ & ~_0823_;
	assign _0825_ = ~(_0824_ | _0800_);
	assign _0826_ = _0792_ | _0789_;
	assign _0827_ = ~(_0796_ & _1867_);
	assign _0828_ = _0793_ & ~_0827_;
	assign _0829_ = _0826_ & ~_0828_;
	assign _0830_ = _0786_ | _0784_;
	assign _0831_ = ~_1876_;
	assign _0832_ = _0782_ | _0831_;
	assign _0833_ = _0787_ & ~_0832_;
	assign _0834_ = _0830_ & ~_0833_;
	assign _0835_ = _0798_ & ~_0834_;
	assign _0836_ = _0829_ & ~_0835_;
	assign _0837_ = _0781_ & ~_0836_;
	assign _0838_ = ~_1849_;
	assign _0839_ = _0778_ | _0838_;
	assign _0840_ = _0774_ & ~_0773_;
	assign _0841_ = _0840_ & ~_0779_;
	assign _0842_ = _0839_ & ~_0841_;
	assign _0843_ = _0772_ & ~_0842_;
	assign _0844_ = ~(_0770_ & _1842_);
	assign _0845_ = _0768_ & ~_0844_;
	assign _0846_ = _1838_ & ~_0767_;
	assign _0847_ = _0846_ | _0845_;
	assign _0848_ = _0847_ | _0843_;
	assign _0849_ = _0848_ | _0837_;
	assign _0850_ = _0849_ | _0825_;
	assign _0851_ = _0801_ & ~_0850_;
	assign _0057_ = _0851_ & _0447_;
	assign _0852_ = _0447_ ^ _0443_;
	assign _0064_ = _0851_ & ~_0852_;
	assign _0853_ = _0443_ & ~_0447_;
	assign _0854_ = _0853_ ^ _0813_;
	assign _0065_ = _0851_ & ~_0854_;
	assign _0855_ = _0853_ & ~_0813_;
	assign _0856_ = _0855_ ^ _0704_;
	assign _0066_ = _0851_ & ~_0856_;
	assign _0857_ = ~(_0436_ & _0432_);
	assign _0858_ = _0853_ & ~_0857_;
	assign _0859_ = _0858_ ^ _0732_;
	assign _0067_ = _0851_ & ~_0859_;
	assign _0860_ = _0858_ & ~_0732_;
	assign _0861_ = _0860_ ^ _0736_;
	assign _0068_ = _0851_ & ~_0861_;
	assign _0862_ = ~(_0420_ & _0418_);
	assign _0863_ = _0858_ & ~_0862_;
	assign _0864_ = _0863_ ^ _0728_;
	assign _0069_ = _0851_ & ~_0864_;
	assign _0865_ = _0863_ & ~_0728_;
	assign _0866_ = _0865_ ^ _0715_;
	assign _0070_ = _0851_ & ~_0866_;
	assign _0867_ = ~(_0411_ & _0407_);
	assign _0868_ = _0867_ | _0862_;
	assign _0869_ = _0858_ & ~_0868_;
	assign _0870_ = _0869_ ^ _0831_;
	assign _0071_ = _0851_ & ~_0870_;
	assign _0871_ = _0869_ & ~_0831_;
	assign _0872_ = _0871_ ^ _0784_;
	assign _0072_ = _0851_ & ~_0872_;
	assign _0873_ = ~(_1876_ & _1874_);
	assign _0874_ = _0869_ & ~_0873_;
	assign _0875_ = _0874_ ^ _0794_;
	assign _0058_ = _0851_ & ~_0875_;
	assign _0876_ = _0874_ & ~_0794_;
	assign _0877_ = _0876_ ^ _0789_;
	assign _0059_ = _0851_ & ~_0877_;
	assign _0878_ = ~(_1867_ & _1863_);
	assign _0879_ = _0878_ | _0873_;
	assign _0880_ = _0869_ & ~_0879_;
	assign _0881_ = _0880_ ^ _0773_;
	assign _0060_ = _0851_ & ~_0881_;
	assign _0882_ = _0880_ & ~_0773_;
	assign _0883_ = _0882_ ^ _0838_;
	assign _0061_ = _0851_ & ~_0883_;
	assign _0884_ = ~(_1851_ & _1849_);
	assign _0885_ = _0880_ & ~_0884_;
	assign _0886_ = _0885_ ^ _0769_;
	assign _0062_ = _0851_ & ~_0886_;
	assign _0887_ = _0885_ & ~_0769_;
	assign _0888_ = _0887_ ^ _0743_;
	assign _0063_ = _0851_ & ~_0888_;
	assign _0889_ = _1617_ | _1613_;
	assign _0890_ = _1612_ & ~_0889_;
	assign _0891_ = _0890_ & ~_1428_;
	assign _0038_ = (_1610_ ? \mchip.M1.M.read_write  : _0891_);
	assign _0892_ = _1607_ & _1437_;
	assign _0893_ = _0890_ & ~_0892_;
	assign _0039_ = (_1610_ ? \mchip.M1.IN_REG.SHIFT.Q [1] : _0893_);
	assign _0894_ = _1560_ ^ _1432_;
	assign _0895_ = _0890_ & ~_0894_;
	assign _0040_ = (_1610_ ? \mchip.M1.IN_REG.SHIFT.Q [2] : _0895_);
	assign _0896_ = _1560_ | _1614_;
	assign _0897_ = _0896_ ^ _1431_;
	assign _0898_ = _0890_ & ~_0897_;
	assign _0041_ = (_1610_ ? \mchip.M1.IN_REG.SHIFT.Q [3] : _0898_);
	assign _0899_ = ~(_1703_ ^ _1427_);
	assign _0900_ = _0890_ & ~_0899_;
	assign _0042_ = (_1610_ ? \mchip.M1.IN_REG.SHIFT.Q [4] : _0900_);
	assign _0037_ = ~\mchip.M1.S2.EDGE.prev ;
	assign _0901_ = _1414_ | _1410_;
	assign _0902_ = _0901_ | _1417_;
	assign _0903_ = io_out[11] & _1664_;
	assign _0904_ = _0406_ & _1665_;
	assign _0905_ = _1837_ & _1666_;
	assign _0906_ = _0905_ | _0904_;
	assign _0907_ = _0906_ | _0903_;
	assign _0908_ = _1667_ & ~_0725_;
	assign _0909_ = _1669_ & ~_0766_;
	assign _0910_ = _0909_ | _0908_;
	assign _0911_ = _1470_ & ~_1671_;
	assign _0912_ = _1779_ & _1684_;
	assign _0913_ = _0912_ | _0911_;
	assign _0914_ = _0913_ | _0910_;
	assign _0915_ = _0914_ | _0907_;
	assign _0916_ = _1726_ & _1687_;
	assign _0917_ = _1716_ & ~_0492_;
	assign _0918_ = _0917_ | _0916_;
	assign _0919_ = _1714_ & ~_0543_;
	assign _0920_ = _1494_ & ~_1712_;
	assign _0921_ = _0920_ | _0919_;
	assign _0922_ = _0921_ | _0918_;
	assign _0923_ = io_in[13] | ~_0284_;
	assign _0924_ = _1710_ & ~_0923_;
	assign _0925_ = io_in[13] | ~_0276_;
	assign _0926_ = _1708_ & ~_0925_;
	assign _0927_ = _0926_ | _0924_;
	assign _0928_ = io_in[13] | ~_0268_;
	assign _0929_ = _1706_ & ~_0928_;
	assign _0930_ = io_in[13] | ~_0260_;
	assign _0931_ = _1704_ & ~_0930_;
	assign _0932_ = _0931_ | _0929_;
	assign _0933_ = _0932_ | _0927_;
	assign _0934_ = _0933_ | _0922_;
	assign _0935_ = io_in[13] | ~_0252_;
	assign _0936_ = _1700_ & ~_0935_;
	assign _0937_ = io_in[13] | ~_0244_;
	assign _0938_ = _1609_ & ~_0937_;
	assign _0939_ = _0938_ | _0936_;
	assign _0940_ = io_in[13] | ~_0236_;
	assign _0941_ = _1439_ & ~_0940_;
	assign _0942_ = io_in[13] | ~_0228_;
	assign _0943_ = _1562_ & ~_0942_;
	assign _0944_ = _0943_ | _0941_;
	assign _0945_ = _0944_ | _0939_;
	assign _0946_ = io_in[13] | ~_0220_;
	assign _0947_ = _1569_ & ~_0946_;
	assign _0948_ = io_in[13] | ~_0212_;
	assign _0949_ = _1701_ & ~_0948_;
	assign _0950_ = _0949_ | _0947_;
	assign _0951_ = io_in[13] | ~_0204_;
	assign _0952_ = _1719_ & ~_0951_;
	assign _0953_ = io_in[13] | ~_0388_;
	assign _0954_ = _1617_ & ~_0953_;
	assign _0955_ = _0954_ | _0952_;
	assign _0956_ = _0955_ | _0950_;
	assign _0957_ = _0956_ | _0945_;
	assign _0958_ = _0957_ | _0934_;
	assign _0959_ = _0958_ | _0915_;
	assign _0960_ = ~(_1719_ | _1617_);
	assign _0961_ = _1701_ | _1569_;
	assign _0962_ = _0960_ & ~_0961_;
	assign _0963_ = _1700_ | _1609_;
	assign _0964_ = _1562_ | _1439_;
	assign _0965_ = _0964_ | _0963_;
	assign _0966_ = _0962_ & ~_0965_;
	assign _0967_ = _1716_ | _1687_;
	assign _0968_ = _1714_ | ~_1712_;
	assign _0969_ = _0968_ | _0967_;
	assign _0970_ = _1710_ | _1708_;
	assign _0971_ = _1706_ | _1704_;
	assign _0972_ = _0971_ | _0970_;
	assign _0973_ = _0972_ | _0969_;
	assign _0974_ = _0966_ & ~_0973_;
	assign _0975_ = _1666_ | _1665_;
	assign _0976_ = _0975_ | _1664_;
	assign _0977_ = _1669_ | _1667_;
	assign _0978_ = _1684_ | ~_1671_;
	assign _0979_ = _0978_ | _0977_;
	assign _0980_ = _0979_ | _0976_;
	assign _0981_ = _0974_ & ~_0980_;
	assign _0982_ = (_0981_ ? \mchip.M1.MEM.registers[0] [7] : _0959_);
	assign _0983_ = io_out[10] & _1664_;
	assign _0984_ = _0410_ & _1665_;
	assign _0985_ = _1841_ & _1666_;
	assign _0986_ = _0985_ | _0984_;
	assign _0987_ = _0986_ | _0983_;
	assign _0988_ = _0722_ & _1667_;
	assign _0989_ = _0763_ & _1669_;
	assign _0990_ = _0989_ | _0988_;
	assign _0991_ = _1473_ & ~_1671_;
	assign _0992_ = _1783_ & _1684_;
	assign _0993_ = _0992_ | _0991_;
	assign _0994_ = _0993_ | _0990_;
	assign _0995_ = _0994_ | _0987_;
	assign _0996_ = _1730_ & _1687_;
	assign _0997_ = _1716_ & ~_0573_;
	assign _0998_ = _0997_ | _0996_;
	assign _0999_ = _0540_ & _1714_;
	assign _1000_ = _1497_ & ~_1712_;
	assign _1001_ = _1000_ | _0999_;
	assign _1002_ = _1001_ | _0998_;
	assign _1003_ = io_in[13] | ~_0283_;
	assign _1004_ = _1710_ & ~_1003_;
	assign _1005_ = io_in[13] | ~_0275_;
	assign _1006_ = _1708_ & ~_1005_;
	assign _1007_ = _1006_ | _1004_;
	assign _1008_ = io_in[13] | ~_0267_;
	assign _1009_ = _1706_ & ~_1008_;
	assign _1010_ = io_in[13] | ~_0259_;
	assign _1011_ = _1704_ & ~_1010_;
	assign _1012_ = _1011_ | _1009_;
	assign _1013_ = _1012_ | _1007_;
	assign _1014_ = _1013_ | _1002_;
	assign _1015_ = io_in[13] | ~_0251_;
	assign _1016_ = _1700_ & ~_1015_;
	assign _1017_ = io_in[13] | ~_0243_;
	assign _1018_ = _1609_ & ~_1017_;
	assign _1019_ = _1018_ | _1016_;
	assign _1020_ = io_in[13] | ~_0235_;
	assign _1021_ = _1439_ & ~_1020_;
	assign _1022_ = io_in[13] | ~_0227_;
	assign _1023_ = _1562_ & ~_1022_;
	assign _1024_ = _1023_ | _1021_;
	assign _1025_ = _1024_ | _1019_;
	assign _1026_ = io_in[13] | ~_0219_;
	assign _1027_ = _1569_ & ~_1026_;
	assign _1028_ = io_in[13] | ~_0211_;
	assign _1029_ = _1701_ & ~_1028_;
	assign _1030_ = _1029_ | _1027_;
	assign _1031_ = io_in[13] | ~_0203_;
	assign _1032_ = _1719_ & ~_1031_;
	assign _1033_ = io_in[13] | ~_0387_;
	assign _1034_ = _1617_ & ~_1033_;
	assign _1035_ = _1034_ | _1032_;
	assign _1036_ = _1035_ | _1030_;
	assign _1037_ = _1036_ | _1025_;
	assign _1038_ = _1037_ | _1014_;
	assign _1039_ = _1038_ | _0995_;
	assign _1040_ = (_0981_ ? \mchip.M1.MEM.registers[0] [6] : _1039_);
	assign _1041_ = (\mchip.M1.MEM.index [0] ? _1040_ : _0982_);
	assign _1042_ = io_out[9] & _1664_;
	assign _1043_ = _0417_ & _1665_;
	assign _1044_ = _1848_ & _1666_;
	assign _1045_ = _1044_ | _1043_;
	assign _1046_ = _1045_ | _1042_;
	assign _1047_ = _0716_ & _1667_;
	assign _1048_ = _0744_ & _1669_;
	assign _1049_ = _1048_ | _1047_;
	assign _1050_ = _1466_ & ~_1671_;
	assign _1051_ = _1790_ & _1684_;
	assign _1052_ = _1051_ | _1050_;
	assign _1053_ = _1052_ | _1049_;
	assign _1054_ = _1053_ | _1046_;
	assign _1055_ = _1737_ & _1687_;
	assign _1056_ = _0495_ & _1716_;
	assign _1057_ = _1056_ | _1055_;
	assign _1058_ = _0532_ & _1714_;
	assign _1059_ = _1504_ & ~_1712_;
	assign _1060_ = _1059_ | _1058_;
	assign _1061_ = _1060_ | _1057_;
	assign _1062_ = io_in[13] | ~_0282_;
	assign _1063_ = _1710_ & ~_1062_;
	assign _1064_ = io_in[13] | ~_0274_;
	assign _1065_ = _1708_ & ~_1064_;
	assign _1066_ = _1065_ | _1063_;
	assign _1067_ = io_in[13] | ~_0266_;
	assign _1068_ = _1706_ & ~_1067_;
	assign _1069_ = io_in[13] | ~_0258_;
	assign _1070_ = _1704_ & ~_1069_;
	assign _1071_ = _1070_ | _1068_;
	assign _1072_ = _1071_ | _1066_;
	assign _1073_ = _1072_ | _1061_;
	assign _1074_ = io_in[13] | ~_0250_;
	assign _1075_ = _1700_ & ~_1074_;
	assign _1076_ = io_in[13] | ~_0242_;
	assign _1077_ = _1609_ & ~_1076_;
	assign _1078_ = _1077_ | _1075_;
	assign _1079_ = io_in[13] | ~_0234_;
	assign _1080_ = _1439_ & ~_1079_;
	assign _1081_ = io_in[13] | ~_0226_;
	assign _1082_ = _1562_ & ~_1081_;
	assign _1083_ = _1082_ | _1080_;
	assign _1084_ = _1083_ | _1078_;
	assign _1085_ = io_in[13] | ~_0218_;
	assign _1086_ = _1569_ & ~_1085_;
	assign _1087_ = io_in[13] | ~_0210_;
	assign _1088_ = _1701_ & ~_1087_;
	assign _1089_ = _1088_ | _1086_;
	assign _1090_ = io_in[13] | ~_0202_;
	assign _1091_ = _1719_ & ~_1090_;
	assign _1092_ = io_in[13] | ~_0386_;
	assign _1093_ = _1617_ & ~_1092_;
	assign _1094_ = _1093_ | _1091_;
	assign _1095_ = _1094_ | _1089_;
	assign _1096_ = _1095_ | _1084_;
	assign _1097_ = _1096_ | _1073_;
	assign _1098_ = _1097_ | _1054_;
	assign _1099_ = (_0981_ ? \mchip.M1.MEM.registers[0] [5] : _1098_);
	assign _1100_ = io_out[8] & _1664_;
	assign _1101_ = _0421_ & _1665_;
	assign _1102_ = _1852_ & _1666_;
	assign _1103_ = _1102_ | _1101_;
	assign _1104_ = _1103_ | _1100_;
	assign _1105_ = _1667_ & ~_0733_;
	assign _1106_ = _1669_ & ~_0776_;
	assign _1107_ = _1106_ | _1105_;
	assign _1108_ = _1463_ & ~_1671_;
	assign _1109_ = _1794_ & _1684_;
	assign _1110_ = _1109_ | _1108_;
	assign _1111_ = _1110_ | _1107_;
	assign _1112_ = _1111_ | _1104_;
	assign _1113_ = _1741_ & _1687_;
	assign _1114_ = _0496_ & _1716_;
	assign _1115_ = _1114_ | _1113_;
	assign _1116_ = _1714_ & ~_0553_;
	assign _1117_ = _1501_ & ~_1712_;
	assign _1118_ = _1117_ | _1116_;
	assign _1119_ = _1118_ | _1115_;
	assign _1120_ = io_in[13] | ~_0281_;
	assign _1121_ = _1710_ & ~_1120_;
	assign _1122_ = io_in[13] | ~_0273_;
	assign _1123_ = _1708_ & ~_1122_;
	assign _1124_ = _1123_ | _1121_;
	assign _1125_ = io_in[13] | ~_0265_;
	assign _1126_ = _1706_ & ~_1125_;
	assign _1127_ = io_in[13] | ~_0257_;
	assign _1128_ = _1704_ & ~_1127_;
	assign _1129_ = _1128_ | _1126_;
	assign _1130_ = _1129_ | _1124_;
	assign _1131_ = _1130_ | _1119_;
	assign _1132_ = io_in[13] | ~_0249_;
	assign _1133_ = _1700_ & ~_1132_;
	assign _1134_ = io_in[13] | ~_0241_;
	assign _1135_ = _1609_ & ~_1134_;
	assign _1136_ = _1135_ | _1133_;
	assign _1137_ = io_in[13] | ~_0233_;
	assign _1138_ = _1439_ & ~_1137_;
	assign _1139_ = io_in[13] | ~_0225_;
	assign _1140_ = _1562_ & ~_1139_;
	assign _1141_ = _1140_ | _1138_;
	assign _1142_ = _1141_ | _1136_;
	assign _1143_ = io_in[13] | ~_0217_;
	assign _1144_ = _1569_ & ~_1143_;
	assign _1145_ = io_in[13] | ~_0209_;
	assign _1146_ = _1701_ & ~_1145_;
	assign _1147_ = _1146_ | _1144_;
	assign _1148_ = io_in[13] | ~_0201_;
	assign _1149_ = _1719_ & ~_1148_;
	assign _1150_ = io_in[13] | ~_0385_;
	assign _1151_ = _1617_ & ~_1150_;
	assign _1152_ = _1151_ | _1149_;
	assign _1153_ = _1152_ | _1147_;
	assign _1154_ = _1153_ | _1142_;
	assign _1155_ = _1154_ | _1131_;
	assign _1156_ = _1155_ | _1112_;
	assign _1157_ = (_0981_ ? \mchip.M1.MEM.registers[0] [4] : _1156_);
	assign _1158_ = (\mchip.M1.MEM.index [0] ? _1157_ : _1099_);
	assign _1159_ = (\mchip.M1.MEM.index [1] ? _1158_ : _1041_);
	assign _1160_ = io_out[7] & _1664_;
	assign _1161_ = _0431_ & _1665_;
	assign _1162_ = _1862_ & _1666_;
	assign _1163_ = _1162_ | _1161_;
	assign _1164_ = _1163_ | _1160_;
	assign _1165_ = _0708_ & _1667_;
	assign _1166_ = _1669_ & ~_0747_;
	assign _1167_ = _1166_ | _1165_;
	assign _1168_ = _1440_ & ~_1671_;
	assign _1169_ = _1804_ & _1684_;
	assign _1170_ = _1169_ | _1168_;
	assign _1171_ = _1170_ | _1167_;
	assign _1172_ = _1171_ | _1164_;
	assign _1173_ = _1751_ & _1687_;
	assign _1174_ = _1716_ & ~_0499_;
	assign _1175_ = _1174_ | _1173_;
	assign _1176_ = _0523_ & _1714_;
	assign _1177_ = _1508_ & ~_1712_;
	assign _1178_ = _1177_ | _1176_;
	assign _1179_ = _1178_ | _1175_;
	assign _1180_ = io_in[13] | ~_0280_;
	assign _1181_ = _1710_ & ~_1180_;
	assign _1182_ = io_in[13] | ~_0272_;
	assign _1183_ = _1708_ & ~_1182_;
	assign _1184_ = _1183_ | _1181_;
	assign _1185_ = io_in[13] | ~_0264_;
	assign _1186_ = _1706_ & ~_1185_;
	assign _1187_ = io_in[13] | ~_0256_;
	assign _1188_ = _1704_ & ~_1187_;
	assign _1189_ = _1188_ | _1186_;
	assign _1190_ = _1189_ | _1184_;
	assign _1191_ = _1190_ | _1179_;
	assign _1192_ = io_in[13] | ~_0248_;
	assign _1193_ = _1700_ & ~_1192_;
	assign _1194_ = io_in[13] | ~_0240_;
	assign _1195_ = _1609_ & ~_1194_;
	assign _1196_ = _1195_ | _1193_;
	assign _1197_ = io_in[13] | ~_0232_;
	assign _1198_ = _1439_ & ~_1197_;
	assign _1199_ = io_in[13] | ~_0224_;
	assign _1200_ = _1562_ & ~_1199_;
	assign _1201_ = _1200_ | _1198_;
	assign _1202_ = _1201_ | _1196_;
	assign _1203_ = io_in[13] | ~_0216_;
	assign _1204_ = _1569_ & ~_1203_;
	assign _1205_ = io_in[13] | ~_0208_;
	assign _1206_ = _1701_ & ~_1205_;
	assign _1207_ = _1206_ | _1204_;
	assign _1208_ = io_in[13] | ~_0200_;
	assign _1209_ = _1719_ & ~_1208_;
	assign _1210_ = io_in[13] | ~_0384_;
	assign _1211_ = _1617_ & ~_1210_;
	assign _1212_ = _1211_ | _1209_;
	assign _1213_ = _1212_ | _1207_;
	assign _1214_ = _1213_ | _1202_;
	assign _1215_ = _1214_ | _1191_;
	assign _1216_ = _1215_ | _1172_;
	assign _1217_ = (_0981_ ? \mchip.M1.MEM.registers[0] [3] : _1216_);
	assign _1218_ = io_out[6] & _1664_;
	assign _1219_ = _0435_ & _1665_;
	assign _1220_ = _1866_ & _1666_;
	assign _1221_ = _1220_ | _1219_;
	assign _1222_ = _1221_ | _1218_;
	assign _1223_ = _0706_ & _1667_;
	assign _1224_ = _1669_ & ~_0795_;
	assign _1225_ = _1224_ | _1223_;
	assign _1226_ = _1444_ & ~_1671_;
	assign _1227_ = _1808_ & _1684_;
	assign _1228_ = _1227_ | _1226_;
	assign _1229_ = _1228_ | _1225_;
	assign _1230_ = _1229_ | _1222_;
	assign _1231_ = _1755_ & _1687_;
	assign _1232_ = _0500_ & _1716_;
	assign _1233_ = _1232_ | _1231_;
	assign _1234_ = _0521_ & _1714_;
	assign _1235_ = _1512_ & ~_1712_;
	assign _1236_ = _1235_ | _1234_;
	assign _1237_ = _1236_ | _1233_;
	assign _1238_ = io_in[13] | ~_0279_;
	assign _1239_ = _1710_ & ~_1238_;
	assign _1240_ = io_in[13] | ~_0271_;
	assign _1241_ = _1708_ & ~_1240_;
	assign _1242_ = _1241_ | _1239_;
	assign _1243_ = io_in[13] | ~_0263_;
	assign _1244_ = _1706_ & ~_1243_;
	assign _1245_ = io_in[13] | ~_0255_;
	assign _1246_ = _1704_ & ~_1245_;
	assign _1247_ = _1246_ | _1244_;
	assign _1248_ = _1247_ | _1242_;
	assign _1249_ = _1248_ | _1237_;
	assign _1250_ = io_in[13] | ~_0247_;
	assign _1251_ = _1700_ & ~_1250_;
	assign _1252_ = io_in[13] | ~_0239_;
	assign _1253_ = _1609_ & ~_1252_;
	assign _1254_ = _1253_ | _1251_;
	assign _1255_ = io_in[13] | ~_0231_;
	assign _1256_ = _1439_ & ~_1255_;
	assign _1257_ = io_in[13] | ~_0223_;
	assign _1258_ = _1562_ & ~_1257_;
	assign _1259_ = _1258_ | _1256_;
	assign _1260_ = _1259_ | _1254_;
	assign _1261_ = io_in[13] | ~_0215_;
	assign _1262_ = _1569_ & ~_1261_;
	assign _1263_ = io_in[13] | ~_0207_;
	assign _1264_ = _1701_ & ~_1263_;
	assign _1265_ = _1264_ | _1262_;
	assign _1266_ = io_in[13] | ~_0199_;
	assign _1267_ = _1719_ & ~_1266_;
	assign _1268_ = io_in[13] | ~_0383_;
	assign _1269_ = _1617_ & ~_1268_;
	assign _1270_ = _1269_ | _1267_;
	assign _1271_ = _1270_ | _1265_;
	assign _1272_ = _1271_ | _1260_;
	assign _1273_ = _1272_ | _1249_;
	assign _1274_ = _1273_ | _1230_;
	assign _1275_ = (_0981_ ? \mchip.M1.MEM.registers[0] [2] : _1274_);
	assign _1276_ = (\mchip.M1.MEM.index [0] ? _1275_ : _1217_);
	assign _1277_ = io_out[5] & _1664_;
	assign _1278_ = _0442_ & _1665_;
	assign _1279_ = _1873_ & _1666_;
	assign _1280_ = _1279_ | _1278_;
	assign _1281_ = _1280_ | _1277_;
	assign _1282_ = _0700_ & _1667_;
	assign _1283_ = _0750_ & _1669_;
	assign _1284_ = _1283_ | _1282_;
	assign _1285_ = _1449_ & ~_1671_;
	assign _1286_ = _1815_ & _1684_;
	assign _1287_ = _1286_ | _1285_;
	assign _1288_ = _1287_ | _1284_;
	assign _1289_ = _1288_ | _1281_;
	assign _1290_ = _1762_ & _1687_;
	assign _1291_ = _0503_ & _1716_;
	assign _1292_ = _1291_ | _1290_;
	assign _1293_ = _0513_ & _1714_;
	assign _1294_ = _1519_ & ~_1712_;
	assign _1295_ = _1294_ | _1293_;
	assign _1296_ = _1295_ | _1292_;
	assign _1297_ = io_in[13] | ~_0278_;
	assign _1298_ = _1710_ & ~_1297_;
	assign _1299_ = io_in[13] | ~_0270_;
	assign _1300_ = _1708_ & ~_1299_;
	assign _1301_ = _1300_ | _1298_;
	assign _1302_ = io_in[13] | ~_0262_;
	assign _1303_ = _1706_ & ~_1302_;
	assign _1304_ = io_in[13] | ~_0254_;
	assign _1305_ = _1704_ & ~_1304_;
	assign _1306_ = _1305_ | _1303_;
	assign _1307_ = _1306_ | _1301_;
	assign _1308_ = _1307_ | _1296_;
	assign _1309_ = io_in[13] | ~_0246_;
	assign _1310_ = _1700_ & ~_1309_;
	assign _1311_ = io_in[13] | ~_0238_;
	assign _1312_ = _1609_ & ~_1311_;
	assign _1313_ = _1312_ | _1310_;
	assign _1314_ = io_in[13] | ~_0230_;
	assign _1315_ = _1439_ & ~_1314_;
	assign _1316_ = io_in[13] | ~_0222_;
	assign _1317_ = _1562_ & ~_1316_;
	assign _1318_ = _1317_ | _1315_;
	assign _1319_ = _1318_ | _1313_;
	assign _1320_ = io_in[13] | ~_0214_;
	assign _1321_ = _1569_ & ~_1320_;
	assign _1322_ = io_in[13] | ~_0206_;
	assign _1323_ = _1701_ & ~_1322_;
	assign _1324_ = _1323_ | _1321_;
	assign _1325_ = io_in[13] | ~_0198_;
	assign _1326_ = _1719_ & ~_1325_;
	assign _1327_ = io_in[13] | ~_0382_;
	assign _1328_ = _1617_ & ~_1327_;
	assign _1329_ = _1328_ | _1326_;
	assign _1330_ = _1329_ | _1324_;
	assign _1331_ = _1330_ | _1319_;
	assign _1332_ = _1331_ | _1308_;
	assign _1333_ = _1332_ | _1289_;
	assign _1334_ = (_0981_ ? \mchip.M1.MEM.registers[0] [1] : _1333_);
	assign _1335_ = io_out[4] & _1664_;
	assign _1336_ = _0446_ & _1665_;
	assign _1337_ = _1877_ & _1666_;
	assign _1338_ = _1337_ | _1336_;
	assign _1339_ = _1338_ | _1335_;
	assign _1340_ = _1667_ & ~_0698_;
	assign _1341_ = _0751_ & _1669_;
	assign _1342_ = _1341_ | _1340_;
	assign _1343_ = _1453_ & ~_1671_;
	assign _1344_ = _1819_ & _1684_;
	assign _1345_ = _1344_ | _1343_;
	assign _1346_ = _1345_ | _1342_;
	assign _1347_ = _1346_ | _1339_;
	assign _1348_ = _1766_ & _1687_;
	assign _1349_ = _0502_ & _1716_;
	assign _1350_ = _1349_ | _1348_;
	assign _1351_ = _0508_ & _1714_;
	assign _1352_ = _1523_ & ~_1712_;
	assign _1353_ = _1352_ | _1351_;
	assign _1354_ = _1353_ | _1350_;
	assign _1355_ = io_in[13] | ~_0277_;
	assign _1356_ = _1710_ & ~_1355_;
	assign _1357_ = io_in[13] | ~_0269_;
	assign _1358_ = _1708_ & ~_1357_;
	assign _1359_ = _1358_ | _1356_;
	assign _1360_ = io_in[13] | ~_0261_;
	assign _1361_ = _1706_ & ~_1360_;
	assign _1362_ = io_in[13] | ~_0253_;
	assign _1363_ = _1704_ & ~_1362_;
	assign _1364_ = _1363_ | _1361_;
	assign _1365_ = _1364_ | _1359_;
	assign _1366_ = _1365_ | _1354_;
	assign _1367_ = io_in[13] | ~_0245_;
	assign _1368_ = _1700_ & ~_1367_;
	assign _1369_ = io_in[13] | ~_0237_;
	assign _1370_ = _1609_ & ~_1369_;
	assign _1371_ = _1370_ | _1368_;
	assign _1372_ = io_in[13] | ~_0229_;
	assign _1373_ = _1439_ & ~_1372_;
	assign _1374_ = io_in[13] | ~_0221_;
	assign _1375_ = _1562_ & ~_1374_;
	assign _1376_ = _1375_ | _1373_;
	assign _1377_ = _1376_ | _1371_;
	assign _1378_ = io_in[13] | ~_0213_;
	assign _1379_ = _1569_ & ~_1378_;
	assign _1380_ = io_in[13] | ~_0205_;
	assign _1381_ = _1701_ & ~_1380_;
	assign _1382_ = _1381_ | _1379_;
	assign _1383_ = io_in[13] | ~_0197_;
	assign _1384_ = _1719_ & ~_1383_;
	assign _1385_ = io_in[13] | ~_0381_;
	assign _1386_ = _1617_ & ~_1385_;
	assign _1387_ = _1386_ | _1384_;
	assign _1388_ = _1387_ | _1382_;
	assign _1389_ = _1388_ | _1377_;
	assign _1390_ = _1389_ | _1366_;
	assign _1391_ = _1390_ | _1347_;
	assign _1392_ = (_0981_ ? \mchip.M1.MEM.registers[0] [0] : _1391_);
	assign _1393_ = (\mchip.M1.MEM.index [0] ? _1392_ : _1334_);
	assign _1394_ = (\mchip.M1.MEM.index [1] ? _1393_ : _1276_);
	assign _1395_ = (\mchip.M1.MEM.index [2] ? _1394_ : _1159_);
	assign _1396_ = ~(_1395_ | _1675_);
	assign \mchip.SDA_out  = _1396_ | _0902_;
	assign _0047_ = \mchip.M1.S1.EDGE.prev  & \mchip.M1.S2.EDGE.sig_negedge ;
	assign _0048_ = \mchip.M1.S2.EDGE.sig_posedge  & \mchip.M1.S1.EDGE.prev ;
	assign _0044_ = \mchip.M1.S1.m1.Q  & ~\mchip.M1.S1.EDGE.prev ;
	assign _0043_ = \mchip.M1.S1.EDGE.prev  & ~\mchip.M1.S1.m1.Q ;
	assign _0046_ = \mchip.M1.S2.m1.Q  & ~\mchip.M1.S2.EDGE.prev ;
	assign _0045_ = \mchip.M1.S2.EDGE.prev  & ~\mchip.M1.S2.m1.Q ;
	assign _0036_ = _1421_ & \mchip.M1.S1.EDGE.sig_posedge ;
	assign _1397_ = ~(_1546_ | _1406_);
	assign _1398_ = _1397_ & ~_1404_;
	assign _1399_ = _1404_ & ~_1408_;
	assign _1400_ = _1397_ & ~_1399_;
	assign _1401_ = _1400_ | _1398_;
	assign \mchip.M1.IN_REG.SHIFT.en  = \mchip.M1.S1.EDGE.sig_posedge  & ~_1401_;
	assign _0000_ = _1589_ & ~_1692_;
	assign _1890_[1] = \mchip.M1.COUNT.count [1] ^ \mchip.M1.COUNT.count [0];
	assign _1402_ = \mchip.M1.COUNT.count [1] & \mchip.M1.COUNT.count [0];
	assign _1890_[2] = _1402_ ^ \mchip.M1.COUNT.count [2];
	assign _1403_ = ~(_1402_ & \mchip.M1.COUNT.count [2]);
	assign _1890_[3] = _1403_ ^ _1421_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0121_ <= 1'h1;
		else
			_0121_ <= 1'h0;
	always @(posedge io_in[12])
		if (io_in[13])
			_0122_ <= 1'h0;
		else
			_0122_ <= _0002_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0123_ <= 1'h0;
		else
			_0123_ <= _0003_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0124_ <= 1'h0;
		else
			_0124_ <= _0000_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0125_ <= 1'h0;
		else
			_0125_ <= _0004_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0126_ <= 1'h0;
		else
			_0126_ <= _0005_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0127_ <= 1'h0;
		else
			_0127_ <= _0006_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0128_ <= 1'h0;
		else
			_0128_ <= _0007_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0129_ <= 1'h0;
		else
			_0129_ <= _0008_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0130_ <= 1'h0;
		else
			_0130_ <= _0009_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0131_ <= 1'h0;
		else
			_0131_ <= _0001_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0132_ <= 1'h0;
		else
			_0132_ <= _0097_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0133_ <= 1'h0;
		else
			_0133_ <= _0098_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0134_ <= 1'h0;
		else
			_0134_ <= _0099_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0135_ <= 1'h0;
		else
			_0135_ <= _0100_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0136_ <= 1'h0;
		else
			_0136_ <= _0101_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0137_ <= 1'h0;
		else
			_0137_ <= _0102_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0138_ <= 1'h1;
		else if (!_0119_)
			_0138_ <= _0081_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0139_ <= 1'h0;
		else if (!_0119_)
			_0139_ <= _0088_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0140_ <= 1'h0;
		else if (!_0119_)
			_0140_ <= _0089_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0141_ <= 1'h0;
		else if (!_0119_)
			_0141_ <= _0090_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0142_ <= 1'h0;
		else if (!_0119_)
			_0142_ <= _0091_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0143_ <= 1'h0;
		else if (!_0119_)
			_0143_ <= _0092_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0144_ <= 1'h0;
		else if (!_0119_)
			_0144_ <= _0093_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0145_ <= 1'h0;
		else if (!_0119_)
			_0145_ <= _0094_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0146_ <= 1'h0;
		else if (!_0119_)
			_0146_ <= _0095_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0147_ <= 1'h0;
		else if (!_0119_)
			_0147_ <= _0096_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0148_ <= 1'h0;
		else if (!_0119_)
			_0148_ <= _0082_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0149_ <= 1'h0;
		else if (!_0119_)
			_0149_ <= _0083_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0150_ <= 1'h0;
		else if (!_0119_)
			_0150_ <= _0084_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0151_ <= 1'h0;
		else if (!_0119_)
			_0151_ <= _0085_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0152_ <= 1'h0;
		else if (!_0119_)
			_0152_ <= _0086_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0153_ <= 1'h0;
		else if (!_0119_)
			_0153_ <= _0087_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0154_ <= 1'h1;
		else if (!_0118_)
			_0154_ <= _0057_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0155_ <= 1'h0;
		else if (!_0118_)
			_0155_ <= _0064_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0156_ <= 1'h0;
		else if (!_0118_)
			_0156_ <= _0065_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0157_ <= 1'h0;
		else if (!_0118_)
			_0157_ <= _0066_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0158_ <= 1'h0;
		else if (!_0118_)
			_0158_ <= _0067_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0159_ <= 1'h0;
		else if (!_0118_)
			_0159_ <= _0068_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0160_ <= 1'h0;
		else if (!_0118_)
			_0160_ <= _0069_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0161_ <= 1'h0;
		else if (!_0118_)
			_0161_ <= _0070_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0162_ <= 1'h0;
		else if (!_0118_)
			_0162_ <= _0071_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0163_ <= 1'h0;
		else if (!_0118_)
			_0163_ <= _0072_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0164_ <= 1'h0;
		else if (!_0118_)
			_0164_ <= _0058_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0165_ <= 1'h0;
		else if (!_0118_)
			_0165_ <= _0059_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0166_ <= 1'h0;
		else if (!_0118_)
			_0166_ <= _0060_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0167_ <= 1'h0;
		else if (!_0118_)
			_0167_ <= _0061_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0168_ <= 1'h0;
		else if (!_0118_)
			_0168_ <= _0062_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0169_ <= 1'h0;
		else if (!_0118_)
			_0169_ <= _0063_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0170_ <= 1'h0;
		else
			_0170_ <= _0073_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0171_ <= 1'h0;
		else
			_0171_ <= _0074_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0172_ <= 1'h0;
		else
			_0172_ <= _0075_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0173_ <= 1'h0;
		else
			_0173_ <= _0076_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0174_ <= 1'h0;
		else
			_0174_ <= _0077_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0175_ <= 1'h0;
		else
			_0175_ <= _0078_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0176_ <= 1'h0;
		else
			_0176_ <= _0079_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0177_ <= 1'h0;
		else
			_0177_ <= _0080_;
	always @(posedge io_in[12])
		if (\mchip.M1.STOP.clear_stop )
			_0178_ <= 1'h0;
		else if (_0048_)
			_0178_ <= 1'h1;
	always @(posedge io_in[12])
		if (io_in[13])
			_0179_ <= 1'h0;
		else
			_0179_ <= _0049_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0180_ <= 1'h0;
		else
			_0180_ <= _0050_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0181_ <= 1'h0;
		else
			_0181_ <= _0051_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0182_ <= 1'h0;
		else
			_0182_ <= _0052_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0183_ <= 1'h0;
		else
			_0183_ <= _0053_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0184_ <= 1'h0;
		else
			_0184_ <= _0054_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0185_ <= 1'h0;
		else
			_0185_ <= _0055_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0186_ <= 1'h0;
		else
			_0186_ <= _0056_;
	always @(posedge io_in[12]) \mchip.M1.S2.m1.Q  <= io_in[1];
	always @(posedge io_in[12]) \mchip.M1.S1.EDGE.sig_posedge  <= _0044_;
	always @(posedge io_in[12]) \mchip.M1.S1.EDGE.sig_negedge  <= _0043_;
	always @(posedge io_in[12]) \mchip.M1.S1.EDGE.prev  <= \mchip.M1.S1.m1.Q ;
	always @(posedge io_in[12]) \mchip.M1.S2.EDGE.sig_posedge  <= _0046_;
	always @(posedge io_in[12]) \mchip.M1.S2.EDGE.sig_negedge  <= _0045_;
	always @(posedge io_in[12]) \mchip.M1.S2.EDGE.prev  <= \mchip.M1.S2.m1.Q ;
	always @(posedge io_in[12])
		if (io_in[13])
			_0187_ <= 1'h0;
		else if (_0010_)
			_0187_ <= _0038_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0188_ <= 1'h0;
		else if (_0010_)
			_0188_ <= _0039_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0189_ <= 1'h0;
		else if (_0010_)
			_0189_ <= _0040_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0190_ <= 1'h0;
		else if (_0010_)
			_0190_ <= _0041_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0191_ <= 1'h0;
		else if (_0010_)
			_0191_ <= _0042_;
	always @(posedge io_in[12])
		if (\mchip.M1.START.clear_start )
			_0192_ <= 1'h0;
		else if (_0047_)
			_0192_ <= 1'h1;
	always @(posedge io_in[12])
		if (\mchip.M1.COUNT.clear )
			_0193_ <= 1'h0;
		else if (_0036_)
			_0193_ <= _1889_[0];
	always @(posedge io_in[12])
		if (\mchip.M1.COUNT.clear )
			_0194_ <= 1'h0;
		else if (_0036_)
			_0194_ <= _1890_[1];
	always @(posedge io_in[12])
		if (\mchip.M1.COUNT.clear )
			_0195_ <= 1'h0;
		else if (_0036_)
			_0195_ <= _1890_[2];
	always @(posedge io_in[12])
		if (\mchip.M1.COUNT.clear )
			_0196_ <= 1'h0;
		else if (_0036_)
			_0196_ <= _1890_[3];
	always @(posedge io_in[12])
		if (\mchip.M1.S1.EDGE.sig_posedge )
			\mchip.M1.READ_ACK.ACK  <= _0037_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0197_ <= 1'h0;
		else if (_0012_)
			_0197_ <= \mchip.M1.M.read_write ;
	always @(posedge io_in[12])
		if (io_in[13])
			_0198_ <= 1'h0;
		else if (_0012_)
			_0198_ <= \mchip.M1.IN_REG.SHIFT.Q [1];
	always @(posedge io_in[12])
		if (io_in[13])
			_0199_ <= 1'h0;
		else if (_0012_)
			_0199_ <= \mchip.M1.IN_REG.SHIFT.Q [2];
	always @(posedge io_in[12])
		if (io_in[13])
			_0200_ <= 1'h0;
		else if (_0012_)
			_0200_ <= \mchip.M1.IN_REG.SHIFT.Q [3];
	always @(posedge io_in[12])
		if (io_in[13])
			_0201_ <= 1'h0;
		else if (_0012_)
			_0201_ <= \mchip.M1.IN_REG.SHIFT.Q [4];
	always @(posedge io_in[12])
		if (io_in[13])
			_0202_ <= 1'h0;
		else if (_0012_)
			_0202_ <= \mchip.M1.IN_REG.SHIFT.Q [5];
	always @(posedge io_in[12])
		if (io_in[13])
			_0203_ <= 1'h0;
		else if (_0012_)
			_0203_ <= \mchip.M1.IN_REG.SHIFT.Q [6];
	always @(posedge io_in[12])
		if (io_in[13])
			_0204_ <= 1'h0;
		else if (_0012_)
			_0204_ <= \mchip.M1.IN_REG.SHIFT.Q [7];
	always @(posedge io_in[12])
		if (io_in[13])
			_0205_ <= 1'h0;
		else if (_0013_)
			_0205_ <= \mchip.M1.M.read_write ;
	always @(posedge io_in[12])
		if (io_in[13])
			_0206_ <= 1'h0;
		else if (_0013_)
			_0206_ <= \mchip.M1.IN_REG.SHIFT.Q [1];
	always @(posedge io_in[12])
		if (io_in[13])
			_0207_ <= 1'h0;
		else if (_0013_)
			_0207_ <= \mchip.M1.IN_REG.SHIFT.Q [2];
	always @(posedge io_in[12])
		if (io_in[13])
			_0208_ <= 1'h0;
		else if (_0013_)
			_0208_ <= \mchip.M1.IN_REG.SHIFT.Q [3];
	always @(posedge io_in[12])
		if (io_in[13])
			_0209_ <= 1'h0;
		else if (_0013_)
			_0209_ <= \mchip.M1.IN_REG.SHIFT.Q [4];
	always @(posedge io_in[12])
		if (io_in[13])
			_0210_ <= 1'h0;
		else if (_0013_)
			_0210_ <= \mchip.M1.IN_REG.SHIFT.Q [5];
	always @(posedge io_in[12])
		if (io_in[13])
			_0211_ <= 1'h0;
		else if (_0013_)
			_0211_ <= \mchip.M1.IN_REG.SHIFT.Q [6];
	always @(posedge io_in[12])
		if (io_in[13])
			_0212_ <= 1'h0;
		else if (_0013_)
			_0212_ <= \mchip.M1.IN_REG.SHIFT.Q [7];
	always @(posedge io_in[12])
		if (io_in[13])
			_0213_ <= 1'h0;
		else if (_0014_)
			_0213_ <= \mchip.M1.M.read_write ;
	always @(posedge io_in[12])
		if (io_in[13])
			_0214_ <= 1'h0;
		else if (_0014_)
			_0214_ <= \mchip.M1.IN_REG.SHIFT.Q [1];
	always @(posedge io_in[12])
		if (io_in[13])
			_0215_ <= 1'h0;
		else if (_0014_)
			_0215_ <= \mchip.M1.IN_REG.SHIFT.Q [2];
	always @(posedge io_in[12])
		if (io_in[13])
			_0216_ <= 1'h0;
		else if (_0014_)
			_0216_ <= \mchip.M1.IN_REG.SHIFT.Q [3];
	always @(posedge io_in[12])
		if (io_in[13])
			_0217_ <= 1'h0;
		else if (_0014_)
			_0217_ <= \mchip.M1.IN_REG.SHIFT.Q [4];
	always @(posedge io_in[12])
		if (io_in[13])
			_0218_ <= 1'h0;
		else if (_0014_)
			_0218_ <= \mchip.M1.IN_REG.SHIFT.Q [5];
	always @(posedge io_in[12])
		if (io_in[13])
			_0219_ <= 1'h0;
		else if (_0014_)
			_0219_ <= \mchip.M1.IN_REG.SHIFT.Q [6];
	always @(posedge io_in[12])
		if (io_in[13])
			_0220_ <= 1'h0;
		else if (_0014_)
			_0220_ <= \mchip.M1.IN_REG.SHIFT.Q [7];
	always @(posedge io_in[12])
		if (io_in[13])
			_0221_ <= 1'h0;
		else if (_0015_)
			_0221_ <= \mchip.M1.M.read_write ;
	always @(posedge io_in[12])
		if (io_in[13])
			_0222_ <= 1'h0;
		else if (_0015_)
			_0222_ <= \mchip.M1.IN_REG.SHIFT.Q [1];
	always @(posedge io_in[12])
		if (io_in[13])
			_0223_ <= 1'h0;
		else if (_0015_)
			_0223_ <= \mchip.M1.IN_REG.SHIFT.Q [2];
	always @(posedge io_in[12])
		if (io_in[13])
			_0224_ <= 1'h0;
		else if (_0015_)
			_0224_ <= \mchip.M1.IN_REG.SHIFT.Q [3];
	always @(posedge io_in[12])
		if (io_in[13])
			_0225_ <= 1'h0;
		else if (_0015_)
			_0225_ <= \mchip.M1.IN_REG.SHIFT.Q [4];
	always @(posedge io_in[12])
		if (io_in[13])
			_0226_ <= 1'h0;
		else if (_0015_)
			_0226_ <= \mchip.M1.IN_REG.SHIFT.Q [5];
	always @(posedge io_in[12])
		if (io_in[13])
			_0227_ <= 1'h0;
		else if (_0015_)
			_0227_ <= \mchip.M1.IN_REG.SHIFT.Q [6];
	always @(posedge io_in[12])
		if (io_in[13])
			_0228_ <= 1'h0;
		else if (_0015_)
			_0228_ <= \mchip.M1.IN_REG.SHIFT.Q [7];
	always @(posedge io_in[12])
		if (io_in[13])
			_0229_ <= 1'h0;
		else if (_0016_)
			_0229_ <= \mchip.M1.M.read_write ;
	always @(posedge io_in[12])
		if (io_in[13])
			_0230_ <= 1'h0;
		else if (_0016_)
			_0230_ <= \mchip.M1.IN_REG.SHIFT.Q [1];
	always @(posedge io_in[12])
		if (io_in[13])
			_0231_ <= 1'h0;
		else if (_0016_)
			_0231_ <= \mchip.M1.IN_REG.SHIFT.Q [2];
	always @(posedge io_in[12])
		if (io_in[13])
			_0232_ <= 1'h0;
		else if (_0016_)
			_0232_ <= \mchip.M1.IN_REG.SHIFT.Q [3];
	always @(posedge io_in[12])
		if (io_in[13])
			_0233_ <= 1'h0;
		else if (_0016_)
			_0233_ <= \mchip.M1.IN_REG.SHIFT.Q [4];
	always @(posedge io_in[12])
		if (io_in[13])
			_0234_ <= 1'h0;
		else if (_0016_)
			_0234_ <= \mchip.M1.IN_REG.SHIFT.Q [5];
	always @(posedge io_in[12])
		if (io_in[13])
			_0235_ <= 1'h0;
		else if (_0016_)
			_0235_ <= \mchip.M1.IN_REG.SHIFT.Q [6];
	always @(posedge io_in[12])
		if (io_in[13])
			_0236_ <= 1'h0;
		else if (_0016_)
			_0236_ <= \mchip.M1.IN_REG.SHIFT.Q [7];
	always @(posedge io_in[12])
		if (io_in[13])
			_0237_ <= 1'h0;
		else if (_0017_)
			_0237_ <= \mchip.M1.M.read_write ;
	always @(posedge io_in[12])
		if (io_in[13])
			_0238_ <= 1'h0;
		else if (_0017_)
			_0238_ <= \mchip.M1.IN_REG.SHIFT.Q [1];
	always @(posedge io_in[12])
		if (io_in[13])
			_0239_ <= 1'h0;
		else if (_0017_)
			_0239_ <= \mchip.M1.IN_REG.SHIFT.Q [2];
	always @(posedge io_in[12])
		if (io_in[13])
			_0240_ <= 1'h0;
		else if (_0017_)
			_0240_ <= \mchip.M1.IN_REG.SHIFT.Q [3];
	always @(posedge io_in[12])
		if (io_in[13])
			_0241_ <= 1'h0;
		else if (_0017_)
			_0241_ <= \mchip.M1.IN_REG.SHIFT.Q [4];
	always @(posedge io_in[12])
		if (io_in[13])
			_0242_ <= 1'h0;
		else if (_0017_)
			_0242_ <= \mchip.M1.IN_REG.SHIFT.Q [5];
	always @(posedge io_in[12])
		if (io_in[13])
			_0243_ <= 1'h0;
		else if (_0017_)
			_0243_ <= \mchip.M1.IN_REG.SHIFT.Q [6];
	always @(posedge io_in[12])
		if (io_in[13])
			_0244_ <= 1'h0;
		else if (_0017_)
			_0244_ <= \mchip.M1.IN_REG.SHIFT.Q [7];
	always @(posedge io_in[12])
		if (io_in[13])
			_0245_ <= 1'h0;
		else if (_0018_)
			_0245_ <= \mchip.M1.M.read_write ;
	always @(posedge io_in[12])
		if (io_in[13])
			_0246_ <= 1'h0;
		else if (_0018_)
			_0246_ <= \mchip.M1.IN_REG.SHIFT.Q [1];
	always @(posedge io_in[12])
		if (io_in[13])
			_0247_ <= 1'h0;
		else if (_0018_)
			_0247_ <= \mchip.M1.IN_REG.SHIFT.Q [2];
	always @(posedge io_in[12])
		if (io_in[13])
			_0248_ <= 1'h0;
		else if (_0018_)
			_0248_ <= \mchip.M1.IN_REG.SHIFT.Q [3];
	always @(posedge io_in[12])
		if (io_in[13])
			_0249_ <= 1'h0;
		else if (_0018_)
			_0249_ <= \mchip.M1.IN_REG.SHIFT.Q [4];
	always @(posedge io_in[12])
		if (io_in[13])
			_0250_ <= 1'h0;
		else if (_0018_)
			_0250_ <= \mchip.M1.IN_REG.SHIFT.Q [5];
	always @(posedge io_in[12])
		if (io_in[13])
			_0251_ <= 1'h0;
		else if (_0018_)
			_0251_ <= \mchip.M1.IN_REG.SHIFT.Q [6];
	always @(posedge io_in[12])
		if (io_in[13])
			_0252_ <= 1'h0;
		else if (_0018_)
			_0252_ <= \mchip.M1.IN_REG.SHIFT.Q [7];
	always @(posedge io_in[12])
		if (io_in[13])
			_0253_ <= 1'h0;
		else if (_0019_)
			_0253_ <= \mchip.M1.M.read_write ;
	always @(posedge io_in[12])
		if (io_in[13])
			_0254_ <= 1'h0;
		else if (_0019_)
			_0254_ <= \mchip.M1.IN_REG.SHIFT.Q [1];
	always @(posedge io_in[12])
		if (io_in[13])
			_0255_ <= 1'h0;
		else if (_0019_)
			_0255_ <= \mchip.M1.IN_REG.SHIFT.Q [2];
	always @(posedge io_in[12])
		if (io_in[13])
			_0256_ <= 1'h0;
		else if (_0019_)
			_0256_ <= \mchip.M1.IN_REG.SHIFT.Q [3];
	always @(posedge io_in[12])
		if (io_in[13])
			_0257_ <= 1'h0;
		else if (_0019_)
			_0257_ <= \mchip.M1.IN_REG.SHIFT.Q [4];
	always @(posedge io_in[12])
		if (io_in[13])
			_0258_ <= 1'h0;
		else if (_0019_)
			_0258_ <= \mchip.M1.IN_REG.SHIFT.Q [5];
	always @(posedge io_in[12])
		if (io_in[13])
			_0259_ <= 1'h0;
		else if (_0019_)
			_0259_ <= \mchip.M1.IN_REG.SHIFT.Q [6];
	always @(posedge io_in[12])
		if (io_in[13])
			_0260_ <= 1'h0;
		else if (_0019_)
			_0260_ <= \mchip.M1.IN_REG.SHIFT.Q [7];
	always @(posedge io_in[12])
		if (io_in[13])
			_0261_ <= 1'h0;
		else if (_0020_)
			_0261_ <= \mchip.M1.M.read_write ;
	always @(posedge io_in[12])
		if (io_in[13])
			_0262_ <= 1'h0;
		else if (_0020_)
			_0262_ <= \mchip.M1.IN_REG.SHIFT.Q [1];
	always @(posedge io_in[12])
		if (io_in[13])
			_0263_ <= 1'h0;
		else if (_0020_)
			_0263_ <= \mchip.M1.IN_REG.SHIFT.Q [2];
	always @(posedge io_in[12])
		if (io_in[13])
			_0264_ <= 1'h0;
		else if (_0020_)
			_0264_ <= \mchip.M1.IN_REG.SHIFT.Q [3];
	always @(posedge io_in[12])
		if (io_in[13])
			_0265_ <= 1'h0;
		else if (_0020_)
			_0265_ <= \mchip.M1.IN_REG.SHIFT.Q [4];
	always @(posedge io_in[12])
		if (io_in[13])
			_0266_ <= 1'h0;
		else if (_0020_)
			_0266_ <= \mchip.M1.IN_REG.SHIFT.Q [5];
	always @(posedge io_in[12])
		if (io_in[13])
			_0267_ <= 1'h0;
		else if (_0020_)
			_0267_ <= \mchip.M1.IN_REG.SHIFT.Q [6];
	always @(posedge io_in[12])
		if (io_in[13])
			_0268_ <= 1'h0;
		else if (_0020_)
			_0268_ <= \mchip.M1.IN_REG.SHIFT.Q [7];
	always @(posedge io_in[12])
		if (io_in[13])
			_0269_ <= 1'h0;
		else if (_0021_)
			_0269_ <= \mchip.M1.M.read_write ;
	always @(posedge io_in[12])
		if (io_in[13])
			_0270_ <= 1'h0;
		else if (_0021_)
			_0270_ <= \mchip.M1.IN_REG.SHIFT.Q [1];
	always @(posedge io_in[12])
		if (io_in[13])
			_0271_ <= 1'h0;
		else if (_0021_)
			_0271_ <= \mchip.M1.IN_REG.SHIFT.Q [2];
	always @(posedge io_in[12])
		if (io_in[13])
			_0272_ <= 1'h0;
		else if (_0021_)
			_0272_ <= \mchip.M1.IN_REG.SHIFT.Q [3];
	always @(posedge io_in[12])
		if (io_in[13])
			_0273_ <= 1'h0;
		else if (_0021_)
			_0273_ <= \mchip.M1.IN_REG.SHIFT.Q [4];
	always @(posedge io_in[12])
		if (io_in[13])
			_0274_ <= 1'h0;
		else if (_0021_)
			_0274_ <= \mchip.M1.IN_REG.SHIFT.Q [5];
	always @(posedge io_in[12])
		if (io_in[13])
			_0275_ <= 1'h0;
		else if (_0021_)
			_0275_ <= \mchip.M1.IN_REG.SHIFT.Q [6];
	always @(posedge io_in[12])
		if (io_in[13])
			_0276_ <= 1'h0;
		else if (_0021_)
			_0276_ <= \mchip.M1.IN_REG.SHIFT.Q [7];
	always @(posedge io_in[12])
		if (io_in[13])
			_0277_ <= 1'h0;
		else if (_0022_)
			_0277_ <= \mchip.M1.M.read_write ;
	always @(posedge io_in[12])
		if (io_in[13])
			_0278_ <= 1'h0;
		else if (_0022_)
			_0278_ <= \mchip.M1.IN_REG.SHIFT.Q [1];
	always @(posedge io_in[12])
		if (io_in[13])
			_0279_ <= 1'h0;
		else if (_0022_)
			_0279_ <= \mchip.M1.IN_REG.SHIFT.Q [2];
	always @(posedge io_in[12])
		if (io_in[13])
			_0280_ <= 1'h0;
		else if (_0022_)
			_0280_ <= \mchip.M1.IN_REG.SHIFT.Q [3];
	always @(posedge io_in[12])
		if (io_in[13])
			_0281_ <= 1'h0;
		else if (_0022_)
			_0281_ <= \mchip.M1.IN_REG.SHIFT.Q [4];
	always @(posedge io_in[12])
		if (io_in[13])
			_0282_ <= 1'h0;
		else if (_0022_)
			_0282_ <= \mchip.M1.IN_REG.SHIFT.Q [5];
	always @(posedge io_in[12])
		if (io_in[13])
			_0283_ <= 1'h0;
		else if (_0022_)
			_0283_ <= \mchip.M1.IN_REG.SHIFT.Q [6];
	always @(posedge io_in[12])
		if (io_in[13])
			_0284_ <= 1'h0;
		else if (_0022_)
			_0284_ <= \mchip.M1.IN_REG.SHIFT.Q [7];
	always @(posedge io_in[12])
		if (io_in[13])
			_0285_ <= 1'h0;
		else if (_0023_)
			_0285_ <= \mchip.M1.M.read_write ;
	always @(posedge io_in[12])
		if (io_in[13])
			_0286_ <= 1'h0;
		else if (_0023_)
			_0286_ <= \mchip.M1.IN_REG.SHIFT.Q [1];
	always @(posedge io_in[12])
		if (io_in[13])
			_0287_ <= 1'h0;
		else if (_0023_)
			_0287_ <= \mchip.M1.IN_REG.SHIFT.Q [2];
	always @(posedge io_in[12])
		if (io_in[13])
			_0288_ <= 1'h0;
		else if (_0023_)
			_0288_ <= \mchip.M1.IN_REG.SHIFT.Q [3];
	always @(posedge io_in[12])
		if (io_in[13])
			_0289_ <= 1'h0;
		else if (_0023_)
			_0289_ <= \mchip.M1.IN_REG.SHIFT.Q [4];
	always @(posedge io_in[12])
		if (io_in[13])
			_0290_ <= 1'h0;
		else if (_0023_)
			_0290_ <= \mchip.M1.IN_REG.SHIFT.Q [5];
	always @(posedge io_in[12])
		if (io_in[13])
			_0291_ <= 1'h0;
		else if (_0023_)
			_0291_ <= \mchip.M1.IN_REG.SHIFT.Q [6];
	always @(posedge io_in[12])
		if (io_in[13])
			_0292_ <= 1'h0;
		else if (_0023_)
			_0292_ <= \mchip.M1.IN_REG.SHIFT.Q [7];
	always @(posedge io_in[12])
		if (io_in[13])
			_0293_ <= 1'h0;
		else if (_0024_)
			_0293_ <= \mchip.M1.M.read_write ;
	always @(posedge io_in[12])
		if (io_in[13])
			_0294_ <= 1'h0;
		else if (_0024_)
			_0294_ <= \mchip.M1.IN_REG.SHIFT.Q [1];
	always @(posedge io_in[12])
		if (io_in[13])
			_0295_ <= 1'h0;
		else if (_0024_)
			_0295_ <= \mchip.M1.IN_REG.SHIFT.Q [2];
	always @(posedge io_in[12])
		if (io_in[13])
			_0296_ <= 1'h0;
		else if (_0024_)
			_0296_ <= \mchip.M1.IN_REG.SHIFT.Q [3];
	always @(posedge io_in[12])
		if (io_in[13])
			_0297_ <= 1'h0;
		else if (_0024_)
			_0297_ <= \mchip.M1.IN_REG.SHIFT.Q [4];
	always @(posedge io_in[12])
		if (io_in[13])
			_0298_ <= 1'h0;
		else if (_0024_)
			_0298_ <= \mchip.M1.IN_REG.SHIFT.Q [5];
	always @(posedge io_in[12])
		if (io_in[13])
			_0299_ <= 1'h0;
		else if (_0024_)
			_0299_ <= \mchip.M1.IN_REG.SHIFT.Q [6];
	always @(posedge io_in[12])
		if (io_in[13])
			_0300_ <= 1'h0;
		else if (_0024_)
			_0300_ <= \mchip.M1.IN_REG.SHIFT.Q [7];
	always @(posedge io_in[12])
		if (io_in[13])
			_0301_ <= 1'h0;
		else if (_0025_)
			_0301_ <= \mchip.M1.M.read_write ;
	always @(posedge io_in[12])
		if (io_in[13])
			_0302_ <= 1'h0;
		else if (_0025_)
			_0302_ <= \mchip.M1.IN_REG.SHIFT.Q [1];
	always @(posedge io_in[12])
		if (io_in[13])
			_0303_ <= 1'h0;
		else if (_0025_)
			_0303_ <= \mchip.M1.IN_REG.SHIFT.Q [2];
	always @(posedge io_in[12])
		if (io_in[13])
			_0304_ <= 1'h0;
		else if (_0025_)
			_0304_ <= \mchip.M1.IN_REG.SHIFT.Q [3];
	always @(posedge io_in[12])
		if (io_in[13])
			_0305_ <= 1'h0;
		else if (_0025_)
			_0305_ <= \mchip.M1.IN_REG.SHIFT.Q [4];
	always @(posedge io_in[12])
		if (io_in[13])
			_0306_ <= 1'h0;
		else if (_0025_)
			_0306_ <= \mchip.M1.IN_REG.SHIFT.Q [5];
	always @(posedge io_in[12])
		if (io_in[13])
			_0307_ <= 1'h0;
		else if (_0025_)
			_0307_ <= \mchip.M1.IN_REG.SHIFT.Q [6];
	always @(posedge io_in[12])
		if (io_in[13])
			_0308_ <= 1'h0;
		else if (_0025_)
			_0308_ <= \mchip.M1.IN_REG.SHIFT.Q [7];
	always @(posedge io_in[12])
		if (io_in[13])
			_0309_ <= 1'h0;
		else if (_0026_)
			_0309_ <= \mchip.M1.M.read_write ;
	always @(posedge io_in[12])
		if (io_in[13])
			_0310_ <= 1'h0;
		else if (_0026_)
			_0310_ <= \mchip.M1.IN_REG.SHIFT.Q [1];
	always @(posedge io_in[12])
		if (io_in[13])
			_0311_ <= 1'h0;
		else if (_0026_)
			_0311_ <= \mchip.M1.IN_REG.SHIFT.Q [2];
	always @(posedge io_in[12])
		if (io_in[13])
			_0312_ <= 1'h0;
		else if (_0026_)
			_0312_ <= \mchip.M1.IN_REG.SHIFT.Q [3];
	always @(posedge io_in[12])
		if (io_in[13])
			_0313_ <= 1'h0;
		else if (_0026_)
			_0313_ <= \mchip.M1.IN_REG.SHIFT.Q [4];
	always @(posedge io_in[12])
		if (io_in[13])
			_0314_ <= 1'h0;
		else if (_0026_)
			_0314_ <= \mchip.M1.IN_REG.SHIFT.Q [5];
	always @(posedge io_in[12])
		if (io_in[13])
			_0315_ <= 1'h0;
		else if (_0026_)
			_0315_ <= \mchip.M1.IN_REG.SHIFT.Q [6];
	always @(posedge io_in[12])
		if (io_in[13])
			_0316_ <= 1'h0;
		else if (_0026_)
			_0316_ <= \mchip.M1.IN_REG.SHIFT.Q [7];
	always @(posedge io_in[12])
		if (io_in[13])
			_0317_ <= 1'h0;
		else if (_0027_)
			_0317_ <= \mchip.M1.M.read_write ;
	always @(posedge io_in[12])
		if (io_in[13])
			_0318_ <= 1'h0;
		else if (_0027_)
			_0318_ <= \mchip.M1.IN_REG.SHIFT.Q [1];
	always @(posedge io_in[12])
		if (io_in[13])
			_0319_ <= 1'h0;
		else if (_0027_)
			_0319_ <= \mchip.M1.IN_REG.SHIFT.Q [2];
	always @(posedge io_in[12])
		if (io_in[13])
			_0320_ <= 1'h0;
		else if (_0027_)
			_0320_ <= \mchip.M1.IN_REG.SHIFT.Q [3];
	always @(posedge io_in[12])
		if (io_in[13])
			_0321_ <= 1'h0;
		else if (_0027_)
			_0321_ <= \mchip.M1.IN_REG.SHIFT.Q [4];
	always @(posedge io_in[12])
		if (io_in[13])
			_0322_ <= 1'h0;
		else if (_0027_)
			_0322_ <= \mchip.M1.IN_REG.SHIFT.Q [5];
	always @(posedge io_in[12])
		if (io_in[13])
			_0323_ <= 1'h0;
		else if (_0027_)
			_0323_ <= \mchip.M1.IN_REG.SHIFT.Q [6];
	always @(posedge io_in[12])
		if (io_in[13])
			_0324_ <= 1'h0;
		else if (_0027_)
			_0324_ <= \mchip.M1.IN_REG.SHIFT.Q [7];
	always @(posedge io_in[12])
		if (io_in[13])
			_0325_ <= 1'h0;
		else if (_0028_)
			_0325_ <= \mchip.M1.M.read_write ;
	always @(posedge io_in[12])
		if (io_in[13])
			_0326_ <= 1'h0;
		else if (_0028_)
			_0326_ <= \mchip.M1.IN_REG.SHIFT.Q [1];
	always @(posedge io_in[12])
		if (io_in[13])
			_0327_ <= 1'h0;
		else if (_0028_)
			_0327_ <= \mchip.M1.IN_REG.SHIFT.Q [2];
	always @(posedge io_in[12])
		if (io_in[13])
			_0328_ <= 1'h0;
		else if (_0028_)
			_0328_ <= \mchip.M1.IN_REG.SHIFT.Q [3];
	always @(posedge io_in[12])
		if (io_in[13])
			_0329_ <= 1'h0;
		else if (_0028_)
			_0329_ <= \mchip.M1.IN_REG.SHIFT.Q [4];
	always @(posedge io_in[12])
		if (io_in[13])
			_0330_ <= 1'h0;
		else if (_0028_)
			_0330_ <= \mchip.M1.IN_REG.SHIFT.Q [5];
	always @(posedge io_in[12])
		if (io_in[13])
			_0331_ <= 1'h0;
		else if (_0028_)
			_0331_ <= \mchip.M1.IN_REG.SHIFT.Q [6];
	always @(posedge io_in[12])
		if (io_in[13])
			_0332_ <= 1'h0;
		else if (_0028_)
			_0332_ <= \mchip.M1.IN_REG.SHIFT.Q [7];
	always @(posedge io_in[12])
		if (io_in[13])
			_0333_ <= 1'h0;
		else if (_0029_)
			_0333_ <= \mchip.M1.M.read_write ;
	always @(posedge io_in[12])
		if (io_in[13])
			_0334_ <= 1'h0;
		else if (_0029_)
			_0334_ <= \mchip.M1.IN_REG.SHIFT.Q [1];
	always @(posedge io_in[12])
		if (io_in[13])
			_0335_ <= 1'h0;
		else if (_0029_)
			_0335_ <= \mchip.M1.IN_REG.SHIFT.Q [2];
	always @(posedge io_in[12])
		if (io_in[13])
			_0336_ <= 1'h0;
		else if (_0029_)
			_0336_ <= \mchip.M1.IN_REG.SHIFT.Q [3];
	always @(posedge io_in[12])
		if (io_in[13])
			_0337_ <= 1'h0;
		else if (_0029_)
			_0337_ <= \mchip.M1.IN_REG.SHIFT.Q [4];
	always @(posedge io_in[12])
		if (io_in[13])
			_0338_ <= 1'h0;
		else if (_0029_)
			_0338_ <= \mchip.M1.IN_REG.SHIFT.Q [5];
	always @(posedge io_in[12])
		if (io_in[13])
			_0339_ <= 1'h0;
		else if (_0029_)
			_0339_ <= \mchip.M1.IN_REG.SHIFT.Q [6];
	always @(posedge io_in[12])
		if (io_in[13])
			_0340_ <= 1'h0;
		else if (_0029_)
			_0340_ <= \mchip.M1.IN_REG.SHIFT.Q [7];
	always @(posedge io_in[12])
		if (io_in[13])
			_0341_ <= 1'h0;
		else if (_0030_)
			_0341_ <= \mchip.M1.M.read_write ;
	always @(posedge io_in[12])
		if (io_in[13])
			_0342_ <= 1'h0;
		else if (_0030_)
			_0342_ <= \mchip.M1.IN_REG.SHIFT.Q [1];
	always @(posedge io_in[12])
		if (io_in[13])
			_0343_ <= 1'h0;
		else if (_0030_)
			_0343_ <= \mchip.M1.IN_REG.SHIFT.Q [2];
	always @(posedge io_in[12])
		if (io_in[13])
			_0344_ <= 1'h0;
		else if (_0030_)
			_0344_ <= \mchip.M1.IN_REG.SHIFT.Q [3];
	always @(posedge io_in[12])
		if (io_in[13])
			_0345_ <= 1'h0;
		else if (_0030_)
			_0345_ <= \mchip.M1.IN_REG.SHIFT.Q [4];
	always @(posedge io_in[12])
		if (io_in[13])
			_0346_ <= 1'h0;
		else if (_0030_)
			_0346_ <= \mchip.M1.IN_REG.SHIFT.Q [5];
	always @(posedge io_in[12])
		if (io_in[13])
			_0347_ <= 1'h0;
		else if (_0030_)
			_0347_ <= \mchip.M1.IN_REG.SHIFT.Q [6];
	always @(posedge io_in[12])
		if (io_in[13])
			_0348_ <= 1'h0;
		else if (_0030_)
			_0348_ <= \mchip.M1.IN_REG.SHIFT.Q [7];
	always @(posedge io_in[12])
		if (io_in[13])
			_0349_ <= 1'h0;
		else if (_0031_)
			_0349_ <= \mchip.M1.M.read_write ;
	always @(posedge io_in[12])
		if (io_in[13])
			_0350_ <= 1'h0;
		else if (_0031_)
			_0350_ <= \mchip.M1.IN_REG.SHIFT.Q [1];
	always @(posedge io_in[12])
		if (io_in[13])
			_0351_ <= 1'h0;
		else if (_0031_)
			_0351_ <= \mchip.M1.IN_REG.SHIFT.Q [2];
	always @(posedge io_in[12])
		if (io_in[13])
			_0352_ <= 1'h0;
		else if (_0031_)
			_0352_ <= \mchip.M1.IN_REG.SHIFT.Q [3];
	always @(posedge io_in[12])
		if (io_in[13])
			_0353_ <= 1'h0;
		else if (_0031_)
			_0353_ <= \mchip.M1.IN_REG.SHIFT.Q [4];
	always @(posedge io_in[12])
		if (io_in[13])
			_0354_ <= 1'h0;
		else if (_0031_)
			_0354_ <= \mchip.M1.IN_REG.SHIFT.Q [5];
	always @(posedge io_in[12])
		if (io_in[13])
			_0355_ <= 1'h0;
		else if (_0031_)
			_0355_ <= \mchip.M1.IN_REG.SHIFT.Q [6];
	always @(posedge io_in[12])
		if (io_in[13])
			_0356_ <= 1'h0;
		else if (_0031_)
			_0356_ <= \mchip.M1.IN_REG.SHIFT.Q [7];
	always @(posedge io_in[12])
		if (io_in[13])
			_0357_ <= 1'h0;
		else if (_0032_)
			_0357_ <= \mchip.M1.M.read_write ;
	always @(posedge io_in[12])
		if (io_in[13])
			_0358_ <= 1'h0;
		else if (_0032_)
			_0358_ <= \mchip.M1.IN_REG.SHIFT.Q [1];
	always @(posedge io_in[12])
		if (io_in[13])
			_0359_ <= 1'h0;
		else if (_0032_)
			_0359_ <= \mchip.M1.IN_REG.SHIFT.Q [2];
	always @(posedge io_in[12])
		if (io_in[13])
			_0360_ <= 1'h0;
		else if (_0032_)
			_0360_ <= \mchip.M1.IN_REG.SHIFT.Q [3];
	always @(posedge io_in[12])
		if (io_in[13])
			_0361_ <= 1'h0;
		else if (_0032_)
			_0361_ <= \mchip.M1.IN_REG.SHIFT.Q [4];
	always @(posedge io_in[12])
		if (io_in[13])
			_0362_ <= 1'h0;
		else if (_0032_)
			_0362_ <= \mchip.M1.IN_REG.SHIFT.Q [5];
	always @(posedge io_in[12])
		if (io_in[13])
			_0363_ <= 1'h0;
		else if (_0032_)
			_0363_ <= \mchip.M1.IN_REG.SHIFT.Q [6];
	always @(posedge io_in[12])
		if (io_in[13])
			_0364_ <= 1'h0;
		else if (_0032_)
			_0364_ <= \mchip.M1.IN_REG.SHIFT.Q [7];
	always @(posedge io_in[12])
		if (io_in[13])
			_0365_ <= 1'h0;
		else if (_0033_)
			_0365_ <= \mchip.M1.M.read_write ;
	always @(posedge io_in[12])
		if (io_in[13])
			_0366_ <= 1'h0;
		else if (_0033_)
			_0366_ <= \mchip.M1.IN_REG.SHIFT.Q [1];
	always @(posedge io_in[12])
		if (io_in[13])
			_0367_ <= 1'h0;
		else if (_0033_)
			_0367_ <= \mchip.M1.IN_REG.SHIFT.Q [2];
	always @(posedge io_in[12])
		if (io_in[13])
			_0368_ <= 1'h0;
		else if (_0033_)
			_0368_ <= \mchip.M1.IN_REG.SHIFT.Q [3];
	always @(posedge io_in[12])
		if (io_in[13])
			_0369_ <= 1'h0;
		else if (_0033_)
			_0369_ <= \mchip.M1.IN_REG.SHIFT.Q [4];
	always @(posedge io_in[12])
		if (io_in[13])
			_0370_ <= 1'h0;
		else if (_0033_)
			_0370_ <= \mchip.M1.IN_REG.SHIFT.Q [5];
	always @(posedge io_in[12])
		if (io_in[13])
			_0371_ <= 1'h0;
		else if (_0033_)
			_0371_ <= \mchip.M1.IN_REG.SHIFT.Q [6];
	always @(posedge io_in[12])
		if (io_in[13])
			_0372_ <= 1'h0;
		else if (_0033_)
			_0372_ <= \mchip.M1.IN_REG.SHIFT.Q [7];
	always @(posedge io_in[12])
		if (!io_in[13])
			\mchip.M1.MEM.registers[0] [0] <= \mchip.M1.MEM.parallel_in_temp [0];
	always @(posedge io_in[12])
		if (!io_in[13])
			\mchip.M1.MEM.registers[0] [1] <= \mchip.M1.MEM.parallel_in_temp [1];
	always @(posedge io_in[12])
		if (!io_in[13])
			\mchip.M1.MEM.registers[0] [2] <= \mchip.M1.MEM.parallel_in_temp [2];
	always @(posedge io_in[12])
		if (!io_in[13])
			\mchip.M1.MEM.registers[0] [3] <= \mchip.M1.MEM.parallel_in_temp [3];
	always @(posedge io_in[12])
		if (!io_in[13])
			\mchip.M1.MEM.registers[0] [4] <= \mchip.M1.MEM.parallel_in_temp [4];
	always @(posedge io_in[12])
		if (!io_in[13])
			\mchip.M1.MEM.registers[0] [5] <= \mchip.M1.MEM.parallel_in_temp [5];
	always @(posedge io_in[12])
		if (!io_in[13])
			\mchip.M1.MEM.registers[0] [6] <= \mchip.M1.MEM.parallel_in_temp [6];
	always @(posedge io_in[12])
		if (!io_in[13])
			\mchip.M1.MEM.registers[0] [7] <= \mchip.M1.MEM.parallel_in_temp [7];
	always @(posedge io_in[12])
		if (!io_in[13])
			\mchip.M1.MEM.parallel_in_temp [0] <= io_in[4];
	always @(posedge io_in[12])
		if (!io_in[13])
			\mchip.M1.MEM.parallel_in_temp [1] <= io_in[5];
	always @(posedge io_in[12])
		if (!io_in[13])
			\mchip.M1.MEM.parallel_in_temp [2] <= io_in[6];
	always @(posedge io_in[12])
		if (!io_in[13])
			\mchip.M1.MEM.parallel_in_temp [3] <= io_in[7];
	always @(posedge io_in[12])
		if (!io_in[13])
			\mchip.M1.MEM.parallel_in_temp [4] <= io_in[8];
	always @(posedge io_in[12])
		if (!io_in[13])
			\mchip.M1.MEM.parallel_in_temp [5] <= io_in[9];
	always @(posedge io_in[12])
		if (!io_in[13])
			\mchip.M1.MEM.parallel_in_temp [6] <= io_in[10];
	always @(posedge io_in[12])
		if (!io_in[13])
			\mchip.M1.MEM.parallel_in_temp [7] <= io_in[11];
	always @(posedge io_in[12])
		if (_0034_)
			\mchip.M1.MEM.index [0] <= \mchip.M1.COUNT.count [0];
	always @(posedge io_in[12])
		if (_0034_)
			\mchip.M1.MEM.index [1] <= \mchip.M1.COUNT.count [1];
	always @(posedge io_in[12])
		if (_0034_)
			\mchip.M1.MEM.index [2] <= \mchip.M1.COUNT.count [2];
	always @(posedge io_in[12])
		if (io_in[13])
			_0373_ <= 1'h0;
		else if (\mchip.M1.IN_REG.SHIFT.en )
			_0373_ <= \mchip.M1.S2.EDGE.prev ;
	always @(posedge io_in[12])
		if (io_in[13])
			_0374_ <= 1'h0;
		else if (\mchip.M1.IN_REG.SHIFT.en )
			_0374_ <= \mchip.M1.M.read_write ;
	always @(posedge io_in[12])
		if (io_in[13])
			_0375_ <= 1'h0;
		else if (\mchip.M1.IN_REG.SHIFT.en )
			_0375_ <= \mchip.M1.IN_REG.SHIFT.Q [1];
	always @(posedge io_in[12])
		if (io_in[13])
			_0376_ <= 1'h0;
		else if (\mchip.M1.IN_REG.SHIFT.en )
			_0376_ <= \mchip.M1.IN_REG.SHIFT.Q [2];
	always @(posedge io_in[12])
		if (io_in[13])
			_0377_ <= 1'h0;
		else if (\mchip.M1.IN_REG.SHIFT.en )
			_0377_ <= \mchip.M1.IN_REG.SHIFT.Q [3];
	always @(posedge io_in[12])
		if (io_in[13])
			_0378_ <= 1'h0;
		else if (\mchip.M1.IN_REG.SHIFT.en )
			_0378_ <= \mchip.M1.IN_REG.SHIFT.Q [4];
	always @(posedge io_in[12])
		if (io_in[13])
			_0379_ <= 1'h0;
		else if (\mchip.M1.IN_REG.SHIFT.en )
			_0379_ <= \mchip.M1.IN_REG.SHIFT.Q [5];
	always @(posedge io_in[12])
		if (io_in[13])
			_0380_ <= 1'h0;
		else if (\mchip.M1.IN_REG.SHIFT.en )
			_0380_ <= \mchip.M1.IN_REG.SHIFT.Q [6];
	always @(posedge io_in[12])
		if (io_in[13])
			_0381_ <= 1'h0;
		else if (_0011_)
			_0381_ <= \mchip.M1.M.read_write ;
	always @(posedge io_in[12])
		if (io_in[13])
			_0382_ <= 1'h0;
		else if (_0011_)
			_0382_ <= \mchip.M1.IN_REG.SHIFT.Q [1];
	always @(posedge io_in[12])
		if (io_in[13])
			_0383_ <= 1'h0;
		else if (_0011_)
			_0383_ <= \mchip.M1.IN_REG.SHIFT.Q [2];
	always @(posedge io_in[12])
		if (io_in[13])
			_0384_ <= 1'h0;
		else if (_0011_)
			_0384_ <= \mchip.M1.IN_REG.SHIFT.Q [3];
	always @(posedge io_in[12])
		if (io_in[13])
			_0385_ <= 1'h0;
		else if (_0011_)
			_0385_ <= \mchip.M1.IN_REG.SHIFT.Q [4];
	always @(posedge io_in[12])
		if (io_in[13])
			_0386_ <= 1'h0;
		else if (_0011_)
			_0386_ <= \mchip.M1.IN_REG.SHIFT.Q [5];
	always @(posedge io_in[12])
		if (io_in[13])
			_0387_ <= 1'h0;
		else if (_0011_)
			_0387_ <= \mchip.M1.IN_REG.SHIFT.Q [6];
	always @(posedge io_in[12])
		if (io_in[13])
			_0388_ <= 1'h0;
		else if (_0011_)
			_0388_ <= \mchip.M1.IN_REG.SHIFT.Q [7];
	always @(posedge io_in[12])
		if (io_in[13])
			_0389_ <= 1'h0;
		else if (!_0120_)
			_0389_ <= _0103_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0390_ <= 1'h0;
		else if (!_0120_)
			_0390_ <= _0109_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0391_ <= 1'h0;
		else if (!_0120_)
			_0391_ <= _0110_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0392_ <= 1'h0;
		else if (!_0120_)
			_0392_ <= _0111_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0393_ <= 1'h0;
		else if (!_0120_)
			_0393_ <= _0112_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0394_ <= 1'h0;
		else if (!_0120_)
			_0394_ <= _0113_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0395_ <= 1'h0;
		else if (!_0120_)
			_0395_ <= _0114_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0396_ <= 1'h0;
		else if (!_0120_)
			_0396_ <= _0115_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0397_ <= 1'h0;
		else if (!_0120_)
			_0397_ <= _0116_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0398_ <= 1'h1;
		else if (!_0120_)
			_0398_ <= _0117_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0399_ <= 1'h1;
		else if (!_0120_)
			_0399_ <= _0104_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0400_ <= 1'h1;
		else if (!_0120_)
			_0400_ <= _0105_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0401_ <= 1'h1;
		else if (!_0120_)
			_0401_ <= _0106_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0402_ <= 1'h1;
		else if (!_0120_)
			_0402_ <= _0107_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0403_ <= 1'h1;
		else if (!_0120_)
			_0403_ <= _0108_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0404_ <= 1'h1;
		else if (!_0120_)
			_0404_ <= _0035_;
	always @(posedge io_in[12]) \mchip.M1.S1.m1.Q  <= io_in[0];
	assign _1889_[3:1] = \mchip.M1.COUNT.count [3:1];
	assign _1890_[0] = _1889_[0];
	assign {io_out[13:12], io_out[3:0]} = {2'h0, \mchip.M2.PWM2 , \mchip.M2.PWM1 , \mchip.M2.UART_DRIVER.tx , \mchip.SDA_out };
	assign \mchip.M1.ACK  = \mchip.M1.READ_ACK.ACK ;
	assign \mchip.M1.ADDR.addr  = 7'h20;
	assign \mchip.M1.ADDR.addr_sel  = io_in[3:2];
	assign \mchip.M1.ADDR.data_in  = \mchip.M1.IN_REG.SHIFT.Q [7:1];
	assign \mchip.M1.COUNT.clock  = io_in[12];
	assign \mchip.M1.COUNT.en  = \mchip.M1.S1.EDGE.sig_posedge ;
	assign \mchip.M1.IN_REG.SCL_posedge  = \mchip.M1.S1.EDGE.sig_posedge ;
	assign \mchip.M1.IN_REG.SDA  = \mchip.M1.S2.EDGE.prev ;
	assign \mchip.M1.IN_REG.SHIFT.Q [0] = \mchip.M1.M.read_write ;
	assign \mchip.M1.IN_REG.SHIFT.clock  = io_in[12];
	assign \mchip.M1.IN_REG.SHIFT.reset  = io_in[13];
	assign \mchip.M1.IN_REG.SHIFT.serial  = \mchip.M1.S2.EDGE.prev ;
	assign \mchip.M1.IN_REG.clock  = io_in[12];
	assign \mchip.M1.IN_REG.data_in  = {\mchip.M1.IN_REG.SHIFT.Q [7:1], \mchip.M1.M.read_write };
	assign \mchip.M1.IN_REG.reset  = io_in[13];
	assign \mchip.M1.M.ACK  = \mchip.M1.READ_ACK.ACK ;
	assign \mchip.M1.M.SCL_negedge  = \mchip.M1.S1.EDGE.sig_negedge ;
	assign \mchip.M1.M.clear_counter  = \mchip.M1.COUNT.clear ;
	assign \mchip.M1.M.clock  = io_in[12];
	assign \mchip.M1.M.currState [10] = 1'h0;
	assign \mchip.M1.M.data_in  = {\mchip.M1.IN_REG.SHIFT.Q [7:1], \mchip.M1.M.read_write };
	assign \mchip.M1.M.out_en  = \mchip.M1.M.currState [1];
	assign \mchip.M1.M.reg_sel_en  = \mchip.M1.M.currState [5];
	assign \mchip.M1.M.reset  = io_in[13];
	assign \mchip.M1.MEM.SCL_negedge  = \mchip.M1.S1.EDGE.sig_negedge ;
	assign \mchip.M1.MEM.clock  = io_in[12];
	assign \mchip.M1.MEM.count  = \mchip.M1.COUNT.count [2:0];
	assign \mchip.M1.MEM.data_in  = {\mchip.M1.IN_REG.SHIFT.Q [7:1], \mchip.M1.M.read_write };
	assign \mchip.M1.MEM.j  = 32'd24;
	assign \mchip.M1.MEM.parallel_in  = io_in[11:4];
	assign \mchip.M1.MEM.reg_out  = io_out[11:4];
	assign \mchip.M1.MEM.registers[1]  = io_out[11:4];
	assign \mchip.M1.MEM.registers_packed [15:0] = {io_out[11:4], \mchip.M1.MEM.registers[0] };
	assign \mchip.M1.MEM.reset  = io_in[13];
	assign \mchip.M1.OUT.out_en  = \mchip.M1.M.currState [1];
	assign \mchip.M1.READ_ACK.SCL_posedge  = \mchip.M1.S1.EDGE.sig_posedge ;
	assign \mchip.M1.READ_ACK.SDA  = \mchip.M1.S2.EDGE.prev ;
	assign \mchip.M1.READ_ACK.clock  = io_in[12];
	assign \mchip.M1.REG.SCL_negedge  = \mchip.M1.S1.EDGE.sig_negedge ;
	assign \mchip.M1.REG.clock  = io_in[12];
	assign \mchip.M1.REG.en  = \mchip.M1.M.currState [5];
	assign \mchip.M1.REG.reset  = io_in[13];
	assign \mchip.M1.REG.sel_in  = {\mchip.M1.IN_REG.SHIFT.Q [4:1], \mchip.M1.M.read_write };
	assign \mchip.M1.S1.EDGE.clock  = io_in[12];
	assign \mchip.M1.S1.EDGE.sig  = \mchip.M1.S1.m1.Q ;
	assign \mchip.M1.S1.EDGE.sig_out  = \mchip.M1.S1.EDGE.prev ;
	assign \mchip.M1.S1.async  = io_in[0];
	assign \mchip.M1.S1.clock  = io_in[12];
	assign \mchip.M1.S1.m1.D  = io_in[0];
	assign \mchip.M1.S1.m1.clock  = io_in[12];
	assign \mchip.M1.S1.sig_negedge  = \mchip.M1.S1.EDGE.sig_negedge ;
	assign \mchip.M1.S1.sig_posedge  = \mchip.M1.S1.EDGE.sig_posedge ;
	assign \mchip.M1.S1.sync  = \mchip.M1.S1.EDGE.prev ;
	assign \mchip.M1.S1.temp  = \mchip.M1.S1.m1.Q ;
	assign \mchip.M1.S2.EDGE.clock  = io_in[12];
	assign \mchip.M1.S2.EDGE.sig  = \mchip.M1.S2.m1.Q ;
	assign \mchip.M1.S2.EDGE.sig_out  = \mchip.M1.S2.EDGE.prev ;
	assign \mchip.M1.S2.async  = io_in[1];
	assign \mchip.M1.S2.clock  = io_in[12];
	assign \mchip.M1.S2.m1.D  = io_in[1];
	assign \mchip.M1.S2.m1.clock  = io_in[12];
	assign \mchip.M1.S2.sig_negedge  = \mchip.M1.S2.EDGE.sig_negedge ;
	assign \mchip.M1.S2.sig_posedge  = \mchip.M1.S2.EDGE.sig_posedge ;
	assign \mchip.M1.S2.sync  = \mchip.M1.S2.EDGE.prev ;
	assign \mchip.M1.S2.temp  = \mchip.M1.S2.m1.Q ;
	assign \mchip.M1.SCL_in  = io_in[0];
	assign \mchip.M1.SCL_negedge  = \mchip.M1.S1.EDGE.sig_negedge ;
	assign \mchip.M1.SCL_posedge  = \mchip.M1.S1.EDGE.sig_posedge ;
	assign \mchip.M1.SCL_sync  = \mchip.M1.S1.EDGE.prev ;
	assign \mchip.M1.SDA_in  = io_in[1];
	assign \mchip.M1.SDA_negedge  = \mchip.M1.S2.EDGE.sig_negedge ;
	assign \mchip.M1.SDA_posedge  = \mchip.M1.S2.EDGE.sig_posedge ;
	assign \mchip.M1.SDA_sync  = \mchip.M1.S2.EDGE.prev ;
	assign \mchip.M1.START.SCL  = \mchip.M1.S1.EDGE.prev ;
	assign \mchip.M1.START.SDA_negedge  = \mchip.M1.S2.EDGE.sig_negedge ;
	assign \mchip.M1.START.clock  = io_in[12];
	assign \mchip.M1.STOP.SCL  = \mchip.M1.S1.EDGE.prev ;
	assign \mchip.M1.STOP.SDA_posedge  = \mchip.M1.S2.EDGE.sig_posedge ;
	assign \mchip.M1.STOP.clock  = io_in[12];
	assign \mchip.M1.addr_sel  = io_in[3:2];
	assign \mchip.M1.clear_counter  = \mchip.M1.COUNT.clear ;
	assign \mchip.M1.clock  = io_in[12];
	assign \mchip.M1.count  = \mchip.M1.COUNT.count ;
	assign \mchip.M1.data_in  = {\mchip.M1.IN_REG.SHIFT.Q [7:1], \mchip.M1.M.read_write };
	assign \mchip.M1.out_en  = \mchip.M1.M.currState [1];
	assign \mchip.M1.parallel_in  = io_in[11:4];
	assign \mchip.M1.reg_out  = io_out[11:4];
	assign \mchip.M1.reg_sel_en  = \mchip.M1.M.currState [5];
	assign \mchip.M1.registers_packed [15:0] = {io_out[11:4], \mchip.M1.MEM.registers[0] };
	assign \mchip.M1.reset  = io_in[13];
	assign \mchip.M2.PWM_DRIVER.P1.PWM_out  = \mchip.M2.PWM1 ;
	assign \mchip.M2.PWM_DRIVER.P1.clock  = io_in[12];
	assign \mchip.M2.PWM_DRIVER.P1.reset  = io_in[13];
	assign \mchip.M2.PWM_DRIVER.P2.PWM_out  = \mchip.M2.PWM2 ;
	assign \mchip.M2.PWM_DRIVER.P2.clock  = io_in[12];
	assign \mchip.M2.PWM_DRIVER.P2.reset  = io_in[13];
	assign \mchip.M2.PWM_DRIVER.PWM1  = \mchip.M2.PWM1 ;
	assign \mchip.M2.PWM_DRIVER.PWM2  = \mchip.M2.PWM2 ;
	assign \mchip.M2.PWM_DRIVER.clock  = io_in[12];
	assign \mchip.M2.PWM_DRIVER.registers_packed [15:0] = {io_out[11:4], \mchip.M1.MEM.registers[0] };
	assign \mchip.M2.PWM_DRIVER.reset  = io_in[13];
	assign \mchip.M2.UART_DRIVER.clock  = io_in[12];
	assign \mchip.M2.UART_DRIVER.data  = io_out[11:4];
	assign \mchip.M2.UART_DRIVER.frame [0] = \mchip.M2.UART_DRIVER.tx ;
	assign \mchip.M2.UART_DRIVER.reset  = io_in[13];
	assign \mchip.M2.clock  = io_in[12];
	assign \mchip.M2.data_out  = {io_out[11:4], \mchip.M2.PWM2 , \mchip.M2.PWM1 , \mchip.M2.UART_DRIVER.tx };
	assign \mchip.M2.reg_out  = io_out[11:4];
	assign \mchip.M2.registers_packed [15:0] = {io_out[11:4], \mchip.M1.MEM.registers[0] };
	assign \mchip.M2.reset  = io_in[13];
	assign \mchip.M2.tx  = \mchip.M2.UART_DRIVER.tx ;
	assign \mchip.SCL_in  = io_in[0];
	assign \mchip.SDA_in  = io_in[1];
	assign \mchip.clock  = io_in[12];
	assign \mchip.data_out  = {io_out[11:4], \mchip.M2.PWM2 , \mchip.M2.PWM1 , \mchip.M2.UART_DRIVER.tx };
	assign \mchip.io_in  = io_in[11:0];
	assign \mchip.io_out  = {io_out[11:4], \mchip.M2.PWM2 , \mchip.M2.PWM1 , \mchip.M2.UART_DRIVER.tx , \mchip.SDA_out };
	assign \mchip.reg_out  = io_out[11:4];
	assign \mchip.registers_packed [15:0] = {io_out[11:4], \mchip.M1.MEM.registers[0] };
	assign \mchip.reset  = io_in[13];
endmodule
module d13_jrduvall_s444 (
	io_in,
	io_out
);
	wire _000_;
	wire _001_;
	wire _002_;
	wire _003_;
	wire _004_;
	wire _005_;
	wire _006_;
	wire _007_;
	wire _008_;
	wire _009_;
	wire _010_;
	wire _011_;
	wire _012_;
	wire _013_;
	wire _014_;
	wire _015_;
	wire _016_;
	wire _017_;
	wire _018_;
	wire _019_;
	wire _020_;
	wire _021_;
	wire _022_;
	wire _023_;
	wire _024_;
	wire _025_;
	wire _026_;
	wire _027_;
	wire _028_;
	wire _029_;
	wire _030_;
	wire _031_;
	wire _032_;
	wire _033_;
	wire _034_;
	wire _035_;
	wire _036_;
	wire _037_;
	wire _038_;
	wire _039_;
	wire _040_;
	wire _041_;
	wire _042_;
	wire _043_;
	wire _044_;
	wire _045_;
	wire _046_;
	wire _047_;
	wire _048_;
	wire _049_;
	wire _050_;
	input wire [13:0] io_in;
	output wire [13:0] io_out;
	wire \mchip.clock ;
	wire [11:0] \mchip.io_in ;
	wire [11:0] \mchip.io_out ;
	wire \mchip.reset ;
	wire \mchip.s444.c_in ;
	wire \mchip.s444.c_out ;
	wire \mchip.s444.carry_logic.c_in ;
	wire \mchip.s444.carry_logic.c_out ;
	wire \mchip.s444.carry_logic.gen ;
	wire \mchip.s444.carry_logic.prop ;
	wire \mchip.s444.carry_logic.sum_out ;
	wire \mchip.s444.clk ;
	wire \mchip.s444.d_flip_flops.clk ;
	wire [1:0] \mchip.s444.d_flip_flops.dff.D ;
	reg [1:0] \mchip.s444.d_flip_flops.dff.Q ;
	wire \mchip.s444.d_flip_flops.dff.clear ;
	wire \mchip.s444.d_flip_flops.dff.clock ;
	wire \mchip.s444.d_flip_flops.dff.en ;
	wire \mchip.s444.d_flip_flops.dff.load ;
	wire \mchip.s444.d_flip_flops.dff0 ;
	wire [3:0] \mchip.s444.d_flip_flops.dff0_mux.D ;
	wire [1:0] \mchip.s444.d_flip_flops.dff0_mux.I ;
	wire \mchip.s444.d_flip_flops.dff0_mux.O ;
	wire \mchip.s444.d_flip_flops.dff0_out ;
	wire [1:0] \mchip.s444.d_flip_flops.dff0_sel ;
	wire \mchip.s444.d_flip_flops.dff1 ;
	wire [3:0] \mchip.s444.d_flip_flops.dff1_mux.D ;
	wire [1:0] \mchip.s444.d_flip_flops.dff1_mux.I ;
	wire \mchip.s444.d_flip_flops.dff1_mux.O ;
	wire \mchip.s444.d_flip_flops.dff1_out ;
	wire [1:0] \mchip.s444.d_flip_flops.dff1_sel ;
	wire \mchip.s444.d_flip_flops.dff_reg.I ;
	wire \mchip.s444.d_flip_flops.dff_reg.O ;
	wire [3:0] \mchip.s444.d_flip_flops.dff_reg.Q ;
	wire \mchip.s444.d_flip_flops.dff_reg.clock ;
	wire \mchip.s444.d_flip_flops.dff_reg.en ;
	wire \mchip.s444.d_flip_flops.dff_reg.highBit ;
	wire \mchip.s444.d_flip_flops.dff_reg.left ;
	wire \mchip.s444.d_flip_flops.dff_reg.lowBit ;
	wire [3:0] \mchip.s444.d_flip_flops.dff_reg.myLatch.D ;
	reg [3:0] \mchip.s444.d_flip_flops.dff_reg.myLatch.Q ;
	wire \mchip.s444.d_flip_flops.dff_reg.myLatch.clear ;
	wire \mchip.s444.d_flip_flops.dff_reg.myLatch.clock ;
	wire \mchip.s444.d_flip_flops.dff_reg.myLatch.en ;
	wire \mchip.s444.d_flip_flops.dff_reg.myLatch.load ;
	wire \mchip.s444.d_flip_flops.dff_reg.reset ;
	wire \mchip.s444.d_flip_flops.dff_reg.shift ;
	wire [3:0] \mchip.s444.d_flip_flops.dff_reg.shiftResult ;
	wire [3:0] \mchip.s444.d_flip_flops.dff_reg.shiftedLeft ;
	wire \mchip.s444.d_flip_flops.en ;
	wire \mchip.s444.d_flip_flops.feed0_0 ;
	wire \mchip.s444.d_flip_flops.feed0_out ;
	wire \mchip.s444.d_flip_flops.feed1_0 ;
	wire \mchip.s444.d_flip_flops.feed1_out ;
	wire \mchip.s444.d_flip_flops.main_out ;
	wire \mchip.s444.d_flip_flops.reset ;
	wire \mchip.s444.d_flip_flops.shift_in ;
	wire \mchip.s444.d_flip_flops.shift_out ;
	wire \mchip.s444.d_flip_flops.sum_out ;
	wire \mchip.s444.dff0_out ;
	wire \mchip.s444.dff1_out ;
	wire \mchip.s444.en ;
	wire [3:0] \mchip.s444.feed0 ;
	wire \mchip.s444.feed0_out ;
	wire [3:0] \mchip.s444.feed1 ;
	wire \mchip.s444.feed1_out ;
	wire \mchip.s444.lut1 ;
	wire \mchip.s444.lut2 ;
	wire \mchip.s444.lut5_mux.clk ;
	wire \mchip.s444.lut5_mux.en ;
	wire \mchip.s444.lut5_mux.feed0_out ;
	wire \mchip.s444.lut5_mux.feed1_3 ;
	wire \mchip.s444.lut5_mux.lut1 ;
	wire \mchip.s444.lut5_mux.lut5_reg.I ;
	wire \mchip.s444.lut5_mux.lut5_reg.O ;
	wire \mchip.s444.lut5_mux.lut5_reg.Q ;
	wire \mchip.s444.lut5_mux.lut5_reg.clock ;
	wire \mchip.s444.lut5_mux.lut5_reg.en ;
	wire \mchip.s444.lut5_mux.lut5_reg.highBit ;
	wire \mchip.s444.lut5_mux.lut5_reg.left ;
	wire \mchip.s444.lut5_mux.lut5_reg.lowBit ;
	wire \mchip.s444.lut5_mux.lut5_reg.myLatch.D ;
	reg \mchip.s444.lut5_mux.lut5_reg.myLatch.Q ;
	wire \mchip.s444.lut5_mux.lut5_reg.myLatch.clear ;
	wire \mchip.s444.lut5_mux.lut5_reg.myLatch.clock ;
	wire \mchip.s444.lut5_mux.lut5_reg.myLatch.en ;
	wire \mchip.s444.lut5_mux.lut5_reg.myLatch.load ;
	wire \mchip.s444.lut5_mux.lut5_reg.reset ;
	wire \mchip.s444.lut5_mux.lut5_reg.shift ;
	wire \mchip.s444.lut5_mux.lut5_reg.shiftResult ;
	wire \mchip.s444.lut5_mux.lut5_reg.shiftedLeft ;
	wire \mchip.s444.lut5_mux.lut5_reg.shiftedRight ;
	wire \mchip.s444.lut5_mux.lut5_sel ;
	wire \mchip.s444.lut5_mux.reset ;
	wire \mchip.s444.lut5_mux.shift_in ;
	wire \mchip.s444.lut5_mux.shift_out ;
	wire [3:0] \mchip.s444.main ;
	wire \mchip.s444.main_out ;
	wire \mchip.s444.reset ;
	wire \mchip.s444.s444_logic.clk ;
	wire \mchip.s444.s444_logic.en ;
	wire [3:0] \mchip.s444.s444_logic.feed0 ;
	wire [3:0] \mchip.s444.s444_logic.feed1 ;
	wire [3:0] \mchip.s444.s444_logic.feed2 ;
	wire [15:0] \mchip.s444.s444_logic.l0.D ;
	wire [3:0] \mchip.s444.s444_logic.l0.I ;
	wire [15:0] \mchip.s444.s444_logic.l0_dat ;
	wire \mchip.s444.s444_logic.l0_reg.I ;
	wire \mchip.s444.s444_logic.l0_reg.O ;
	wire [15:0] \mchip.s444.s444_logic.l0_reg.Q ;
	wire \mchip.s444.s444_logic.l0_reg.clock ;
	wire \mchip.s444.s444_logic.l0_reg.en ;
	wire \mchip.s444.s444_logic.l0_reg.highBit ;
	wire \mchip.s444.s444_logic.l0_reg.left ;
	wire \mchip.s444.s444_logic.l0_reg.lowBit ;
	wire [15:0] \mchip.s444.s444_logic.l0_reg.myLatch.D ;
	reg [15:0] \mchip.s444.s444_logic.l0_reg.myLatch.Q ;
	wire \mchip.s444.s444_logic.l0_reg.myLatch.clear ;
	wire \mchip.s444.s444_logic.l0_reg.myLatch.clock ;
	wire \mchip.s444.s444_logic.l0_reg.myLatch.en ;
	wire \mchip.s444.s444_logic.l0_reg.myLatch.load ;
	wire \mchip.s444.s444_logic.l0_reg.reset ;
	wire \mchip.s444.s444_logic.l0_reg.shift ;
	wire [15:0] \mchip.s444.s444_logic.l0_reg.shiftResult ;
	wire [15:0] \mchip.s444.s444_logic.l0_reg.shiftedLeft ;
	wire [15:0] \mchip.s444.s444_logic.l1.D ;
	wire [3:0] \mchip.s444.s444_logic.l1.I ;
	wire \mchip.s444.s444_logic.l1.O ;
	wire [15:0] \mchip.s444.s444_logic.l1_dat ;
	wire \mchip.s444.s444_logic.l1_reg.I ;
	wire \mchip.s444.s444_logic.l1_reg.O ;
	wire [15:0] \mchip.s444.s444_logic.l1_reg.Q ;
	wire \mchip.s444.s444_logic.l1_reg.clock ;
	wire \mchip.s444.s444_logic.l1_reg.en ;
	wire \mchip.s444.s444_logic.l1_reg.highBit ;
	wire \mchip.s444.s444_logic.l1_reg.left ;
	wire \mchip.s444.s444_logic.l1_reg.lowBit ;
	wire [15:0] \mchip.s444.s444_logic.l1_reg.myLatch.D ;
	reg [15:0] \mchip.s444.s444_logic.l1_reg.myLatch.Q ;
	wire \mchip.s444.s444_logic.l1_reg.myLatch.clear ;
	wire \mchip.s444.s444_logic.l1_reg.myLatch.clock ;
	wire \mchip.s444.s444_logic.l1_reg.myLatch.en ;
	wire \mchip.s444.s444_logic.l1_reg.myLatch.load ;
	wire \mchip.s444.s444_logic.l1_reg.reset ;
	wire \mchip.s444.s444_logic.l1_reg.shift ;
	wire [15:0] \mchip.s444.s444_logic.l1_reg.shiftResult ;
	wire [15:0] \mchip.s444.s444_logic.l1_reg.shiftedLeft ;
	wire [15:0] \mchip.s444.s444_logic.l2.D ;
	wire [3:0] \mchip.s444.s444_logic.l2.I ;
	wire \mchip.s444.s444_logic.l2.O ;
	wire [15:0] \mchip.s444.s444_logic.l2_dat ;
	wire \mchip.s444.s444_logic.l2_reg.I ;
	wire \mchip.s444.s444_logic.l2_reg.O ;
	wire [15:0] \mchip.s444.s444_logic.l2_reg.Q ;
	wire \mchip.s444.s444_logic.l2_reg.clock ;
	wire \mchip.s444.s444_logic.l2_reg.en ;
	wire \mchip.s444.s444_logic.l2_reg.highBit ;
	wire \mchip.s444.s444_logic.l2_reg.left ;
	wire \mchip.s444.s444_logic.l2_reg.lowBit ;
	wire [15:0] \mchip.s444.s444_logic.l2_reg.myLatch.D ;
	reg [15:0] \mchip.s444.s444_logic.l2_reg.myLatch.Q ;
	wire \mchip.s444.s444_logic.l2_reg.myLatch.clear ;
	wire \mchip.s444.s444_logic.l2_reg.myLatch.clock ;
	wire \mchip.s444.s444_logic.l2_reg.myLatch.en ;
	wire \mchip.s444.s444_logic.l2_reg.myLatch.load ;
	wire \mchip.s444.s444_logic.l2_reg.reset ;
	wire \mchip.s444.s444_logic.l2_reg.shift ;
	wire [15:0] \mchip.s444.s444_logic.l2_reg.shiftResult ;
	wire [15:0] \mchip.s444.s444_logic.l2_reg.shiftedLeft ;
	wire \mchip.s444.s444_logic.lut1 ;
	wire \mchip.s444.s444_logic.lut2 ;
	wire \mchip.s444.s444_logic.m0_reg.I ;
	wire \mchip.s444.s444_logic.m0_reg.O ;
	wire \mchip.s444.s444_logic.m0_reg.Q ;
	wire \mchip.s444.s444_logic.m0_reg.clock ;
	wire \mchip.s444.s444_logic.m0_reg.en ;
	wire \mchip.s444.s444_logic.m0_reg.highBit ;
	wire \mchip.s444.s444_logic.m0_reg.left ;
	wire \mchip.s444.s444_logic.m0_reg.lowBit ;
	wire \mchip.s444.s444_logic.m0_reg.myLatch.D ;
	reg \mchip.s444.s444_logic.m0_reg.myLatch.Q ;
	wire \mchip.s444.s444_logic.m0_reg.myLatch.clear ;
	wire \mchip.s444.s444_logic.m0_reg.myLatch.clock ;
	wire \mchip.s444.s444_logic.m0_reg.myLatch.en ;
	wire \mchip.s444.s444_logic.m0_reg.myLatch.load ;
	wire \mchip.s444.s444_logic.m0_reg.reset ;
	wire \mchip.s444.s444_logic.m0_reg.shift ;
	wire \mchip.s444.s444_logic.m0_reg.shiftResult ;
	wire \mchip.s444.s444_logic.m0_reg.shiftedLeft ;
	wire \mchip.s444.s444_logic.m0_reg.shiftedRight ;
	wire \mchip.s444.s444_logic.m0_sel ;
	wire \mchip.s444.s444_logic.m1_reg.I ;
	wire \mchip.s444.s444_logic.m1_reg.O ;
	wire \mchip.s444.s444_logic.m1_reg.Q ;
	wire \mchip.s444.s444_logic.m1_reg.clock ;
	wire \mchip.s444.s444_logic.m1_reg.en ;
	wire \mchip.s444.s444_logic.m1_reg.highBit ;
	wire \mchip.s444.s444_logic.m1_reg.left ;
	wire \mchip.s444.s444_logic.m1_reg.lowBit ;
	wire \mchip.s444.s444_logic.m1_reg.myLatch.D ;
	reg \mchip.s444.s444_logic.m1_reg.myLatch.Q ;
	wire \mchip.s444.s444_logic.m1_reg.myLatch.clear ;
	wire \mchip.s444.s444_logic.m1_reg.myLatch.clock ;
	wire \mchip.s444.s444_logic.m1_reg.myLatch.en ;
	wire \mchip.s444.s444_logic.m1_reg.myLatch.load ;
	wire \mchip.s444.s444_logic.m1_reg.reset ;
	wire \mchip.s444.s444_logic.m1_reg.shift ;
	wire \mchip.s444.s444_logic.m1_reg.shiftResult ;
	wire \mchip.s444.s444_logic.m1_reg.shiftedLeft ;
	wire \mchip.s444.s444_logic.m1_reg.shiftedRight ;
	wire \mchip.s444.s444_logic.m1_sel ;
	wire \mchip.s444.s444_logic.m2_reg.I ;
	wire \mchip.s444.s444_logic.m2_reg.O ;
	wire \mchip.s444.s444_logic.m2_reg.Q ;
	wire \mchip.s444.s444_logic.m2_reg.clock ;
	wire \mchip.s444.s444_logic.m2_reg.en ;
	wire \mchip.s444.s444_logic.m2_reg.highBit ;
	wire \mchip.s444.s444_logic.m2_reg.left ;
	wire \mchip.s444.s444_logic.m2_reg.lowBit ;
	wire \mchip.s444.s444_logic.m2_reg.myLatch.D ;
	reg \mchip.s444.s444_logic.m2_reg.myLatch.Q ;
	wire \mchip.s444.s444_logic.m2_reg.myLatch.clear ;
	wire \mchip.s444.s444_logic.m2_reg.myLatch.clock ;
	wire \mchip.s444.s444_logic.m2_reg.myLatch.en ;
	wire \mchip.s444.s444_logic.m2_reg.myLatch.load ;
	wire \mchip.s444.s444_logic.m2_reg.reset ;
	wire \mchip.s444.s444_logic.m2_reg.shift ;
	wire \mchip.s444.s444_logic.m2_reg.shiftResult ;
	wire \mchip.s444.s444_logic.m2_reg.shiftedLeft ;
	wire \mchip.s444.s444_logic.m2_reg.shiftedRight ;
	wire \mchip.s444.s444_logic.m2_sel ;
	wire [3:0] \mchip.s444.s444_logic.main ;
	wire \mchip.s444.s444_logic.reset ;
	wire \mchip.s444.s444_logic.shift_in ;
	wire \mchip.s444.s444_logic.shift_l0 ;
	wire \mchip.s444.s444_logic.shift_l1 ;
	wire \mchip.s444.s444_logic.shift_l2 ;
	wire \mchip.s444.s444_logic.shift_m0 ;
	wire \mchip.s444.s444_logic.shift_m1 ;
	wire \mchip.s444.s444_logic.shift_m2 ;
	wire \mchip.s444.s444_logic.shift_out ;
	wire \mchip.s444.shift0 ;
	wire \mchip.s444.shift1 ;
	wire \mchip.s444.shift_in ;
	wire \mchip.s444.shift_out ;
	wire \mchip.s444.sum_out ;
	assign _029_ = (io_in[0] ? \mchip.s444.s444_logic.l1_reg.myLatch.Q [1] : \mchip.s444.s444_logic.l1_reg.myLatch.Q [0]);
	assign _030_ = (io_in[0] ? \mchip.s444.s444_logic.l1_reg.myLatch.Q [3] : \mchip.s444.s444_logic.l1_reg.myLatch.Q [2]);
	assign _031_ = (io_in[1] ? _030_ : _029_);
	assign _032_ = (io_in[0] ? \mchip.s444.s444_logic.l1_reg.myLatch.Q [5] : \mchip.s444.s444_logic.l1_reg.myLatch.Q [4]);
	assign _033_ = (io_in[0] ? \mchip.s444.s444_logic.l1_reg.myLatch.Q [7] : \mchip.s444.s444_logic.l1_reg.myLatch.Q [6]);
	assign _034_ = (io_in[1] ? _033_ : _032_);
	assign _035_ = (io_in[2] ? _034_ : _031_);
	assign _036_ = (\mchip.s444.s444_logic.m2_reg.myLatch.Q  ? io_in[3] : io_in[4]);
	assign _037_ = (io_in[0] ? \mchip.s444.s444_logic.l1_reg.myLatch.Q [9] : \mchip.s444.s444_logic.l1_reg.myLatch.Q [8]);
	assign _038_ = (io_in[0] ? \mchip.s444.s444_logic.l1_reg.myLatch.Q [11] : \mchip.s444.s444_logic.l1_reg.myLatch.Q [10]);
	assign _039_ = (io_in[1] ? _038_ : _037_);
	assign _040_ = (io_in[0] ? \mchip.s444.s444_logic.l1_reg.myLatch.Q [13] : \mchip.s444.s444_logic.l1_reg.myLatch.Q [12]);
	assign _041_ = (io_in[0] ? \mchip.s444.s444_logic.l1_reg.myLatch.Q [15] : \mchip.s444.s444_logic.l1_reg.myLatch.Q [14]);
	assign _042_ = (io_in[1] ? _041_ : _040_);
	assign _043_ = (io_in[2] ? _042_ : _039_);
	assign \mchip.s444.carry_logic.prop  = (_036_ ? _043_ : _035_);
	assign _044_ = (io_in[5] ? \mchip.s444.s444_logic.l2_reg.myLatch.Q [1] : \mchip.s444.s444_logic.l2_reg.myLatch.Q [0]);
	assign _045_ = (io_in[5] ? \mchip.s444.s444_logic.l2_reg.myLatch.Q [3] : \mchip.s444.s444_logic.l2_reg.myLatch.Q [2]);
	assign _046_ = (io_in[6] ? _045_ : _044_);
	assign _047_ = (\mchip.s444.s444_logic.m1_reg.myLatch.Q  ? io_in[7] : \mchip.s444.carry_logic.prop );
	assign _048_ = (io_in[5] ? \mchip.s444.s444_logic.l2_reg.myLatch.Q [5] : \mchip.s444.s444_logic.l2_reg.myLatch.Q [4]);
	assign _049_ = (io_in[5] ? \mchip.s444.s444_logic.l2_reg.myLatch.Q [7] : \mchip.s444.s444_logic.l2_reg.myLatch.Q [6]);
	assign _050_ = (io_in[6] ? _049_ : _048_);
	assign _000_ = (_047_ ? _050_ : _046_);
	assign _001_ = (io_in[0] ? \mchip.s444.s444_logic.l0_reg.myLatch.Q [1] : \mchip.s444.s444_logic.l0_reg.myLatch.Q [0]);
	assign _002_ = (io_in[0] ? \mchip.s444.s444_logic.l0_reg.myLatch.Q [3] : \mchip.s444.s444_logic.l0_reg.myLatch.Q [2]);
	assign _003_ = (io_in[1] ? _002_ : _001_);
	assign _004_ = (io_in[0] ? \mchip.s444.s444_logic.l0_reg.myLatch.Q [5] : \mchip.s444.s444_logic.l0_reg.myLatch.Q [4]);
	assign _005_ = (io_in[0] ? \mchip.s444.s444_logic.l0_reg.myLatch.Q [7] : \mchip.s444.s444_logic.l0_reg.myLatch.Q [6]);
	assign _006_ = (io_in[1] ? _005_ : _004_);
	assign _007_ = (io_in[2] ? _006_ : _003_);
	assign _008_ = (io_in[0] ? \mchip.s444.s444_logic.l0_reg.myLatch.Q [9] : \mchip.s444.s444_logic.l0_reg.myLatch.Q [8]);
	assign _009_ = (io_in[0] ? \mchip.s444.s444_logic.l0_reg.myLatch.Q [11] : \mchip.s444.s444_logic.l0_reg.myLatch.Q [10]);
	assign _010_ = (io_in[1] ? _009_ : _008_);
	assign _011_ = (io_in[0] ? \mchip.s444.s444_logic.l0_reg.myLatch.Q [13] : \mchip.s444.s444_logic.l0_reg.myLatch.Q [12]);
	assign _012_ = (io_in[0] ? \mchip.s444.s444_logic.l0_reg.myLatch.Q [15] : \mchip.s444.s444_logic.l0_reg.myLatch.Q [14]);
	assign _013_ = (io_in[1] ? _012_ : _011_);
	assign _014_ = (io_in[2] ? _013_ : _010_);
	assign _015_ = (io_in[3] ? _014_ : _007_);
	assign _016_ = (\mchip.s444.s444_logic.m0_reg.myLatch.Q  ? io_in[8] : _015_);
	assign _017_ = (io_in[5] ? \mchip.s444.s444_logic.l2_reg.myLatch.Q [9] : \mchip.s444.s444_logic.l2_reg.myLatch.Q [8]);
	assign _018_ = (io_in[5] ? \mchip.s444.s444_logic.l2_reg.myLatch.Q [11] : \mchip.s444.s444_logic.l2_reg.myLatch.Q [10]);
	assign _019_ = (io_in[6] ? _018_ : _017_);
	assign _020_ = (io_in[5] ? \mchip.s444.s444_logic.l2_reg.myLatch.Q [13] : \mchip.s444.s444_logic.l2_reg.myLatch.Q [12]);
	assign _021_ = (io_in[5] ? \mchip.s444.s444_logic.l2_reg.myLatch.Q [15] : \mchip.s444.s444_logic.l2_reg.myLatch.Q [14]);
	assign _022_ = (io_in[6] ? _021_ : _020_);
	assign _023_ = (_047_ ? _022_ : _019_);
	assign \mchip.s444.carry_logic.gen  = (_016_ ? _023_ : _000_);
	assign \mchip.s444.c_out  = (\mchip.s444.carry_logic.prop  ? io_in[9] : \mchip.s444.carry_logic.gen );
	assign _024_ = \mchip.s444.lut5_mux.lut5_reg.myLatch.Q  & io_in[4];
	assign \mchip.s444.d_flip_flops.feed0_out  = (_024_ ? \mchip.s444.carry_logic.prop  : _015_);
	assign \mchip.s444.carry_logic.sum_out  = \mchip.s444.carry_logic.prop  ^ io_in[9];
	assign _025_ = \mchip.s444.carry_logic.prop  & ~\mchip.s444.d_flip_flops.dff_reg.myLatch.Q [2];
	assign _026_ = (\mchip.s444.d_flip_flops.dff_reg.myLatch.Q [2] ? \mchip.s444.carry_logic.sum_out  : io_in[0]);
	assign \mchip.s444.d_flip_flops.dff1  = (\mchip.s444.d_flip_flops.dff_reg.myLatch.Q [3] ? _026_ : _025_);
	assign _027_ = \mchip.s444.d_flip_flops.feed0_out  & ~\mchip.s444.d_flip_flops.dff_reg.myLatch.Q [0];
	assign _028_ = (\mchip.s444.d_flip_flops.dff_reg.myLatch.Q [0] ? \mchip.s444.carry_logic.sum_out  : io_in[0]);
	assign \mchip.s444.d_flip_flops.dff0  = (\mchip.s444.d_flip_flops.dff_reg.myLatch.Q [1] ? _028_ : _027_);
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.s444.d_flip_flops.dff.Q [0] <= 1'h0;
		else
			\mchip.s444.d_flip_flops.dff.Q [0] <= \mchip.s444.d_flip_flops.dff0 ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.s444.d_flip_flops.dff.Q [1] <= 1'h0;
		else
			\mchip.s444.d_flip_flops.dff.Q [1] <= \mchip.s444.d_flip_flops.dff1 ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.s444.s444_logic.l2_reg.myLatch.Q [0] <= 1'h0;
		else if (io_in[11])
			\mchip.s444.s444_logic.l2_reg.myLatch.Q [0] <= \mchip.s444.s444_logic.l1_reg.myLatch.Q [15];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.s444.s444_logic.l2_reg.myLatch.Q [1] <= 1'h0;
		else if (io_in[11])
			\mchip.s444.s444_logic.l2_reg.myLatch.Q [1] <= \mchip.s444.s444_logic.l2_reg.myLatch.Q [0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.s444.s444_logic.l2_reg.myLatch.Q [2] <= 1'h0;
		else if (io_in[11])
			\mchip.s444.s444_logic.l2_reg.myLatch.Q [2] <= \mchip.s444.s444_logic.l2_reg.myLatch.Q [1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.s444.s444_logic.l2_reg.myLatch.Q [3] <= 1'h0;
		else if (io_in[11])
			\mchip.s444.s444_logic.l2_reg.myLatch.Q [3] <= \mchip.s444.s444_logic.l2_reg.myLatch.Q [2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.s444.s444_logic.l2_reg.myLatch.Q [4] <= 1'h0;
		else if (io_in[11])
			\mchip.s444.s444_logic.l2_reg.myLatch.Q [4] <= \mchip.s444.s444_logic.l2_reg.myLatch.Q [3];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.s444.s444_logic.l2_reg.myLatch.Q [5] <= 1'h0;
		else if (io_in[11])
			\mchip.s444.s444_logic.l2_reg.myLatch.Q [5] <= \mchip.s444.s444_logic.l2_reg.myLatch.Q [4];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.s444.s444_logic.l2_reg.myLatch.Q [6] <= 1'h0;
		else if (io_in[11])
			\mchip.s444.s444_logic.l2_reg.myLatch.Q [6] <= \mchip.s444.s444_logic.l2_reg.myLatch.Q [5];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.s444.s444_logic.l2_reg.myLatch.Q [7] <= 1'h0;
		else if (io_in[11])
			\mchip.s444.s444_logic.l2_reg.myLatch.Q [7] <= \mchip.s444.s444_logic.l2_reg.myLatch.Q [6];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.s444.s444_logic.l2_reg.myLatch.Q [8] <= 1'h0;
		else if (io_in[11])
			\mchip.s444.s444_logic.l2_reg.myLatch.Q [8] <= \mchip.s444.s444_logic.l2_reg.myLatch.Q [7];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.s444.s444_logic.l2_reg.myLatch.Q [9] <= 1'h0;
		else if (io_in[11])
			\mchip.s444.s444_logic.l2_reg.myLatch.Q [9] <= \mchip.s444.s444_logic.l2_reg.myLatch.Q [8];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.s444.s444_logic.l2_reg.myLatch.Q [10] <= 1'h0;
		else if (io_in[11])
			\mchip.s444.s444_logic.l2_reg.myLatch.Q [10] <= \mchip.s444.s444_logic.l2_reg.myLatch.Q [9];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.s444.s444_logic.l2_reg.myLatch.Q [11] <= 1'h0;
		else if (io_in[11])
			\mchip.s444.s444_logic.l2_reg.myLatch.Q [11] <= \mchip.s444.s444_logic.l2_reg.myLatch.Q [10];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.s444.s444_logic.l2_reg.myLatch.Q [12] <= 1'h0;
		else if (io_in[11])
			\mchip.s444.s444_logic.l2_reg.myLatch.Q [12] <= \mchip.s444.s444_logic.l2_reg.myLatch.Q [11];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.s444.s444_logic.l2_reg.myLatch.Q [13] <= 1'h0;
		else if (io_in[11])
			\mchip.s444.s444_logic.l2_reg.myLatch.Q [13] <= \mchip.s444.s444_logic.l2_reg.myLatch.Q [12];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.s444.s444_logic.l2_reg.myLatch.Q [14] <= 1'h0;
		else if (io_in[11])
			\mchip.s444.s444_logic.l2_reg.myLatch.Q [14] <= \mchip.s444.s444_logic.l2_reg.myLatch.Q [13];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.s444.s444_logic.l2_reg.myLatch.Q [15] <= 1'h0;
		else if (io_in[11])
			\mchip.s444.s444_logic.l2_reg.myLatch.Q [15] <= \mchip.s444.s444_logic.l2_reg.myLatch.Q [14];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.s444.s444_logic.l1_reg.myLatch.Q [0] <= 1'h0;
		else if (io_in[11])
			\mchip.s444.s444_logic.l1_reg.myLatch.Q [0] <= \mchip.s444.s444_logic.l0_reg.myLatch.Q [15];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.s444.s444_logic.l1_reg.myLatch.Q [1] <= 1'h0;
		else if (io_in[11])
			\mchip.s444.s444_logic.l1_reg.myLatch.Q [1] <= \mchip.s444.s444_logic.l1_reg.myLatch.Q [0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.s444.s444_logic.l1_reg.myLatch.Q [2] <= 1'h0;
		else if (io_in[11])
			\mchip.s444.s444_logic.l1_reg.myLatch.Q [2] <= \mchip.s444.s444_logic.l1_reg.myLatch.Q [1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.s444.s444_logic.l1_reg.myLatch.Q [3] <= 1'h0;
		else if (io_in[11])
			\mchip.s444.s444_logic.l1_reg.myLatch.Q [3] <= \mchip.s444.s444_logic.l1_reg.myLatch.Q [2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.s444.s444_logic.l1_reg.myLatch.Q [4] <= 1'h0;
		else if (io_in[11])
			\mchip.s444.s444_logic.l1_reg.myLatch.Q [4] <= \mchip.s444.s444_logic.l1_reg.myLatch.Q [3];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.s444.s444_logic.l1_reg.myLatch.Q [5] <= 1'h0;
		else if (io_in[11])
			\mchip.s444.s444_logic.l1_reg.myLatch.Q [5] <= \mchip.s444.s444_logic.l1_reg.myLatch.Q [4];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.s444.s444_logic.l1_reg.myLatch.Q [6] <= 1'h0;
		else if (io_in[11])
			\mchip.s444.s444_logic.l1_reg.myLatch.Q [6] <= \mchip.s444.s444_logic.l1_reg.myLatch.Q [5];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.s444.s444_logic.l1_reg.myLatch.Q [7] <= 1'h0;
		else if (io_in[11])
			\mchip.s444.s444_logic.l1_reg.myLatch.Q [7] <= \mchip.s444.s444_logic.l1_reg.myLatch.Q [6];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.s444.s444_logic.l1_reg.myLatch.Q [8] <= 1'h0;
		else if (io_in[11])
			\mchip.s444.s444_logic.l1_reg.myLatch.Q [8] <= \mchip.s444.s444_logic.l1_reg.myLatch.Q [7];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.s444.s444_logic.l1_reg.myLatch.Q [9] <= 1'h0;
		else if (io_in[11])
			\mchip.s444.s444_logic.l1_reg.myLatch.Q [9] <= \mchip.s444.s444_logic.l1_reg.myLatch.Q [8];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.s444.s444_logic.l1_reg.myLatch.Q [10] <= 1'h0;
		else if (io_in[11])
			\mchip.s444.s444_logic.l1_reg.myLatch.Q [10] <= \mchip.s444.s444_logic.l1_reg.myLatch.Q [9];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.s444.s444_logic.l1_reg.myLatch.Q [11] <= 1'h0;
		else if (io_in[11])
			\mchip.s444.s444_logic.l1_reg.myLatch.Q [11] <= \mchip.s444.s444_logic.l1_reg.myLatch.Q [10];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.s444.s444_logic.l1_reg.myLatch.Q [12] <= 1'h0;
		else if (io_in[11])
			\mchip.s444.s444_logic.l1_reg.myLatch.Q [12] <= \mchip.s444.s444_logic.l1_reg.myLatch.Q [11];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.s444.s444_logic.l1_reg.myLatch.Q [13] <= 1'h0;
		else if (io_in[11])
			\mchip.s444.s444_logic.l1_reg.myLatch.Q [13] <= \mchip.s444.s444_logic.l1_reg.myLatch.Q [12];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.s444.s444_logic.l1_reg.myLatch.Q [14] <= 1'h0;
		else if (io_in[11])
			\mchip.s444.s444_logic.l1_reg.myLatch.Q [14] <= \mchip.s444.s444_logic.l1_reg.myLatch.Q [13];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.s444.s444_logic.l1_reg.myLatch.Q [15] <= 1'h0;
		else if (io_in[11])
			\mchip.s444.s444_logic.l1_reg.myLatch.Q [15] <= \mchip.s444.s444_logic.l1_reg.myLatch.Q [14];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.s444.s444_logic.l0_reg.myLatch.Q [0] <= 1'h0;
		else if (io_in[11])
			\mchip.s444.s444_logic.l0_reg.myLatch.Q [0] <= \mchip.s444.s444_logic.m2_reg.myLatch.Q ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.s444.s444_logic.l0_reg.myLatch.Q [1] <= 1'h0;
		else if (io_in[11])
			\mchip.s444.s444_logic.l0_reg.myLatch.Q [1] <= \mchip.s444.s444_logic.l0_reg.myLatch.Q [0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.s444.s444_logic.l0_reg.myLatch.Q [2] <= 1'h0;
		else if (io_in[11])
			\mchip.s444.s444_logic.l0_reg.myLatch.Q [2] <= \mchip.s444.s444_logic.l0_reg.myLatch.Q [1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.s444.s444_logic.l0_reg.myLatch.Q [3] <= 1'h0;
		else if (io_in[11])
			\mchip.s444.s444_logic.l0_reg.myLatch.Q [3] <= \mchip.s444.s444_logic.l0_reg.myLatch.Q [2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.s444.s444_logic.l0_reg.myLatch.Q [4] <= 1'h0;
		else if (io_in[11])
			\mchip.s444.s444_logic.l0_reg.myLatch.Q [4] <= \mchip.s444.s444_logic.l0_reg.myLatch.Q [3];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.s444.s444_logic.l0_reg.myLatch.Q [5] <= 1'h0;
		else if (io_in[11])
			\mchip.s444.s444_logic.l0_reg.myLatch.Q [5] <= \mchip.s444.s444_logic.l0_reg.myLatch.Q [4];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.s444.s444_logic.l0_reg.myLatch.Q [6] <= 1'h0;
		else if (io_in[11])
			\mchip.s444.s444_logic.l0_reg.myLatch.Q [6] <= \mchip.s444.s444_logic.l0_reg.myLatch.Q [5];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.s444.s444_logic.l0_reg.myLatch.Q [7] <= 1'h0;
		else if (io_in[11])
			\mchip.s444.s444_logic.l0_reg.myLatch.Q [7] <= \mchip.s444.s444_logic.l0_reg.myLatch.Q [6];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.s444.s444_logic.l0_reg.myLatch.Q [8] <= 1'h0;
		else if (io_in[11])
			\mchip.s444.s444_logic.l0_reg.myLatch.Q [8] <= \mchip.s444.s444_logic.l0_reg.myLatch.Q [7];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.s444.s444_logic.l0_reg.myLatch.Q [9] <= 1'h0;
		else if (io_in[11])
			\mchip.s444.s444_logic.l0_reg.myLatch.Q [9] <= \mchip.s444.s444_logic.l0_reg.myLatch.Q [8];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.s444.s444_logic.l0_reg.myLatch.Q [10] <= 1'h0;
		else if (io_in[11])
			\mchip.s444.s444_logic.l0_reg.myLatch.Q [10] <= \mchip.s444.s444_logic.l0_reg.myLatch.Q [9];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.s444.s444_logic.l0_reg.myLatch.Q [11] <= 1'h0;
		else if (io_in[11])
			\mchip.s444.s444_logic.l0_reg.myLatch.Q [11] <= \mchip.s444.s444_logic.l0_reg.myLatch.Q [10];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.s444.s444_logic.l0_reg.myLatch.Q [12] <= 1'h0;
		else if (io_in[11])
			\mchip.s444.s444_logic.l0_reg.myLatch.Q [12] <= \mchip.s444.s444_logic.l0_reg.myLatch.Q [11];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.s444.s444_logic.l0_reg.myLatch.Q [13] <= 1'h0;
		else if (io_in[11])
			\mchip.s444.s444_logic.l0_reg.myLatch.Q [13] <= \mchip.s444.s444_logic.l0_reg.myLatch.Q [12];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.s444.s444_logic.l0_reg.myLatch.Q [14] <= 1'h0;
		else if (io_in[11])
			\mchip.s444.s444_logic.l0_reg.myLatch.Q [14] <= \mchip.s444.s444_logic.l0_reg.myLatch.Q [13];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.s444.s444_logic.l0_reg.myLatch.Q [15] <= 1'h0;
		else if (io_in[11])
			\mchip.s444.s444_logic.l0_reg.myLatch.Q [15] <= \mchip.s444.s444_logic.l0_reg.myLatch.Q [14];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.s444.s444_logic.m2_reg.myLatch.Q  <= 1'h0;
		else if (io_in[11])
			\mchip.s444.s444_logic.m2_reg.myLatch.Q  <= \mchip.s444.s444_logic.m1_reg.myLatch.Q ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.s444.s444_logic.m1_reg.myLatch.Q  <= 1'h0;
		else if (io_in[11])
			\mchip.s444.s444_logic.m1_reg.myLatch.Q  <= \mchip.s444.s444_logic.m0_reg.myLatch.Q ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.s444.s444_logic.m0_reg.myLatch.Q  <= 1'h0;
		else if (io_in[11])
			\mchip.s444.s444_logic.m0_reg.myLatch.Q  <= io_in[10];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.s444.lut5_mux.lut5_reg.myLatch.Q  <= 1'h0;
		else if (io_in[11])
			\mchip.s444.lut5_mux.lut5_reg.myLatch.Q  <= \mchip.s444.s444_logic.l2_reg.myLatch.Q [15];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.s444.d_flip_flops.dff_reg.myLatch.Q [0] <= 1'h0;
		else if (io_in[11])
			\mchip.s444.d_flip_flops.dff_reg.myLatch.Q [0] <= \mchip.s444.lut5_mux.lut5_reg.myLatch.Q ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.s444.d_flip_flops.dff_reg.myLatch.Q [1] <= 1'h0;
		else if (io_in[11])
			\mchip.s444.d_flip_flops.dff_reg.myLatch.Q [1] <= \mchip.s444.d_flip_flops.dff_reg.myLatch.Q [0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.s444.d_flip_flops.dff_reg.myLatch.Q [2] <= 1'h0;
		else if (io_in[11])
			\mchip.s444.d_flip_flops.dff_reg.myLatch.Q [2] <= \mchip.s444.d_flip_flops.dff_reg.myLatch.Q [1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.s444.d_flip_flops.dff_reg.myLatch.Q [3] <= 1'h0;
		else if (io_in[11])
			\mchip.s444.d_flip_flops.dff_reg.myLatch.Q [3] <= \mchip.s444.d_flip_flops.dff_reg.myLatch.Q [2];
	assign io_out = {3'h0, \mchip.s444.d_flip_flops.dff_reg.myLatch.Q [3], \mchip.s444.c_out , \mchip.s444.carry_logic.sum_out , 3'h0, \mchip.s444.d_flip_flops.dff.Q , \mchip.s444.carry_logic.gen , \mchip.s444.carry_logic.prop , \mchip.s444.d_flip_flops.feed0_out };
	assign \mchip.clock  = io_in[12];
	assign \mchip.io_in  = io_in[11:0];
	assign \mchip.io_out  = {1'h0, \mchip.s444.d_flip_flops.dff_reg.myLatch.Q [3], \mchip.s444.c_out , \mchip.s444.carry_logic.sum_out , 3'h0, \mchip.s444.d_flip_flops.dff.Q , \mchip.s444.carry_logic.gen , \mchip.s444.carry_logic.prop , \mchip.s444.d_flip_flops.feed0_out };
	assign \mchip.reset  = io_in[13];
	assign \mchip.s444.c_in  = io_in[9];
	assign \mchip.s444.carry_logic.c_in  = io_in[9];
	assign \mchip.s444.carry_logic.c_out  = \mchip.s444.c_out ;
	assign \mchip.s444.clk  = io_in[12];
	assign \mchip.s444.d_flip_flops.clk  = io_in[12];
	assign \mchip.s444.d_flip_flops.dff.D  = {\mchip.s444.d_flip_flops.dff1 , \mchip.s444.d_flip_flops.dff0 };
	assign \mchip.s444.d_flip_flops.dff.clear  = io_in[13];
	assign \mchip.s444.d_flip_flops.dff.clock  = io_in[12];
	assign \mchip.s444.d_flip_flops.dff.en  = 1'h1;
	assign \mchip.s444.d_flip_flops.dff.load  = 1'h1;
	assign \mchip.s444.d_flip_flops.dff0_mux.D  = {\mchip.s444.carry_logic.sum_out , io_in[0], 1'h0, \mchip.s444.d_flip_flops.feed0_out };
	assign \mchip.s444.d_flip_flops.dff0_mux.I  = \mchip.s444.d_flip_flops.dff_reg.myLatch.Q [1:0];
	assign \mchip.s444.d_flip_flops.dff0_mux.O  = \mchip.s444.d_flip_flops.dff0 ;
	assign \mchip.s444.d_flip_flops.dff0_out  = \mchip.s444.d_flip_flops.dff.Q [0];
	assign \mchip.s444.d_flip_flops.dff0_sel  = \mchip.s444.d_flip_flops.dff_reg.myLatch.Q [1:0];
	assign \mchip.s444.d_flip_flops.dff1_mux.D  = {\mchip.s444.carry_logic.sum_out , io_in[0], 1'h0, \mchip.s444.carry_logic.prop };
	assign \mchip.s444.d_flip_flops.dff1_mux.I  = \mchip.s444.d_flip_flops.dff_reg.myLatch.Q [3:2];
	assign \mchip.s444.d_flip_flops.dff1_mux.O  = \mchip.s444.d_flip_flops.dff1 ;
	assign \mchip.s444.d_flip_flops.dff1_out  = \mchip.s444.d_flip_flops.dff.Q [1];
	assign \mchip.s444.d_flip_flops.dff1_sel  = \mchip.s444.d_flip_flops.dff_reg.myLatch.Q [3:2];
	assign \mchip.s444.d_flip_flops.dff_reg.I  = \mchip.s444.lut5_mux.lut5_reg.myLatch.Q ;
	assign \mchip.s444.d_flip_flops.dff_reg.O  = \mchip.s444.d_flip_flops.dff_reg.myLatch.Q [3];
	assign \mchip.s444.d_flip_flops.dff_reg.Q  = \mchip.s444.d_flip_flops.dff_reg.myLatch.Q ;
	assign \mchip.s444.d_flip_flops.dff_reg.clock  = io_in[12];
	assign \mchip.s444.d_flip_flops.dff_reg.en  = 1'h1;
	assign \mchip.s444.d_flip_flops.dff_reg.highBit  = \mchip.s444.d_flip_flops.dff_reg.myLatch.Q [3];
	assign \mchip.s444.d_flip_flops.dff_reg.left  = 1'h1;
	assign \mchip.s444.d_flip_flops.dff_reg.lowBit  = \mchip.s444.d_flip_flops.dff_reg.myLatch.Q [0];
	assign \mchip.s444.d_flip_flops.dff_reg.myLatch.D  = {\mchip.s444.d_flip_flops.dff_reg.myLatch.Q [2:0], \mchip.s444.lut5_mux.lut5_reg.myLatch.Q };
	assign \mchip.s444.d_flip_flops.dff_reg.myLatch.clear  = io_in[13];
	assign \mchip.s444.d_flip_flops.dff_reg.myLatch.clock  = io_in[12];
	assign \mchip.s444.d_flip_flops.dff_reg.myLatch.en  = 1'h1;
	assign \mchip.s444.d_flip_flops.dff_reg.myLatch.load  = io_in[11];
	assign \mchip.s444.d_flip_flops.dff_reg.reset  = io_in[13];
	assign \mchip.s444.d_flip_flops.dff_reg.shift  = io_in[11];
	assign \mchip.s444.d_flip_flops.dff_reg.shiftResult  = {\mchip.s444.d_flip_flops.dff_reg.myLatch.Q [2:0], \mchip.s444.lut5_mux.lut5_reg.myLatch.Q };
	assign \mchip.s444.d_flip_flops.dff_reg.shiftedLeft  = {\mchip.s444.d_flip_flops.dff_reg.myLatch.Q [2:0], \mchip.s444.lut5_mux.lut5_reg.myLatch.Q };
	assign \mchip.s444.d_flip_flops.en  = io_in[11];
	assign \mchip.s444.d_flip_flops.feed0_0  = io_in[0];
	assign \mchip.s444.d_flip_flops.feed1_0  = io_in[0];
	assign \mchip.s444.d_flip_flops.feed1_out  = \mchip.s444.carry_logic.prop ;
	assign \mchip.s444.d_flip_flops.main_out  = 1'h0;
	assign \mchip.s444.d_flip_flops.reset  = io_in[13];
	assign \mchip.s444.d_flip_flops.shift_in  = \mchip.s444.lut5_mux.lut5_reg.myLatch.Q ;
	assign \mchip.s444.d_flip_flops.shift_out  = \mchip.s444.d_flip_flops.dff_reg.myLatch.Q [3];
	assign \mchip.s444.d_flip_flops.sum_out  = \mchip.s444.carry_logic.sum_out ;
	assign \mchip.s444.dff0_out  = \mchip.s444.d_flip_flops.dff.Q [0];
	assign \mchip.s444.dff1_out  = \mchip.s444.d_flip_flops.dff.Q [1];
	assign \mchip.s444.en  = io_in[11];
	assign \mchip.s444.feed0  = io_in[3:0];
	assign \mchip.s444.feed0_out  = \mchip.s444.d_flip_flops.feed0_out ;
	assign \mchip.s444.feed1  = {io_in[4], io_in[2:0]};
	assign \mchip.s444.feed1_out  = \mchip.s444.carry_logic.prop ;
	assign \mchip.s444.lut1  = \mchip.s444.carry_logic.prop ;
	assign \mchip.s444.lut2  = \mchip.s444.carry_logic.gen ;
	assign \mchip.s444.lut5_mux.clk  = io_in[12];
	assign \mchip.s444.lut5_mux.en  = io_in[11];
	assign \mchip.s444.lut5_mux.feed0_out  = \mchip.s444.d_flip_flops.feed0_out ;
	assign \mchip.s444.lut5_mux.feed1_3  = io_in[4];
	assign \mchip.s444.lut5_mux.lut1  = \mchip.s444.carry_logic.prop ;
	assign \mchip.s444.lut5_mux.lut5_reg.I  = \mchip.s444.s444_logic.l2_reg.myLatch.Q [15];
	assign \mchip.s444.lut5_mux.lut5_reg.O  = \mchip.s444.lut5_mux.lut5_reg.myLatch.Q ;
	assign \mchip.s444.lut5_mux.lut5_reg.Q  = \mchip.s444.lut5_mux.lut5_reg.myLatch.Q ;
	assign \mchip.s444.lut5_mux.lut5_reg.clock  = io_in[12];
	assign \mchip.s444.lut5_mux.lut5_reg.en  = 1'h1;
	assign \mchip.s444.lut5_mux.lut5_reg.highBit  = \mchip.s444.lut5_mux.lut5_reg.myLatch.Q ;
	assign \mchip.s444.lut5_mux.lut5_reg.left  = 1'h1;
	assign \mchip.s444.lut5_mux.lut5_reg.lowBit  = \mchip.s444.lut5_mux.lut5_reg.myLatch.Q ;
	assign \mchip.s444.lut5_mux.lut5_reg.myLatch.D  = \mchip.s444.s444_logic.l2_reg.myLatch.Q [15];
	assign \mchip.s444.lut5_mux.lut5_reg.myLatch.clear  = io_in[13];
	assign \mchip.s444.lut5_mux.lut5_reg.myLatch.clock  = io_in[12];
	assign \mchip.s444.lut5_mux.lut5_reg.myLatch.en  = 1'h1;
	assign \mchip.s444.lut5_mux.lut5_reg.myLatch.load  = io_in[11];
	assign \mchip.s444.lut5_mux.lut5_reg.reset  = io_in[13];
	assign \mchip.s444.lut5_mux.lut5_reg.shift  = io_in[11];
	assign \mchip.s444.lut5_mux.lut5_reg.shiftResult  = \mchip.s444.s444_logic.l2_reg.myLatch.Q [15];
	assign \mchip.s444.lut5_mux.lut5_reg.shiftedLeft  = \mchip.s444.s444_logic.l2_reg.myLatch.Q [15];
	assign \mchip.s444.lut5_mux.lut5_reg.shiftedRight  = \mchip.s444.s444_logic.l2_reg.myLatch.Q [15];
	assign \mchip.s444.lut5_mux.lut5_sel  = \mchip.s444.lut5_mux.lut5_reg.myLatch.Q ;
	assign \mchip.s444.lut5_mux.reset  = io_in[13];
	assign \mchip.s444.lut5_mux.shift_in  = \mchip.s444.s444_logic.l2_reg.myLatch.Q [15];
	assign \mchip.s444.lut5_mux.shift_out  = \mchip.s444.lut5_mux.lut5_reg.myLatch.Q ;
	assign \mchip.s444.main  = io_in[8:5];
	assign \mchip.s444.main_out  = \mchip.s444.carry_logic.gen ;
	assign \mchip.s444.reset  = io_in[13];
	assign \mchip.s444.s444_logic.clk  = io_in[12];
	assign \mchip.s444.s444_logic.en  = io_in[11];
	assign \mchip.s444.s444_logic.feed0  = io_in[3:0];
	assign \mchip.s444.s444_logic.feed1  = {io_in[4], io_in[2:0]};
	assign \mchip.s444.s444_logic.feed2  = {2'h0, io_in[6:5]};
	assign \mchip.s444.s444_logic.l0.D  = \mchip.s444.s444_logic.l0_reg.myLatch.Q ;
	assign \mchip.s444.s444_logic.l0.I  = io_in[3:0];
	assign \mchip.s444.s444_logic.l0_dat  = \mchip.s444.s444_logic.l0_reg.myLatch.Q ;
	assign \mchip.s444.s444_logic.l0_reg.I  = \mchip.s444.s444_logic.m2_reg.myLatch.Q ;
	assign \mchip.s444.s444_logic.l0_reg.O  = \mchip.s444.s444_logic.l0_reg.myLatch.Q [15];
	assign \mchip.s444.s444_logic.l0_reg.Q  = \mchip.s444.s444_logic.l0_reg.myLatch.Q ;
	assign \mchip.s444.s444_logic.l0_reg.clock  = io_in[12];
	assign \mchip.s444.s444_logic.l0_reg.en  = 1'h1;
	assign \mchip.s444.s444_logic.l0_reg.highBit  = \mchip.s444.s444_logic.l0_reg.myLatch.Q [15];
	assign \mchip.s444.s444_logic.l0_reg.left  = 1'h1;
	assign \mchip.s444.s444_logic.l0_reg.lowBit  = \mchip.s444.s444_logic.l0_reg.myLatch.Q [0];
	assign \mchip.s444.s444_logic.l0_reg.myLatch.D  = {\mchip.s444.s444_logic.l0_reg.myLatch.Q [14:0], \mchip.s444.s444_logic.m2_reg.myLatch.Q };
	assign \mchip.s444.s444_logic.l0_reg.myLatch.clear  = io_in[13];
	assign \mchip.s444.s444_logic.l0_reg.myLatch.clock  = io_in[12];
	assign \mchip.s444.s444_logic.l0_reg.myLatch.en  = 1'h1;
	assign \mchip.s444.s444_logic.l0_reg.myLatch.load  = io_in[11];
	assign \mchip.s444.s444_logic.l0_reg.reset  = io_in[13];
	assign \mchip.s444.s444_logic.l0_reg.shift  = io_in[11];
	assign \mchip.s444.s444_logic.l0_reg.shiftResult  = {\mchip.s444.s444_logic.l0_reg.myLatch.Q [14:0], \mchip.s444.s444_logic.m2_reg.myLatch.Q };
	assign \mchip.s444.s444_logic.l0_reg.shiftedLeft  = {\mchip.s444.s444_logic.l0_reg.myLatch.Q [14:0], \mchip.s444.s444_logic.m2_reg.myLatch.Q };
	assign \mchip.s444.s444_logic.l1.D  = \mchip.s444.s444_logic.l1_reg.myLatch.Q ;
	assign \mchip.s444.s444_logic.l1.I  = {1'h0, io_in[2:0]};
	assign \mchip.s444.s444_logic.l1.O  = \mchip.s444.carry_logic.prop ;
	assign \mchip.s444.s444_logic.l1_dat  = \mchip.s444.s444_logic.l1_reg.myLatch.Q ;
	assign \mchip.s444.s444_logic.l1_reg.I  = \mchip.s444.s444_logic.l0_reg.myLatch.Q [15];
	assign \mchip.s444.s444_logic.l1_reg.O  = \mchip.s444.s444_logic.l1_reg.myLatch.Q [15];
	assign \mchip.s444.s444_logic.l1_reg.Q  = \mchip.s444.s444_logic.l1_reg.myLatch.Q ;
	assign \mchip.s444.s444_logic.l1_reg.clock  = io_in[12];
	assign \mchip.s444.s444_logic.l1_reg.en  = 1'h1;
	assign \mchip.s444.s444_logic.l1_reg.highBit  = \mchip.s444.s444_logic.l1_reg.myLatch.Q [15];
	assign \mchip.s444.s444_logic.l1_reg.left  = 1'h1;
	assign \mchip.s444.s444_logic.l1_reg.lowBit  = \mchip.s444.s444_logic.l1_reg.myLatch.Q [0];
	assign \mchip.s444.s444_logic.l1_reg.myLatch.D  = {\mchip.s444.s444_logic.l1_reg.myLatch.Q [14:0], \mchip.s444.s444_logic.l0_reg.myLatch.Q [15]};
	assign \mchip.s444.s444_logic.l1_reg.myLatch.clear  = io_in[13];
	assign \mchip.s444.s444_logic.l1_reg.myLatch.clock  = io_in[12];
	assign \mchip.s444.s444_logic.l1_reg.myLatch.en  = 1'h1;
	assign \mchip.s444.s444_logic.l1_reg.myLatch.load  = io_in[11];
	assign \mchip.s444.s444_logic.l1_reg.reset  = io_in[13];
	assign \mchip.s444.s444_logic.l1_reg.shift  = io_in[11];
	assign \mchip.s444.s444_logic.l1_reg.shiftResult  = {\mchip.s444.s444_logic.l1_reg.myLatch.Q [14:0], \mchip.s444.s444_logic.l0_reg.myLatch.Q [15]};
	assign \mchip.s444.s444_logic.l1_reg.shiftedLeft  = {\mchip.s444.s444_logic.l1_reg.myLatch.Q [14:0], \mchip.s444.s444_logic.l0_reg.myLatch.Q [15]};
	assign \mchip.s444.s444_logic.l2.D  = \mchip.s444.s444_logic.l2_reg.myLatch.Q ;
	assign \mchip.s444.s444_logic.l2.I  = {2'h0, io_in[6:5]};
	assign \mchip.s444.s444_logic.l2.O  = \mchip.s444.carry_logic.gen ;
	assign \mchip.s444.s444_logic.l2_dat  = \mchip.s444.s444_logic.l2_reg.myLatch.Q ;
	assign \mchip.s444.s444_logic.l2_reg.I  = \mchip.s444.s444_logic.l1_reg.myLatch.Q [15];
	assign \mchip.s444.s444_logic.l2_reg.O  = \mchip.s444.s444_logic.l2_reg.myLatch.Q [15];
	assign \mchip.s444.s444_logic.l2_reg.Q  = \mchip.s444.s444_logic.l2_reg.myLatch.Q ;
	assign \mchip.s444.s444_logic.l2_reg.clock  = io_in[12];
	assign \mchip.s444.s444_logic.l2_reg.en  = 1'h1;
	assign \mchip.s444.s444_logic.l2_reg.highBit  = \mchip.s444.s444_logic.l2_reg.myLatch.Q [15];
	assign \mchip.s444.s444_logic.l2_reg.left  = 1'h1;
	assign \mchip.s444.s444_logic.l2_reg.lowBit  = \mchip.s444.s444_logic.l2_reg.myLatch.Q [0];
	assign \mchip.s444.s444_logic.l2_reg.myLatch.D  = {\mchip.s444.s444_logic.l2_reg.myLatch.Q [14:0], \mchip.s444.s444_logic.l1_reg.myLatch.Q [15]};
	assign \mchip.s444.s444_logic.l2_reg.myLatch.clear  = io_in[13];
	assign \mchip.s444.s444_logic.l2_reg.myLatch.clock  = io_in[12];
	assign \mchip.s444.s444_logic.l2_reg.myLatch.en  = 1'h1;
	assign \mchip.s444.s444_logic.l2_reg.myLatch.load  = io_in[11];
	assign \mchip.s444.s444_logic.l2_reg.reset  = io_in[13];
	assign \mchip.s444.s444_logic.l2_reg.shift  = io_in[11];
	assign \mchip.s444.s444_logic.l2_reg.shiftResult  = {\mchip.s444.s444_logic.l2_reg.myLatch.Q [14:0], \mchip.s444.s444_logic.l1_reg.myLatch.Q [15]};
	assign \mchip.s444.s444_logic.l2_reg.shiftedLeft  = {\mchip.s444.s444_logic.l2_reg.myLatch.Q [14:0], \mchip.s444.s444_logic.l1_reg.myLatch.Q [15]};
	assign \mchip.s444.s444_logic.lut1  = \mchip.s444.carry_logic.prop ;
	assign \mchip.s444.s444_logic.lut2  = \mchip.s444.carry_logic.gen ;
	assign \mchip.s444.s444_logic.m0_reg.I  = io_in[10];
	assign \mchip.s444.s444_logic.m0_reg.O  = \mchip.s444.s444_logic.m0_reg.myLatch.Q ;
	assign \mchip.s444.s444_logic.m0_reg.Q  = \mchip.s444.s444_logic.m0_reg.myLatch.Q ;
	assign \mchip.s444.s444_logic.m0_reg.clock  = io_in[12];
	assign \mchip.s444.s444_logic.m0_reg.en  = 1'h1;
	assign \mchip.s444.s444_logic.m0_reg.highBit  = \mchip.s444.s444_logic.m0_reg.myLatch.Q ;
	assign \mchip.s444.s444_logic.m0_reg.left  = 1'h1;
	assign \mchip.s444.s444_logic.m0_reg.lowBit  = \mchip.s444.s444_logic.m0_reg.myLatch.Q ;
	assign \mchip.s444.s444_logic.m0_reg.myLatch.D  = io_in[10];
	assign \mchip.s444.s444_logic.m0_reg.myLatch.clear  = io_in[13];
	assign \mchip.s444.s444_logic.m0_reg.myLatch.clock  = io_in[12];
	assign \mchip.s444.s444_logic.m0_reg.myLatch.en  = 1'h1;
	assign \mchip.s444.s444_logic.m0_reg.myLatch.load  = io_in[11];
	assign \mchip.s444.s444_logic.m0_reg.reset  = io_in[13];
	assign \mchip.s444.s444_logic.m0_reg.shift  = io_in[11];
	assign \mchip.s444.s444_logic.m0_reg.shiftResult  = io_in[10];
	assign \mchip.s444.s444_logic.m0_reg.shiftedLeft  = io_in[10];
	assign \mchip.s444.s444_logic.m0_reg.shiftedRight  = io_in[10];
	assign \mchip.s444.s444_logic.m0_sel  = \mchip.s444.s444_logic.m0_reg.myLatch.Q ;
	assign \mchip.s444.s444_logic.m1_reg.I  = \mchip.s444.s444_logic.m0_reg.myLatch.Q ;
	assign \mchip.s444.s444_logic.m1_reg.O  = \mchip.s444.s444_logic.m1_reg.myLatch.Q ;
	assign \mchip.s444.s444_logic.m1_reg.Q  = \mchip.s444.s444_logic.m1_reg.myLatch.Q ;
	assign \mchip.s444.s444_logic.m1_reg.clock  = io_in[12];
	assign \mchip.s444.s444_logic.m1_reg.en  = 1'h1;
	assign \mchip.s444.s444_logic.m1_reg.highBit  = \mchip.s444.s444_logic.m1_reg.myLatch.Q ;
	assign \mchip.s444.s444_logic.m1_reg.left  = 1'h1;
	assign \mchip.s444.s444_logic.m1_reg.lowBit  = \mchip.s444.s444_logic.m1_reg.myLatch.Q ;
	assign \mchip.s444.s444_logic.m1_reg.myLatch.D  = \mchip.s444.s444_logic.m0_reg.myLatch.Q ;
	assign \mchip.s444.s444_logic.m1_reg.myLatch.clear  = io_in[13];
	assign \mchip.s444.s444_logic.m1_reg.myLatch.clock  = io_in[12];
	assign \mchip.s444.s444_logic.m1_reg.myLatch.en  = 1'h1;
	assign \mchip.s444.s444_logic.m1_reg.myLatch.load  = io_in[11];
	assign \mchip.s444.s444_logic.m1_reg.reset  = io_in[13];
	assign \mchip.s444.s444_logic.m1_reg.shift  = io_in[11];
	assign \mchip.s444.s444_logic.m1_reg.shiftResult  = \mchip.s444.s444_logic.m0_reg.myLatch.Q ;
	assign \mchip.s444.s444_logic.m1_reg.shiftedLeft  = \mchip.s444.s444_logic.m0_reg.myLatch.Q ;
	assign \mchip.s444.s444_logic.m1_reg.shiftedRight  = \mchip.s444.s444_logic.m0_reg.myLatch.Q ;
	assign \mchip.s444.s444_logic.m1_sel  = \mchip.s444.s444_logic.m1_reg.myLatch.Q ;
	assign \mchip.s444.s444_logic.m2_reg.I  = \mchip.s444.s444_logic.m1_reg.myLatch.Q ;
	assign \mchip.s444.s444_logic.m2_reg.O  = \mchip.s444.s444_logic.m2_reg.myLatch.Q ;
	assign \mchip.s444.s444_logic.m2_reg.Q  = \mchip.s444.s444_logic.m2_reg.myLatch.Q ;
	assign \mchip.s444.s444_logic.m2_reg.clock  = io_in[12];
	assign \mchip.s444.s444_logic.m2_reg.en  = 1'h1;
	assign \mchip.s444.s444_logic.m2_reg.highBit  = \mchip.s444.s444_logic.m2_reg.myLatch.Q ;
	assign \mchip.s444.s444_logic.m2_reg.left  = 1'h1;
	assign \mchip.s444.s444_logic.m2_reg.lowBit  = \mchip.s444.s444_logic.m2_reg.myLatch.Q ;
	assign \mchip.s444.s444_logic.m2_reg.myLatch.D  = \mchip.s444.s444_logic.m1_reg.myLatch.Q ;
	assign \mchip.s444.s444_logic.m2_reg.myLatch.clear  = io_in[13];
	assign \mchip.s444.s444_logic.m2_reg.myLatch.clock  = io_in[12];
	assign \mchip.s444.s444_logic.m2_reg.myLatch.en  = 1'h1;
	assign \mchip.s444.s444_logic.m2_reg.myLatch.load  = io_in[11];
	assign \mchip.s444.s444_logic.m2_reg.reset  = io_in[13];
	assign \mchip.s444.s444_logic.m2_reg.shift  = io_in[11];
	assign \mchip.s444.s444_logic.m2_reg.shiftResult  = \mchip.s444.s444_logic.m1_reg.myLatch.Q ;
	assign \mchip.s444.s444_logic.m2_reg.shiftedLeft  = \mchip.s444.s444_logic.m1_reg.myLatch.Q ;
	assign \mchip.s444.s444_logic.m2_reg.shiftedRight  = \mchip.s444.s444_logic.m1_reg.myLatch.Q ;
	assign \mchip.s444.s444_logic.m2_sel  = \mchip.s444.s444_logic.m2_reg.myLatch.Q ;
	assign \mchip.s444.s444_logic.main  = io_in[8:5];
	assign \mchip.s444.s444_logic.reset  = io_in[13];
	assign \mchip.s444.s444_logic.shift_in  = io_in[10];
	assign \mchip.s444.s444_logic.shift_l0  = \mchip.s444.s444_logic.l0_reg.myLatch.Q [15];
	assign \mchip.s444.s444_logic.shift_l1  = \mchip.s444.s444_logic.l1_reg.myLatch.Q [15];
	assign \mchip.s444.s444_logic.shift_l2  = \mchip.s444.s444_logic.l2_reg.myLatch.Q [15];
	assign \mchip.s444.s444_logic.shift_m0  = \mchip.s444.s444_logic.m0_reg.myLatch.Q ;
	assign \mchip.s444.s444_logic.shift_m1  = \mchip.s444.s444_logic.m1_reg.myLatch.Q ;
	assign \mchip.s444.s444_logic.shift_m2  = \mchip.s444.s444_logic.m2_reg.myLatch.Q ;
	assign \mchip.s444.s444_logic.shift_out  = \mchip.s444.s444_logic.l2_reg.myLatch.Q [15];
	assign \mchip.s444.shift0  = \mchip.s444.s444_logic.l2_reg.myLatch.Q [15];
	assign \mchip.s444.shift1  = \mchip.s444.lut5_mux.lut5_reg.myLatch.Q ;
	assign \mchip.s444.shift_in  = io_in[10];
	assign \mchip.s444.shift_out  = \mchip.s444.d_flip_flops.dff_reg.myLatch.Q [3];
	assign \mchip.s444.sum_out  = \mchip.s444.carry_logic.sum_out ;
endmodule
module d14_jessief_trafficlight (
	io_in,
	io_out
);
	wire [10:0] _000_;
	wire _001_;
	wire _002_;
	wire _003_;
	wire _004_;
	wire _005_;
	wire _006_;
	wire _007_;
	wire _008_;
	wire _009_;
	wire _010_;
	wire _011_;
	wire _012_;
	wire _013_;
	wire _014_;
	wire _015_;
	wire _016_;
	wire _017_;
	wire _018_;
	wire _019_;
	wire _020_;
	wire _021_;
	wire _022_;
	wire _023_;
	wire _024_;
	wire _025_;
	wire _026_;
	wire _027_;
	wire _028_;
	wire _029_;
	wire _030_;
	wire _031_;
	wire _032_;
	wire _033_;
	wire _034_;
	wire _035_;
	wire _036_;
	wire _037_;
	wire _038_;
	wire _039_;
	wire _040_;
	wire _041_;
	wire _042_;
	wire _043_;
	wire _044_;
	wire _045_;
	wire _046_;
	wire _047_;
	wire _048_;
	wire _049_;
	wire _050_;
	wire _051_;
	wire _052_;
	wire _053_;
	wire _054_;
	wire _055_;
	wire _056_;
	wire _057_;
	wire _058_;
	wire _059_;
	wire _060_;
	wire _061_;
	wire _062_;
	wire _063_;
	wire _064_;
	wire _065_;
	wire _066_;
	wire _067_;
	wire _068_;
	wire _069_;
	wire _070_;
	wire _071_;
	wire _072_;
	wire _073_;
	wire _074_;
	wire _075_;
	wire _076_;
	wire _077_;
	wire _078_;
	wire _079_;
	wire _080_;
	wire _081_;
	wire _082_;
	wire _083_;
	wire _084_;
	wire _085_;
	wire _086_;
	wire _087_;
	wire _088_;
	wire _089_;
	wire _090_;
	wire _091_;
	wire _092_;
	wire _093_;
	wire _094_;
	wire _095_;
	wire _096_;
	wire _097_;
	wire _098_;
	wire _099_;
	wire _100_;
	wire _101_;
	wire _102_;
	wire _103_;
	wire _104_;
	wire _105_;
	wire _106_;
	wire _107_;
	wire _108_;
	wire _109_;
	wire _110_;
	wire _111_;
	wire _112_;
	wire _113_;
	wire _114_;
	wire _115_;
	wire _116_;
	wire _117_;
	wire _118_;
	wire _119_;
	wire _120_;
	wire _121_;
	wire _122_;
	wire _123_;
	wire _124_;
	wire _125_;
	wire _126_;
	wire _127_;
	wire _128_;
	wire _129_;
	wire _130_;
	wire _131_;
	wire _132_;
	wire _133_;
	wire _134_;
	wire _135_;
	wire _136_;
	wire _137_;
	wire [7:0] _138_;
	wire [7:0] _139_;
	wire [7:0] _140_;
	input wire [13:0] io_in;
	output wire [13:0] io_out;
	wire \mchip.button ;
	wire \mchip.car1 ;
	wire \mchip.car2 ;
	wire \mchip.car3 ;
	wire \mchip.car4 ;
	wire \mchip.clock ;
	wire \mchip.control.car1 ;
	wire \mchip.control.car2 ;
	wire \mchip.control.car3 ;
	wire \mchip.control.car4 ;
	wire \mchip.control.clock ;
	reg \mchip.control.five_clr ;
	reg \mchip.control.five_en ;
	wire \mchip.control.green1 ;
	wire \mchip.control.green2 ;
	wire \mchip.control.green3 ;
	wire [3:0] \mchip.control.nextState ;
	wire \mchip.control.orange ;
	wire \mchip.control.ped ;
	reg \mchip.control.ped_clr ;
	wire \mchip.control.red1 ;
	wire \mchip.control.red2 ;
	wire \mchip.control.red3 ;
	wire \mchip.control.reset ;
	reg [3:0] \mchip.control.state ;
	reg \mchip.control.stop_clr ;
	reg \mchip.control.stop_en ;
	wire \mchip.control.stop_five ;
	wire \mchip.control.stop_ped ;
	wire \mchip.control.stop_yellow ;
	wire \mchip.control.turn ;
	wire \mchip.control.white ;
	wire \mchip.control.yellow1 ;
	wire \mchip.control.yellow2 ;
	wire \mchip.control.yellow3 ;
	reg \mchip.control.yellow_clr ;
	reg \mchip.control.yellow_en ;
	wire [7:0] \mchip.five.D ;
	wire [7:0] \mchip.five.Q ;
	wire \mchip.five.clear ;
	wire \mchip.five.clock ;
	wire \mchip.five.en ;
	wire \mchip.five.load ;
	wire \mchip.five_clr ;
	wire \mchip.five_en ;
	wire \mchip.green1 ;
	wire \mchip.green2 ;
	wire \mchip.green3 ;
	wire [11:0] \mchip.io_in ;
	wire [11:0] \mchip.io_out ;
	wire \mchip.orange ;
	wire \mchip.ped ;
	wire \mchip.ped_clr ;
	wire \mchip.pedestrian.button ;
	wire \mchip.pedestrian.clock ;
	reg \mchip.pedestrian.ped ;
	wire \mchip.pedestrian.ped_clr ;
	wire \mchip.red1 ;
	wire \mchip.red2 ;
	wire \mchip.red3 ;
	wire \mchip.reset ;
	wire [7:0] \mchip.stop.D ;
	wire [7:0] \mchip.stop.Q ;
	wire \mchip.stop.clear ;
	wire \mchip.stop.clock ;
	wire \mchip.stop.en ;
	wire \mchip.stop.load ;
	wire \mchip.stop_clr ;
	wire \mchip.stop_en ;
	wire \mchip.stop_five ;
	wire \mchip.stop_ped ;
	wire \mchip.stop_yellow ;
	wire \mchip.turn ;
	wire \mchip.white ;
	wire [7:0] \mchip.yellow.D ;
	wire [7:0] \mchip.yellow.Q ;
	wire \mchip.yellow.clear ;
	wire \mchip.yellow.clock ;
	wire \mchip.yellow.en ;
	wire \mchip.yellow.load ;
	wire \mchip.yellow1 ;
	wire \mchip.yellow2 ;
	wire \mchip.yellow3 ;
	wire \mchip.yellow_clr ;
	wire \mchip.yellow_en ;
	assign _138_[0] = ~\mchip.five.Q [0];
	assign _139_[0] = ~\mchip.stop.Q [0];
	assign _083_ = \mchip.control.state [3] & ~\mchip.control.state [2];
	assign _084_ = \mchip.control.state [1] | \mchip.control.state [0];
	assign _085_ = _083_ & ~_084_;
	assign _086_ = \mchip.control.state [2] & ~\mchip.control.state [3];
	assign _087_ = \mchip.control.state [1] & \mchip.control.state [0];
	assign _088_ = _087_ & _086_;
	assign _089_ = ~(_088_ | _085_);
	assign _090_ = \mchip.control.state [1] | ~\mchip.control.state [0];
	assign _091_ = _086_ & ~_090_;
	assign _092_ = \mchip.control.state [0] | ~\mchip.control.state [1];
	assign _093_ = _086_ & ~_092_;
	assign _094_ = _093_ | _091_;
	assign _095_ = _089_ & ~_094_;
	assign _096_ = \mchip.control.state [3] | \mchip.control.state [2];
	assign _097_ = ~(_096_ | _090_);
	assign _098_ = _096_ | _092_;
	assign _099_ = _097_ | ~_098_;
	assign _100_ = _087_ & ~_096_;
	assign _101_ = _086_ & ~_084_;
	assign _102_ = _101_ | _100_;
	assign _103_ = _102_ | _099_;
	assign _104_ = _095_ & ~_103_;
	assign _105_ = ~(_101_ & \mchip.stop.Q [0]);
	assign _106_ = _085_ & ~\mchip.five.Q [0];
	assign _107_ = _105_ & ~_106_;
	assign \mchip.control.nextState [3] = ~(_107_ | _104_);
	assign _000_[10] = \mchip.control.nextState [3] & ~io_in[13];
	assign _140_[0] = ~\mchip.yellow.Q [0];
	assign _108_ = ~io_in[4];
	assign _109_ = ~io_in[3];
	assign _110_ = _109_ & ~_098_;
	assign _111_ = io_in[2] | io_in[1];
	assign _112_ = _100_ & ~_111_;
	assign _113_ = _112_ | _110_;
	assign _114_ = _098_ & ~_100_;
	assign _115_ = (_114_ ? _108_ : _113_);
	assign _116_ = _139_[0] & ~_115_;
	assign _117_ = _116_ | ~_097_;
	assign _118_ = ~(_116_ | _098_);
	assign _119_ = _117_ & ~_118_;
	assign _120_ = _100_ & ~_116_;
	assign _121_ = _101_ & ~\mchip.stop.Q [0];
	assign _122_ = _121_ | _120_;
	assign _123_ = _119_ & ~_122_;
	assign _124_ = _109_ & ~_111_;
	assign _125_ = _124_ & ~io_in[4];
	assign _126_ = ~(_125_ & \mchip.five.Q [0]);
	assign _127_ = _085_ & ~_126_;
	assign _128_ = _125_ | \mchip.pedestrian.ped ;
	assign _129_ = \mchip.yellow.Q [0] & ~_128_;
	assign _130_ = _088_ & ~_129_;
	assign _131_ = _130_ | _127_;
	assign _132_ = io_in[4] & ~\mchip.pedestrian.ped ;
	assign _133_ = ~(_132_ | _111_);
	assign _134_ = _133_ & ~io_in[3];
	assign _135_ = \mchip.yellow.Q [0] & ~_134_;
	assign _136_ = _091_ & ~_135_;
	assign _137_ = ~(io_in[2] | io_in[1]);
	assign _019_ = ~\mchip.pedestrian.ped ;
	assign _020_ = ~(io_in[4] | io_in[3]);
	assign _021_ = _019_ & ~_020_;
	assign _022_ = _137_ & ~_021_;
	assign _023_ = \mchip.yellow.Q [0] & ~_022_;
	assign _024_ = _093_ & ~_023_;
	assign _025_ = _024_ | _136_;
	assign _026_ = _025_ | _131_;
	assign _027_ = _026_ | ~_123_;
	assign _028_ = _111_ | _019_;
	assign _029_ = _028_ | io_in[3];
	assign _030_ = _108_ & ~_029_;
	assign \mchip.control.nextState [2] = (_104_ ? _030_ : _027_);
	assign _031_ = \mchip.control.nextState [2] & ~io_in[13];
	assign _032_ = ~io_in[13];
	assign _033_ = _124_ | io_in[4];
	assign _034_ = _033_ | _138_[0];
	assign _035_ = _085_ & ~_034_;
	assign _036_ = _019_ & ~_033_;
	assign _037_ = \mchip.yellow.Q [0] & ~_036_;
	assign _038_ = _088_ & ~_037_;
	assign _039_ = _038_ | _035_;
	assign _040_ = _124_ | _140_[0];
	assign _041_ = _091_ & ~_040_;
	assign _042_ = io_in[4] | ~io_in[3];
	assign _043_ = _019_ & ~_042_;
	assign _044_ = _043_ | _111_;
	assign _045_ = \mchip.yellow.Q [0] & ~_044_;
	assign _046_ = _093_ & ~_045_;
	assign _047_ = _046_ | _041_;
	assign _048_ = _047_ | _039_;
	assign _049_ = _114_ & ~_048_;
	assign _050_ = (_104_ ? _033_ : _049_);
	assign _051_ = _032_ & ~_050_;
	assign _052_ = _051_ | _031_;
	assign _004_ = _052_ | _000_[10];
	assign _053_ = _051_ | _000_[10];
	assign _003_ = _053_ | ~_031_;
	assign _006_ = _031_ | _000_[10];
	assign _007_ = _050_ | io_in[13];
	assign _002_ = _006_ | _007_;
	assign _005_ = _000_[10] | ~_031_;
	assign _001_ = _005_ | _007_;
	assign _054_ = _109_ & ~_137_;
	assign _055_ = _108_ & ~_054_;
	assign _056_ = _055_ | _138_[0];
	assign _057_ = _056_ | ~_085_;
	assign _058_ = _019_ & ~_055_;
	assign _059_ = \mchip.yellow.Q [0] & ~_058_;
	assign _060_ = _088_ & ~_059_;
	assign _061_ = _057_ & ~_060_;
	assign _062_ = _109_ & ~_133_;
	assign _063_ = \mchip.yellow.Q [0] & ~_062_;
	assign _064_ = _091_ & ~_063_;
	assign _065_ = _133_ | _140_[0];
	assign _066_ = _093_ & ~_065_;
	assign _067_ = _066_ | _064_;
	assign _068_ = _061_ & ~_067_;
	assign _069_ = _100_ | _097_;
	assign _070_ = _068_ & ~_069_;
	assign _071_ = (_104_ ? _055_ : _070_);
	assign \mchip.control.nextState [0] = ~_071_;
	assign \mchip.control.nextState [1] = ~_050_;
	assign _008_ = _032_ & ~_071_;
	assign _017_ = _008_ | _051_;
	assign _016_ = _007_ & ~_008_;
	assign _015_ = _017_ ^ _031_;
	assign _018_ = ~_008_;
	assign _072_ = _031_ & ~_017_;
	assign _073_ = _008_ & ~_051_;
	assign _074_ = ~(_073_ | _031_);
	assign _009_ = _074_ | _072_;
	assign _010_ = _016_ ^ _031_;
	assign _075_ = _031_ & ~_073_;
	assign _011_ = _075_ | _074_;
	assign _076_ = _051_ & ~_008_;
	assign _077_ = _031_ & ~_076_;
	assign _078_ = ~(_076_ | _031_);
	assign _012_ = _078_ | _077_;
	assign _079_ = _017_ & ~_076_;
	assign _080_ = _031_ & ~_079_;
	assign _081_ = ~(_079_ | _031_);
	assign _013_ = _081_ | _080_;
	assign _082_ = _016_ & ~_031_;
	assign _014_ = _082_ | _072_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.control.state [0] <= 1'h0;
		else
			\mchip.control.state [0] <= \mchip.control.nextState [0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.control.state [1] <= 1'h0;
		else
			\mchip.control.state [1] <= \mchip.control.nextState [1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.control.state [2] <= 1'h0;
		else
			\mchip.control.state [2] <= \mchip.control.nextState [2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.control.state [3] <= 1'h0;
		else
			\mchip.control.state [3] <= \mchip.control.nextState [3];
	reg \io_out_reg[3] ;
	always @(posedge io_in[12])
		if (_006_)
			\io_out_reg[3]  <= 1'h0;
		else
			\io_out_reg[3]  <= _008_;
	assign io_out[3] = \io_out_reg[3] ;
	always @(posedge io_in[12])
		if (_006_)
			\mchip.control.five_clr  <= 1'h0;
		else
			\mchip.control.five_clr  <= _007_;
	reg \io_out_reg[7] ;
	always @(posedge io_in[12])
		if (_001_)
			\io_out_reg[7]  <= 1'h0;
		else
			\io_out_reg[7]  <= _018_;
	assign io_out[7] = \io_out_reg[7] ;
	always @(posedge io_in[12]) \mchip.control.five_en  <= _000_[10];
	reg \io_out_reg[4] ;
	always @(posedge io_in[12])
		if (_005_)
			\io_out_reg[4]  <= 1'h0;
		else
			\io_out_reg[4]  <= _008_;
	assign io_out[4] = \io_out_reg[4] ;
	reg \io_out_reg[0] ;
	always @(posedge io_in[12])
		if (_005_)
			\io_out_reg[0]  <= 1'h0;
		else
			\io_out_reg[0]  <= _016_;
	assign io_out[0] = \io_out_reg[0] ;
	always @(posedge io_in[12])
		if (_005_)
			\mchip.control.yellow_en  <= 1'h0;
		else
			\mchip.control.yellow_en  <= _017_;
	reg \io_out_reg[1] ;
	always @(posedge io_in[12])
		if (_005_)
			\io_out_reg[1]  <= 1'h1;
		else
			\io_out_reg[1]  <= _017_;
	assign io_out[1] = \io_out_reg[1] ;
	reg \io_out_reg[9] ;
	always @(posedge io_in[12])
		if (_004_)
			\io_out_reg[9]  <= 1'h0;
		else
			\io_out_reg[9]  <= _008_;
	assign io_out[9] = \io_out_reg[9] ;
	always @(posedge io_in[12])
		if (_000_[10])
			\mchip.control.stop_en  <= 1'h0;
		else
			\mchip.control.stop_en  <= _015_;
	always @(posedge io_in[12])
		if (_000_[10])
			\mchip.control.yellow_clr  <= 1'h0;
		else
			\mchip.control.yellow_clr  <= _009_;
	always @(posedge io_in[12])
		if (_000_[10])
			\mchip.control.stop_clr  <= 1'h1;
		else
			\mchip.control.stop_clr  <= _010_;
	reg \io_out_reg[11] ;
	always @(posedge io_in[12])
		if (_000_[10])
			\io_out_reg[11]  <= 1'h1;
		else
			\io_out_reg[11]  <= _011_;
	assign io_out[11] = \io_out_reg[11] ;
	reg \io_out_reg[8] ;
	always @(posedge io_in[12])
		if (_000_[10])
			\io_out_reg[8]  <= 1'h1;
		else
			\io_out_reg[8]  <= _012_;
	assign io_out[8] = \io_out_reg[8] ;
	reg \io_out_reg[5] ;
	always @(posedge io_in[12])
		if (_000_[10])
			\io_out_reg[5]  <= 1'h1;
		else
			\io_out_reg[5]  <= _013_;
	assign io_out[5] = \io_out_reg[5] ;
	always @(posedge io_in[12])
		if (_000_[10])
			\mchip.control.ped_clr  <= 1'h0;
		else
			\mchip.control.ped_clr  <= _014_;
	reg \io_out_reg[10] ;
	always @(posedge io_in[12])
		if (_003_)
			\io_out_reg[10]  <= 1'h0;
		else
			\io_out_reg[10]  <= _008_;
	assign io_out[10] = \io_out_reg[10] ;
	reg \io_out_reg[6] ;
	always @(posedge io_in[12])
		if (_002_)
			\io_out_reg[6]  <= 1'h0;
		else
			\io_out_reg[6]  <= _018_;
	assign io_out[6] = \io_out_reg[6] ;
	reg \io_out_reg[2] ;
	always @(posedge io_in[12])
		if (_002_)
			\io_out_reg[2]  <= 1'h0;
		else
			\io_out_reg[2]  <= _008_;
	assign io_out[2] = \io_out_reg[2] ;
	always @(posedge io_in[12])
		if (io_in[0])
			\mchip.pedestrian.ped  <= 1'h1;
		else if (\mchip.control.ped_clr )
			\mchip.pedestrian.ped  <= 1'h0;
	reg \mchip.five.Q_reg[0] ;
	always @(posedge io_in[12])
		if (\mchip.control.five_clr )
			\mchip.five.Q_reg[0]  <= 1'h0;
		else if (\mchip.control.five_en )
			\mchip.five.Q_reg[0]  <= _138_[0];
	assign \mchip.five.Q [0] = \mchip.five.Q_reg[0] ;
	reg \mchip.stop.Q_reg[0] ;
	always @(posedge io_in[12])
		if (\mchip.control.stop_clr )
			\mchip.stop.Q_reg[0]  <= 1'h0;
		else if (\mchip.control.stop_en )
			\mchip.stop.Q_reg[0]  <= _139_[0];
	assign \mchip.stop.Q [0] = \mchip.stop.Q_reg[0] ;
	reg \mchip.yellow.Q_reg[0] ;
	always @(posedge io_in[12])
		if (\mchip.control.yellow_clr )
			\mchip.yellow.Q_reg[0]  <= 1'h0;
		else if (\mchip.control.yellow_en )
			\mchip.yellow.Q_reg[0]  <= _140_[0];
	assign \mchip.yellow.Q [0] = \mchip.yellow.Q_reg[0] ;
	assign _000_[9:0] = 10'h000;
	assign _138_[7:1] = 7'h00;
	assign _139_[7:1] = 7'h00;
	assign _140_[7:1] = 7'h00;
	assign io_out[13:12] = 2'h0;
	assign \mchip.button  = io_in[0];
	assign \mchip.car1  = io_in[4];
	assign \mchip.car2  = io_in[3];
	assign \mchip.car3  = io_in[2];
	assign \mchip.car4  = io_in[1];
	assign \mchip.clock  = io_in[12];
	assign \mchip.control.car1  = io_in[4];
	assign \mchip.control.car2  = io_in[3];
	assign \mchip.control.car3  = io_in[2];
	assign \mchip.control.car4  = io_in[1];
	assign \mchip.control.clock  = io_in[12];
	assign \mchip.control.green1  = io_out[9];
	assign \mchip.control.green2  = io_out[6];
	assign \mchip.control.green3  = io_out[3];
	assign \mchip.control.orange  = io_out[1];
	assign \mchip.control.ped  = \mchip.pedestrian.ped ;
	assign \mchip.control.red1  = io_out[11];
	assign \mchip.control.red2  = io_out[8];
	assign \mchip.control.red3  = io_out[5];
	assign \mchip.control.reset  = io_in[13];
	assign \mchip.control.stop_five  = \mchip.five.Q [0];
	assign \mchip.control.stop_ped  = \mchip.stop.Q [0];
	assign \mchip.control.stop_yellow  = \mchip.yellow.Q [0];
	assign \mchip.control.turn  = io_out[2];
	assign \mchip.control.white  = io_out[0];
	assign \mchip.control.yellow1  = io_out[10];
	assign \mchip.control.yellow2  = io_out[7];
	assign \mchip.control.yellow3  = io_out[4];
	assign \mchip.five.D  = 8'h00;
	assign \mchip.five.Q [7:1] = 7'h00;
	assign \mchip.five.clear  = \mchip.control.five_clr ;
	assign \mchip.five.clock  = io_in[12];
	assign \mchip.five.en  = \mchip.control.five_en ;
	assign \mchip.five.load  = 1'h0;
	assign \mchip.five_clr  = \mchip.control.five_clr ;
	assign \mchip.five_en  = \mchip.control.five_en ;
	assign \mchip.green1  = io_out[9];
	assign \mchip.green2  = io_out[6];
	assign \mchip.green3  = io_out[3];
	assign \mchip.io_in  = io_in[11:0];
	assign \mchip.io_out  = io_out[11:0];
	assign \mchip.orange  = io_out[1];
	assign \mchip.ped  = \mchip.pedestrian.ped ;
	assign \mchip.ped_clr  = \mchip.control.ped_clr ;
	assign \mchip.pedestrian.button  = io_in[0];
	assign \mchip.pedestrian.clock  = io_in[12];
	assign \mchip.pedestrian.ped_clr  = \mchip.control.ped_clr ;
	assign \mchip.red1  = io_out[11];
	assign \mchip.red2  = io_out[8];
	assign \mchip.red3  = io_out[5];
	assign \mchip.reset  = io_in[13];
	assign \mchip.stop.D  = 8'h00;
	assign \mchip.stop.Q [7:1] = 7'h00;
	assign \mchip.stop.clear  = \mchip.control.stop_clr ;
	assign \mchip.stop.clock  = io_in[12];
	assign \mchip.stop.en  = \mchip.control.stop_en ;
	assign \mchip.stop.load  = 1'h0;
	assign \mchip.stop_clr  = \mchip.control.stop_clr ;
	assign \mchip.stop_en  = \mchip.control.stop_en ;
	assign \mchip.stop_five  = \mchip.five.Q [0];
	assign \mchip.stop_ped  = \mchip.stop.Q [0];
	assign \mchip.stop_yellow  = \mchip.yellow.Q [0];
	assign \mchip.turn  = io_out[2];
	assign \mchip.white  = io_out[0];
	assign \mchip.yellow.D  = 8'h00;
	assign \mchip.yellow.Q [7:1] = 7'h00;
	assign \mchip.yellow.clear  = \mchip.control.yellow_clr ;
	assign \mchip.yellow.clock  = io_in[12];
	assign \mchip.yellow.en  = \mchip.control.yellow_en ;
	assign \mchip.yellow.load  = 1'h0;
	assign \mchip.yellow1  = io_out[10];
	assign \mchip.yellow2  = io_out[7];
	assign \mchip.yellow3  = io_out[4];
	assign \mchip.yellow_clr  = \mchip.control.yellow_clr ;
	assign \mchip.yellow_en  = \mchip.control.yellow_en ;
endmodule
module d15_jerryfen_prng (
	io_in,
	io_out
);
	wire _000_;
	wire _001_;
	wire _002_;
	wire _003_;
	wire _004_;
	wire _005_;
	wire _006_;
	wire _007_;
	wire _008_;
	wire _009_;
	wire _010_;
	wire _011_;
	wire _012_;
	wire _013_;
	wire _014_;
	wire _015_;
	wire _016_;
	wire _017_;
	wire _018_;
	wire _019_;
	wire _020_;
	wire _021_;
	wire _022_;
	wire _023_;
	wire _024_;
	wire _025_;
	wire _026_;
	wire _027_;
	wire _028_;
	wire _029_;
	reg _030_;
	reg _031_;
	reg _032_;
	reg _033_;
	reg _034_;
	reg _035_;
	reg _036_;
	reg _037_;
	wire _038_;
	wire _039_;
	wire _040_;
	wire _041_;
	wire _042_;
	wire _043_;
	wire _044_;
	wire _045_;
	wire _046_;
	wire _047_;
	wire _048_;
	wire _049_;
	wire _050_;
	wire _051_;
	wire _052_;
	wire _053_;
	wire _054_;
	wire _055_;
	wire _056_;
	wire _057_;
	wire _058_;
	wire _059_;
	wire _060_;
	wire _061_;
	wire _062_;
	wire _063_;
	wire _064_;
	wire _065_;
	wire _066_;
	wire _067_;
	wire _068_;
	wire _069_;
	wire _070_;
	wire _071_;
	wire _072_;
	wire _073_;
	wire _074_;
	wire _075_;
	wire _076_;
	wire _077_;
	wire _078_;
	wire _079_;
	wire _080_;
	wire _081_;
	wire _082_;
	wire _083_;
	wire _084_;
	wire _085_;
	wire _086_;
	wire _087_;
	wire _088_;
	wire _089_;
	wire _090_;
	wire _091_;
	wire _092_;
	wire _093_;
	wire _094_;
	wire _095_;
	wire _096_;
	wire _097_;
	wire _098_;
	wire _099_;
	wire _100_;
	wire _101_;
	wire _102_;
	wire _103_;
	wire _104_;
	wire _105_;
	wire _106_;
	wire _107_;
	wire _108_;
	wire _109_;
	wire _110_;
	wire _111_;
	wire _112_;
	wire _113_;
	wire _114_;
	wire _115_;
	wire _116_;
	wire _117_;
	wire _118_;
	wire _119_;
	wire _120_;
	wire _121_;
	wire _122_;
	wire _123_;
	wire _124_;
	wire _125_;
	wire _126_;
	wire _127_;
	wire _128_;
	wire _129_;
	wire _130_;
	wire _131_;
	wire _132_;
	wire _133_;
	wire _134_;
	wire _135_;
	wire _136_;
	wire _137_;
	wire _138_;
	wire _139_;
	wire _140_;
	wire _141_;
	wire _142_;
	wire _143_;
	wire _144_;
	wire _145_;
	wire _146_;
	wire _147_;
	wire _148_;
	wire _149_;
	wire _150_;
	wire _151_;
	wire _152_;
	wire _153_;
	wire _154_;
	wire _155_;
	wire _156_;
	wire _157_;
	wire _158_;
	wire _159_;
	wire _160_;
	wire _161_;
	wire _162_;
	wire _163_;
	wire _164_;
	wire _165_;
	wire _166_;
	wire _167_;
	wire _168_;
	wire _169_;
	wire _170_;
	wire _171_;
	wire _172_;
	wire _173_;
	wire _174_;
	wire _175_;
	wire _176_;
	wire _177_;
	wire _178_;
	wire _179_;
	wire _180_;
	wire _181_;
	wire _182_;
	wire _183_;
	wire _184_;
	wire _185_;
	wire _186_;
	wire _187_;
	wire _188_;
	wire _189_;
	wire _190_;
	wire _191_;
	wire _192_;
	wire _193_;
	wire _194_;
	wire _195_;
	wire _196_;
	wire _197_;
	wire _198_;
	wire _199_;
	wire _200_;
	wire _201_;
	wire _202_;
	input wire [13:0] io_in;
	output wire [13:0] io_out;
	wire \mchip.clock ;
	wire [11:0] \mchip.io_in ;
	wire [11:0] \mchip.io_out ;
	wire [7:0] \mchip.prng_chip_one.AES_out_num ;
	wire \mchip.prng_chip_one.Sbox1.S0 ;
	wire \mchip.prng_chip_one.Sbox1.S1 ;
	wire \mchip.prng_chip_one.Sbox1.S2 ;
	wire \mchip.prng_chip_one.Sbox1.S3 ;
	wire \mchip.prng_chip_one.Sbox1.S4 ;
	wire \mchip.prng_chip_one.Sbox1.S5 ;
	wire \mchip.prng_chip_one.Sbox1.S6 ;
	wire \mchip.prng_chip_one.Sbox1.S7 ;
	wire \mchip.prng_chip_one.Sbox1.U0 ;
	wire \mchip.prng_chip_one.Sbox1.U1 ;
	wire \mchip.prng_chip_one.Sbox1.U2 ;
	wire \mchip.prng_chip_one.Sbox1.U3 ;
	wire \mchip.prng_chip_one.Sbox1.U4 ;
	wire \mchip.prng_chip_one.Sbox1.U5 ;
	wire \mchip.prng_chip_one.Sbox1.U6 ;
	wire \mchip.prng_chip_one.Sbox1.U7 ;
	wire [7:0] \mchip.prng_chip_one.Sbox1.input_num ;
	wire [7:0] \mchip.prng_chip_one.Sbox1.output_num ;
	wire \mchip.prng_chip_one.clk ;
	wire \mchip.prng_chip_one.cnt_en ;
	wire [7:0] \mchip.prng_chip_one.counter1.D ;
	wire \mchip.prng_chip_one.counter1.clear ;
	wire \mchip.prng_chip_one.counter1.clock ;
	wire \mchip.prng_chip_one.counter1.en ;
	wire \mchip.prng_chip_one.counter1.up ;
	wire \mchip.prng_chip_one.ctrl_pth1.clock ;
	wire \mchip.prng_chip_one.ctrl_pth1.cnt_en ;
	reg [3:0] \mchip.prng_chip_one.ctrl_pth1.curr_state ;
	wire \mchip.prng_chip_one.ctrl_pth1.enable ;
	wire \mchip.prng_chip_one.ctrl_pth1.reg_en ;
	wire \mchip.prng_chip_one.ctrl_pth1.reset ;
	wire \mchip.prng_chip_one.ctrl_pth1.sipo_en ;
	wire \mchip.prng_chip_one.ctrl_pth1.valid ;
	wire \mchip.prng_chip_one.en ;
	wire \mchip.prng_chip_one.fibo1.clk ;
	wire \mchip.prng_chip_one.fibo1.reset ;
	reg [7:0] \mchip.prng_chip_one.fibo1.state_out ;
	wire \mchip.prng_chip_one.galo1.clk ;
	wire \mchip.prng_chip_one.galo1.feedback ;
	wire \mchip.prng_chip_one.galo1.out_num ;
	wire \mchip.prng_chip_one.galo1.reset ;
	reg [7:0] \mchip.prng_chip_one.galo1.state_out ;
	wire \mchip.prng_chip_one.galo_out ;
	wire [7:0] \mchip.prng_chip_one.lsfr_rand_num ;
	wire [7:0] \mchip.prng_chip_one.magcomp1.B ;
	wire \mchip.prng_chip_one.mux1.I1 ;
	wire \mchip.prng_chip_one.mux1.S ;
	wire \mchip.prng_chip_one.mux1.Y ;
	wire [7:0] \mchip.prng_chip_one.rand_num ;
	wire [7:0] \mchip.prng_chip_one.reg1.D ;
	reg [7:0] \mchip.prng_chip_one.reg1.Q ;
	wire \mchip.prng_chip_one.reg1.clear ;
	wire \mchip.prng_chip_one.reg1.clock ;
	wire \mchip.prng_chip_one.reg1.en ;
	wire \mchip.prng_chip_one.reg_en ;
	wire [7:0] \mchip.prng_chip_one.reg_rand_num ;
	wire \mchip.prng_chip_one.reset ;
	wire [7:0] \mchip.prng_chip_one.seed ;
	wire \mchip.prng_chip_one.sel ;
	wire \mchip.prng_chip_one.serial_input ;
	wire \mchip.prng_chip_one.sipo_en ;
	wire [7:0] \mchip.prng_chip_one.sr_sipo1.D ;
	reg [7:0] \mchip.prng_chip_one.sr_sipo1.Q ;
	wire \mchip.prng_chip_one.sr_sipo1.clock ;
	wire \mchip.prng_chip_one.sr_sipo1.en ;
	wire \mchip.prng_chip_one.sr_sipo1.left ;
	wire \mchip.prng_chip_one.sr_sipo1.serial ;
	wire \mchip.prng_chip_one.valid ;
	wire \mchip.reset ;
	assign _193_ = io_in[0] | io_in[13];
	assign _194_ = \mchip.prng_chip_one.ctrl_pth1.curr_state [2] & ~_193_;
	assign _195_ = \mchip.prng_chip_one.ctrl_pth1.curr_state [0] & ~io_in[13];
	assign _003_ = _195_ | _194_;
	assign _196_ = io_in[13] | ~io_in[0];
	assign _197_ = \mchip.prng_chip_one.ctrl_pth1.curr_state [2] & ~_196_;
	assign _198_ = io_in[13] | ~_031_;
	assign _199_ = _030_ & ~io_in[13];
	assign _200_ = _198_ & ~_199_;
	assign _201_ = _032_ & ~io_in[13];
	assign _202_ = io_in[13] | ~_033_;
	assign _038_ = _202_ | _201_;
	assign _039_ = _200_ & ~_038_;
	assign _040_ = _037_ & ~io_in[13];
	assign _041_ = _036_ & ~io_in[13];
	assign _042_ = _041_ | _040_;
	assign _043_ = _035_ & ~io_in[13];
	assign _044_ = _034_ & ~io_in[13];
	assign _045_ = _044_ | _043_;
	assign _046_ = _045_ | _042_;
	assign _047_ = _039_ & ~_046_;
	assign _048_ = _047_ | io_in[13];
	assign _049_ = \mchip.prng_chip_one.ctrl_pth1.curr_state [1] & ~_048_;
	assign _002_ = _049_ | _197_;
	assign _050_ = \mchip.prng_chip_one.fibo1.state_out [4] ^ \mchip.prng_chip_one.fibo1.state_out [7];
	assign _051_ = _050_ ^ \mchip.prng_chip_one.fibo1.state_out [2];
	assign \mchip.prng_chip_one.sr_sipo1.serial  = (io_in[1] ? \mchip.prng_chip_one.galo1.state_out [7] : _051_);
	assign _052_ = \mchip.prng_chip_one.reg1.Q [0] ^ io_in[2];
	assign _053_ = \mchip.prng_chip_one.ctrl_pth1.curr_state [0] | \mchip.prng_chip_one.ctrl_pth1.curr_state [1];
	assign _054_ = ~(_053_ | \mchip.prng_chip_one.ctrl_pth1.curr_state [3]);
	assign _055_ = ~(_054_ & io_in[0]);
	assign _014_ = (_055_ ? _051_ : _052_);
	assign _056_ = \mchip.prng_chip_one.reg1.Q [1] ^ io_in[3];
	assign _015_ = (_055_ ? \mchip.prng_chip_one.fibo1.state_out [0] : _056_);
	assign _057_ = \mchip.prng_chip_one.reg1.Q [2] ^ io_in[4];
	assign _016_ = (_055_ ? \mchip.prng_chip_one.fibo1.state_out [1] : _057_);
	assign _058_ = \mchip.prng_chip_one.reg1.Q [3] ^ io_in[5];
	assign _017_ = (_055_ ? \mchip.prng_chip_one.fibo1.state_out [2] : _058_);
	assign _059_ = \mchip.prng_chip_one.reg1.Q [4] ^ io_in[6];
	assign _018_ = (_055_ ? \mchip.prng_chip_one.fibo1.state_out [3] : _059_);
	assign _060_ = \mchip.prng_chip_one.reg1.Q [5] ^ io_in[7];
	assign _019_ = (_055_ ? \mchip.prng_chip_one.fibo1.state_out [4] : _060_);
	assign _061_ = \mchip.prng_chip_one.reg1.Q [6] ^ io_in[8];
	assign _020_ = (_055_ ? \mchip.prng_chip_one.fibo1.state_out [5] : _061_);
	assign _062_ = \mchip.prng_chip_one.reg1.Q [7] ^ io_in[9];
	assign _021_ = (_055_ ? \mchip.prng_chip_one.fibo1.state_out [6] : _062_);
	assign _029_ = (_055_ ? \mchip.prng_chip_one.galo1.state_out [6] : _062_);
	assign _063_ = \mchip.prng_chip_one.galo1.state_out [5] ^ \mchip.prng_chip_one.galo1.state_out [7];
	assign _028_ = (_055_ ? _063_ : _061_);
	assign _064_ = \mchip.prng_chip_one.galo1.state_out [4] ^ \mchip.prng_chip_one.galo1.state_out [7];
	assign _027_ = (_055_ ? _064_ : _060_);
	assign _023_ = (_055_ ? \mchip.prng_chip_one.galo1.state_out [7] : _052_);
	assign _024_ = (_055_ ? \mchip.prng_chip_one.galo1.state_out [0] : _056_);
	assign _025_ = (_055_ ? \mchip.prng_chip_one.galo1.state_out [1] : _057_);
	assign _026_ = (_055_ ? \mchip.prng_chip_one.galo1.state_out [2] : _058_);
	assign _065_ = \mchip.prng_chip_one.galo1.state_out [3] ^ \mchip.prng_chip_one.galo1.state_out [7];
	assign _022_ = (_055_ ? _065_ : _059_);
	assign _006_ = _055_ & ~_199_;
	assign _066_ = _199_ & ~_198_;
	assign _067_ = _066_ | _200_;
	assign _007_ = _055_ & ~_067_;
	assign _068_ = ~_201_;
	assign _069_ = _066_ ^ _068_;
	assign _008_ = _055_ & ~_069_;
	assign _070_ = _066_ & ~_068_;
	assign _071_ = _070_ ^ _202_;
	assign _009_ = _055_ & ~_071_;
	assign _072_ = ~_044_;
	assign _073_ = _202_ | ~_201_;
	assign _074_ = _066_ & ~_073_;
	assign _075_ = _074_ ^ _072_;
	assign _010_ = _055_ & ~_075_;
	assign _076_ = ~(_074_ & _044_);
	assign _077_ = _076_ ^ _043_;
	assign _011_ = _055_ & ~_077_;
	assign _078_ = ~(_044_ & _043_);
	assign _079_ = _074_ & ~_078_;
	assign _080_ = ~(_079_ ^ _041_);
	assign _012_ = _055_ & ~_080_;
	assign _081_ = ~(_079_ & _041_);
	assign _082_ = _081_ ^ _040_;
	assign _013_ = _055_ & ~_082_;
	assign _083_ = ~(\mchip.prng_chip_one.reg1.Q [7] ^ \mchip.prng_chip_one.reg1.Q [2]);
	assign _084_ = \mchip.prng_chip_one.reg1.Q [7] ^ \mchip.prng_chip_one.reg1.Q [1];
	assign _085_ = \mchip.prng_chip_one.reg1.Q [4] ^ \mchip.prng_chip_one.reg1.Q [2];
	assign _086_ = _085_ ^ _084_;
	assign _087_ = _086_ ^ \mchip.prng_chip_one.reg1.Q [3];
	assign _088_ = ~(_087_ ^ \mchip.prng_chip_one.reg1.Q [6]);
	assign _089_ = \mchip.prng_chip_one.reg1.Q [7] ^ \mchip.prng_chip_one.reg1.Q [4];
	assign _090_ = _089_ ^ _088_;
	assign _091_ = \mchip.prng_chip_one.reg1.Q [6] ^ \mchip.prng_chip_one.reg1.Q [5];
	assign _092_ = _091_ ^ _090_;
	assign _093_ = _092_ ^ _084_;
	assign _094_ = _084_ & ~_092_;
	assign _095_ = _091_ ^ \mchip.prng_chip_one.reg1.Q [0];
	assign _096_ = \mchip.prng_chip_one.reg1.Q [1] | ~_095_;
	assign _097_ = _096_ ^ _094_;
	assign _098_ = _087_ ^ \mchip.prng_chip_one.reg1.Q [2];
	assign _099_ = _098_ ^ _091_;
	assign _100_ = _099_ ^ _090_;
	assign _101_ = _085_ & ~_100_;
	assign _102_ = ~(_089_ & _088_);
	assign _103_ = ~(_102_ ^ _101_);
	assign _104_ = _103_ ^ _097_;
	assign _105_ = _104_ ^ _093_;
	assign _106_ = _095_ ^ \mchip.prng_chip_one.reg1.Q [1];
	assign _107_ = _106_ ^ _083_;
	assign _108_ = ~\mchip.prng_chip_one.reg1.Q [0];
	assign _109_ = _098_ ^ _108_;
	assign _110_ = _109_ | _107_;
	assign _111_ = _098_ & _086_;
	assign _112_ = _111_ ^ _110_;
	assign _113_ = _112_ ^ _088_;
	assign _114_ = ~(_113_ ^ _103_);
	assign _115_ = _105_ & ~_114_;
	assign _116_ = _099_ ^ _083_;
	assign _117_ = _099_ & ~_083_;
	assign _118_ = _117_ ^ _102_;
	assign _119_ = ~(_095_ ^ \mchip.prng_chip_one.reg1.Q [4]);
	assign _120_ = \mchip.prng_chip_one.reg1.Q [0] & ~_119_;
	assign _121_ = _120_ ^ _111_;
	assign _122_ = _121_ ^ _118_;
	assign _123_ = _122_ ^ _116_;
	assign _124_ = _123_ ^ _115_;
	assign _125_ = _092_ ^ \mchip.prng_chip_one.reg1.Q [7];
	assign _126_ = _095_ ^ \mchip.prng_chip_one.reg1.Q [7];
	assign _127_ = _090_ ^ \mchip.prng_chip_one.reg1.Q [0];
	assign _128_ = _126_ & ~_127_;
	assign _129_ = _128_ ^ _094_;
	assign _130_ = _129_ ^ _118_;
	assign _131_ = _130_ ^ _125_;
	assign _132_ = (_124_ ? _105_ : _131_);
	assign _133_ = _132_ ^ _105_;
	assign _134_ = ~_105_;
	assign _135_ = ~_131_;
	assign _136_ = (_124_ ? _134_ : _135_);
	assign _137_ = _131_ ^ _115_;
	assign _138_ = _137_ ^ _136_;
	assign _139_ = _131_ & ~_138_;
	assign _140_ = ~(_139_ ^ _133_);
	assign _141_ = ~_123_;
	assign _142_ = (_137_ ? _114_ : _141_);
	assign _143_ = (_131_ ? _132_ : _137_);
	assign _144_ = _143_ & ~_142_;
	assign _145_ = ~(_123_ ^ _114_);
	assign _146_ = _145_ ^ _144_;
	assign _147_ = _146_ ^ _140_;
	assign _148_ = _147_ | _083_;
	assign _149_ = _142_ ^ _132_;
	assign _150_ = ~(_149_ | _090_);
	assign _151_ = ~(_146_ & _095_);
	assign _152_ = _146_ ^ _142_;
	assign _153_ = ~(_152_ | _092_);
	assign _154_ = ~(_153_ ^ _151_);
	assign _155_ = ~(_149_ ^ _147_);
	assign _156_ = ~(_155_ | _100_);
	assign _157_ = _156_ ^ _154_;
	assign _158_ = _157_ ^ _150_;
	assign _159_ = _089_ & ~_149_;
	assign _160_ = _159_ ^ _158_;
	assign _161_ = _132_ & ~_108_;
	assign _162_ = ~(_140_ ^ _136_);
	assign _163_ = _098_ & ~_162_;
	assign _164_ = _163_ ^ _161_;
	assign _165_ = _084_ & ~_152_;
	assign _166_ = _165_ ^ _164_;
	assign _167_ = _099_ & ~_147_;
	assign _168_ = _167_ ^ _166_;
	assign _169_ = ~(_168_ ^ _157_);
	assign _170_ = _142_ | ~_126_;
	assign _171_ = _170_ ^ _169_;
	assign _172_ = _171_ ^ _160_;
	assign \mchip.prng_chip_one.Sbox1.S2  = _172_ ^ _148_;
	assign _173_ = ~(_140_ | _109_);
	assign _174_ = _173_ ^ _163_;
	assign _175_ = ~(_174_ ^ _154_);
	assign _176_ = _085_ & ~_155_;
	assign _177_ = ~(_176_ ^ _159_);
	assign _178_ = _140_ | _107_;
	assign _179_ = _178_ ^ _177_;
	assign _180_ = _086_ & ~_162_;
	assign _181_ = _180_ ^ _179_;
	assign \mchip.prng_chip_one.Sbox1.S3  = ~(_181_ ^ _175_);
	assign \mchip.prng_chip_one.Sbox1.S1  = ~(\mchip.prng_chip_one.Sbox1.S3  ^ _158_);
	assign _182_ = ~(_142_ | _127_);
	assign _183_ = _182_ ^ _153_;
	assign _184_ = _183_ ^ _164_;
	assign _185_ = _146_ & _106_;
	assign _186_ = ~(_185_ ^ _177_);
	assign _187_ = _186_ ^ _184_;
	assign \mchip.prng_chip_one.Sbox1.S6  = _187_ ^ _169_;
	assign \mchip.prng_chip_one.Sbox1.S7  = ~(_187_ ^ _165_);
	assign _188_ = io_in[13] | ~_047_;
	assign _000_ = \mchip.prng_chip_one.ctrl_pth1.curr_state [1] & ~_188_;
	assign _189_ = ~(_136_ | _119_);
	assign _190_ = _189_ ^ _179_;
	assign \mchip.prng_chip_one.Sbox1.S5  = _190_ ^ _171_;
	assign \mchip.prng_chip_one.Sbox1.S4  = _184_ ^ \mchip.prng_chip_one.Sbox1.S3 ;
	assign \mchip.prng_chip_one.Sbox1.S0  = _181_ ^ _158_;
	assign _191_ = \mchip.prng_chip_one.ctrl_pth1.curr_state [0] | \mchip.prng_chip_one.ctrl_pth1.curr_state [2];
	assign _192_ = _191_ | \mchip.prng_chip_one.ctrl_pth1.curr_state [3];
	assign \mchip.prng_chip_one.counter1.en  = ~(_192_ | _047_);
	assign _005_ = \mchip.prng_chip_one.counter1.en  | ~_055_;
	assign \mchip.prng_chip_one.ctrl_pth1.reg_en  = _047_ & ~_192_;
	assign _004_ = \mchip.prng_chip_one.ctrl_pth1.reg_en  | io_in[13];
	assign _001_ = \mchip.prng_chip_one.ctrl_pth1.curr_state [3] | io_in[13];
	always @(posedge io_in[12])
		if (!\mchip.prng_chip_one.counter1.en )
			\mchip.prng_chip_one.sr_sipo1.Q [0] <= 1'h0;
		else
			\mchip.prng_chip_one.sr_sipo1.Q [0] <= \mchip.prng_chip_one.sr_sipo1.serial ;
	always @(posedge io_in[12])
		if (!\mchip.prng_chip_one.counter1.en )
			\mchip.prng_chip_one.sr_sipo1.Q [1] <= 1'h0;
		else
			\mchip.prng_chip_one.sr_sipo1.Q [1] <= \mchip.prng_chip_one.sr_sipo1.Q [0];
	always @(posedge io_in[12])
		if (!\mchip.prng_chip_one.counter1.en )
			\mchip.prng_chip_one.sr_sipo1.Q [2] <= 1'h0;
		else
			\mchip.prng_chip_one.sr_sipo1.Q [2] <= \mchip.prng_chip_one.sr_sipo1.Q [1];
	always @(posedge io_in[12])
		if (!\mchip.prng_chip_one.counter1.en )
			\mchip.prng_chip_one.sr_sipo1.Q [3] <= 1'h0;
		else
			\mchip.prng_chip_one.sr_sipo1.Q [3] <= \mchip.prng_chip_one.sr_sipo1.Q [2];
	always @(posedge io_in[12])
		if (!\mchip.prng_chip_one.counter1.en )
			\mchip.prng_chip_one.sr_sipo1.Q [4] <= 1'h0;
		else
			\mchip.prng_chip_one.sr_sipo1.Q [4] <= \mchip.prng_chip_one.sr_sipo1.Q [3];
	always @(posedge io_in[12])
		if (!\mchip.prng_chip_one.counter1.en )
			\mchip.prng_chip_one.sr_sipo1.Q [5] <= 1'h0;
		else
			\mchip.prng_chip_one.sr_sipo1.Q [5] <= \mchip.prng_chip_one.sr_sipo1.Q [4];
	always @(posedge io_in[12])
		if (!\mchip.prng_chip_one.counter1.en )
			\mchip.prng_chip_one.sr_sipo1.Q [6] <= 1'h0;
		else
			\mchip.prng_chip_one.sr_sipo1.Q [6] <= \mchip.prng_chip_one.sr_sipo1.Q [5];
	always @(posedge io_in[12])
		if (!\mchip.prng_chip_one.counter1.en )
			\mchip.prng_chip_one.sr_sipo1.Q [7] <= 1'h0;
		else
			\mchip.prng_chip_one.sr_sipo1.Q [7] <= \mchip.prng_chip_one.sr_sipo1.Q [6];
	always @(posedge io_in[12])
		if (io_in[13])
			_030_ <= 1'h0;
		else if (_005_)
			_030_ <= _006_;
	always @(posedge io_in[12])
		if (io_in[13])
			_031_ <= 1'h0;
		else if (_005_)
			_031_ <= _007_;
	always @(posedge io_in[12])
		if (io_in[13])
			_032_ <= 1'h0;
		else if (_005_)
			_032_ <= _008_;
	always @(posedge io_in[12])
		if (io_in[13])
			_033_ <= 1'h0;
		else if (_005_)
			_033_ <= _009_;
	always @(posedge io_in[12])
		if (io_in[13])
			_034_ <= 1'h0;
		else if (_005_)
			_034_ <= _010_;
	always @(posedge io_in[12])
		if (io_in[13])
			_035_ <= 1'h0;
		else if (_005_)
			_035_ <= _011_;
	always @(posedge io_in[12])
		if (io_in[13])
			_036_ <= 1'h0;
		else if (_005_)
			_036_ <= _012_;
	always @(posedge io_in[12])
		if (io_in[13])
			_037_ <= 1'h0;
		else if (_005_)
			_037_ <= _013_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.prng_chip_one.fibo1.state_out [0] <= 1'h0;
		else
			\mchip.prng_chip_one.fibo1.state_out [0] <= _014_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.prng_chip_one.fibo1.state_out [1] <= 1'h0;
		else
			\mchip.prng_chip_one.fibo1.state_out [1] <= _015_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.prng_chip_one.fibo1.state_out [2] <= 1'h0;
		else
			\mchip.prng_chip_one.fibo1.state_out [2] <= _016_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.prng_chip_one.fibo1.state_out [3] <= 1'h0;
		else
			\mchip.prng_chip_one.fibo1.state_out [3] <= _017_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.prng_chip_one.fibo1.state_out [4] <= 1'h0;
		else
			\mchip.prng_chip_one.fibo1.state_out [4] <= _018_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.prng_chip_one.fibo1.state_out [5] <= 1'h0;
		else
			\mchip.prng_chip_one.fibo1.state_out [5] <= _019_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.prng_chip_one.fibo1.state_out [6] <= 1'h0;
		else
			\mchip.prng_chip_one.fibo1.state_out [6] <= _020_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.prng_chip_one.fibo1.state_out [7] <= 1'h0;
		else
			\mchip.prng_chip_one.fibo1.state_out [7] <= _021_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.prng_chip_one.galo1.state_out [0] <= 1'h0;
		else
			\mchip.prng_chip_one.galo1.state_out [0] <= _023_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.prng_chip_one.galo1.state_out [1] <= 1'h0;
		else
			\mchip.prng_chip_one.galo1.state_out [1] <= _024_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.prng_chip_one.galo1.state_out [2] <= 1'h0;
		else
			\mchip.prng_chip_one.galo1.state_out [2] <= _025_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.prng_chip_one.galo1.state_out [3] <= 1'h0;
		else
			\mchip.prng_chip_one.galo1.state_out [3] <= _026_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.prng_chip_one.galo1.state_out [4] <= 1'h0;
		else
			\mchip.prng_chip_one.galo1.state_out [4] <= _022_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.prng_chip_one.galo1.state_out [5] <= 1'h0;
		else
			\mchip.prng_chip_one.galo1.state_out [5] <= _027_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.prng_chip_one.galo1.state_out [6] <= 1'h0;
		else
			\mchip.prng_chip_one.galo1.state_out [6] <= _028_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.prng_chip_one.galo1.state_out [7] <= 1'h0;
		else
			\mchip.prng_chip_one.galo1.state_out [7] <= _029_;
	always @(posedge io_in[12])
		if (_004_)
			if (!\mchip.prng_chip_one.ctrl_pth1.reg_en )
				\mchip.prng_chip_one.reg1.Q [0] <= 1'h0;
			else
				\mchip.prng_chip_one.reg1.Q [0] <= \mchip.prng_chip_one.sr_sipo1.Q [0];
	always @(posedge io_in[12])
		if (_004_)
			if (!\mchip.prng_chip_one.ctrl_pth1.reg_en )
				\mchip.prng_chip_one.reg1.Q [1] <= 1'h0;
			else
				\mchip.prng_chip_one.reg1.Q [1] <= \mchip.prng_chip_one.sr_sipo1.Q [1];
	always @(posedge io_in[12])
		if (_004_)
			if (!\mchip.prng_chip_one.ctrl_pth1.reg_en )
				\mchip.prng_chip_one.reg1.Q [2] <= 1'h0;
			else
				\mchip.prng_chip_one.reg1.Q [2] <= \mchip.prng_chip_one.sr_sipo1.Q [2];
	always @(posedge io_in[12])
		if (_004_)
			if (!\mchip.prng_chip_one.ctrl_pth1.reg_en )
				\mchip.prng_chip_one.reg1.Q [3] <= 1'h0;
			else
				\mchip.prng_chip_one.reg1.Q [3] <= \mchip.prng_chip_one.sr_sipo1.Q [3];
	always @(posedge io_in[12])
		if (_004_)
			if (!\mchip.prng_chip_one.ctrl_pth1.reg_en )
				\mchip.prng_chip_one.reg1.Q [4] <= 1'h0;
			else
				\mchip.prng_chip_one.reg1.Q [4] <= \mchip.prng_chip_one.sr_sipo1.Q [4];
	always @(posedge io_in[12])
		if (_004_)
			if (!\mchip.prng_chip_one.ctrl_pth1.reg_en )
				\mchip.prng_chip_one.reg1.Q [5] <= 1'h0;
			else
				\mchip.prng_chip_one.reg1.Q [5] <= \mchip.prng_chip_one.sr_sipo1.Q [5];
	always @(posedge io_in[12])
		if (_004_)
			if (!\mchip.prng_chip_one.ctrl_pth1.reg_en )
				\mchip.prng_chip_one.reg1.Q [6] <= 1'h0;
			else
				\mchip.prng_chip_one.reg1.Q [6] <= \mchip.prng_chip_one.sr_sipo1.Q [6];
	always @(posedge io_in[12])
		if (_004_)
			if (!\mchip.prng_chip_one.ctrl_pth1.reg_en )
				\mchip.prng_chip_one.reg1.Q [7] <= 1'h0;
			else
				\mchip.prng_chip_one.reg1.Q [7] <= \mchip.prng_chip_one.sr_sipo1.Q [7];
	always @(posedge io_in[12]) \mchip.prng_chip_one.ctrl_pth1.curr_state [0] <= _001_;
	always @(posedge io_in[12]) \mchip.prng_chip_one.ctrl_pth1.curr_state [1] <= _002_;
	always @(posedge io_in[12]) \mchip.prng_chip_one.ctrl_pth1.curr_state [2] <= _003_;
	always @(posedge io_in[12]) \mchip.prng_chip_one.ctrl_pth1.curr_state [3] <= _000_;
	assign io_out = {5'h00, \mchip.prng_chip_one.ctrl_pth1.curr_state [3], \mchip.prng_chip_one.Sbox1.S3 , \mchip.prng_chip_one.Sbox1.S7 , \mchip.prng_chip_one.Sbox1.S0 , \mchip.prng_chip_one.Sbox1.S6 , \mchip.prng_chip_one.Sbox1.S4 , \mchip.prng_chip_one.Sbox1.S1 , \mchip.prng_chip_one.Sbox1.S2 , \mchip.prng_chip_one.Sbox1.S5 };
	assign \mchip.clock  = io_in[12];
	assign \mchip.io_in  = io_in[11:0];
	assign \mchip.io_out  = {3'h0, \mchip.prng_chip_one.ctrl_pth1.curr_state [3], \mchip.prng_chip_one.Sbox1.S3 , \mchip.prng_chip_one.Sbox1.S7 , \mchip.prng_chip_one.Sbox1.S0 , \mchip.prng_chip_one.Sbox1.S6 , \mchip.prng_chip_one.Sbox1.S4 , \mchip.prng_chip_one.Sbox1.S1 , \mchip.prng_chip_one.Sbox1.S2 , \mchip.prng_chip_one.Sbox1.S5 };
	assign \mchip.prng_chip_one.AES_out_num  = {\mchip.prng_chip_one.Sbox1.S3 , \mchip.prng_chip_one.Sbox1.S7 , \mchip.prng_chip_one.Sbox1.S0 , \mchip.prng_chip_one.Sbox1.S6 , \mchip.prng_chip_one.Sbox1.S4 , \mchip.prng_chip_one.Sbox1.S1 , \mchip.prng_chip_one.Sbox1.S2 , \mchip.prng_chip_one.Sbox1.S5 };
	assign \mchip.prng_chip_one.Sbox1.U0  = \mchip.prng_chip_one.reg1.Q [7];
	assign \mchip.prng_chip_one.Sbox1.U1  = \mchip.prng_chip_one.reg1.Q [6];
	assign \mchip.prng_chip_one.Sbox1.U2  = \mchip.prng_chip_one.reg1.Q [5];
	assign \mchip.prng_chip_one.Sbox1.U3  = \mchip.prng_chip_one.reg1.Q [4];
	assign \mchip.prng_chip_one.Sbox1.U4  = \mchip.prng_chip_one.reg1.Q [3];
	assign \mchip.prng_chip_one.Sbox1.U5  = \mchip.prng_chip_one.reg1.Q [2];
	assign \mchip.prng_chip_one.Sbox1.U6  = \mchip.prng_chip_one.reg1.Q [1];
	assign \mchip.prng_chip_one.Sbox1.U7  = \mchip.prng_chip_one.reg1.Q [0];
	assign \mchip.prng_chip_one.Sbox1.input_num  = \mchip.prng_chip_one.reg1.Q ;
	assign \mchip.prng_chip_one.Sbox1.output_num  = {\mchip.prng_chip_one.Sbox1.S3 , \mchip.prng_chip_one.Sbox1.S7 , \mchip.prng_chip_one.Sbox1.S0 , \mchip.prng_chip_one.Sbox1.S6 , \mchip.prng_chip_one.Sbox1.S4 , \mchip.prng_chip_one.Sbox1.S1 , \mchip.prng_chip_one.Sbox1.S2 , \mchip.prng_chip_one.Sbox1.S5 };
	assign \mchip.prng_chip_one.clk  = io_in[12];
	assign \mchip.prng_chip_one.cnt_en  = \mchip.prng_chip_one.counter1.en ;
	assign \mchip.prng_chip_one.counter1.D  = 8'h00;
	assign \mchip.prng_chip_one.counter1.clear  = io_in[13];
	assign \mchip.prng_chip_one.counter1.clock  = io_in[12];
	assign \mchip.prng_chip_one.counter1.up  = 1'h1;
	assign \mchip.prng_chip_one.ctrl_pth1.clock  = io_in[12];
	assign \mchip.prng_chip_one.ctrl_pth1.cnt_en  = \mchip.prng_chip_one.counter1.en ;
	assign \mchip.prng_chip_one.ctrl_pth1.enable  = io_in[0];
	assign \mchip.prng_chip_one.ctrl_pth1.reset  = io_in[13];
	assign \mchip.prng_chip_one.ctrl_pth1.sipo_en  = \mchip.prng_chip_one.counter1.en ;
	assign \mchip.prng_chip_one.ctrl_pth1.valid  = \mchip.prng_chip_one.ctrl_pth1.curr_state [3];
	assign \mchip.prng_chip_one.en  = io_in[0];
	assign \mchip.prng_chip_one.fibo1.clk  = io_in[12];
	assign \mchip.prng_chip_one.fibo1.reset  = io_in[13];
	assign \mchip.prng_chip_one.galo1.clk  = io_in[12];
	assign \mchip.prng_chip_one.galo1.feedback  = \mchip.prng_chip_one.galo1.state_out [7];
	assign \mchip.prng_chip_one.galo1.out_num  = \mchip.prng_chip_one.galo1.state_out [7];
	assign \mchip.prng_chip_one.galo1.reset  = io_in[13];
	assign \mchip.prng_chip_one.galo_out  = \mchip.prng_chip_one.galo1.state_out [7];
	assign \mchip.prng_chip_one.lsfr_rand_num  = \mchip.prng_chip_one.sr_sipo1.Q ;
	assign \mchip.prng_chip_one.magcomp1.B  = 8'h08;
	assign \mchip.prng_chip_one.mux1.I1  = \mchip.prng_chip_one.galo1.state_out [7];
	assign \mchip.prng_chip_one.mux1.S  = io_in[1];
	assign \mchip.prng_chip_one.mux1.Y  = \mchip.prng_chip_one.sr_sipo1.serial ;
	assign \mchip.prng_chip_one.rand_num  = {\mchip.prng_chip_one.Sbox1.S3 , \mchip.prng_chip_one.Sbox1.S7 , \mchip.prng_chip_one.Sbox1.S0 , \mchip.prng_chip_one.Sbox1.S6 , \mchip.prng_chip_one.Sbox1.S4 , \mchip.prng_chip_one.Sbox1.S1 , \mchip.prng_chip_one.Sbox1.S2 , \mchip.prng_chip_one.Sbox1.S5 };
	assign \mchip.prng_chip_one.reg1.D  = \mchip.prng_chip_one.sr_sipo1.Q ;
	assign \mchip.prng_chip_one.reg1.clear  = io_in[13];
	assign \mchip.prng_chip_one.reg1.clock  = io_in[12];
	assign \mchip.prng_chip_one.reg1.en  = \mchip.prng_chip_one.ctrl_pth1.reg_en ;
	assign \mchip.prng_chip_one.reg_en  = \mchip.prng_chip_one.ctrl_pth1.reg_en ;
	assign \mchip.prng_chip_one.reg_rand_num  = \mchip.prng_chip_one.reg1.Q ;
	assign \mchip.prng_chip_one.reset  = io_in[13];
	assign \mchip.prng_chip_one.seed  = io_in[9:2];
	assign \mchip.prng_chip_one.sel  = io_in[1];
	assign \mchip.prng_chip_one.serial_input  = \mchip.prng_chip_one.sr_sipo1.serial ;
	assign \mchip.prng_chip_one.sipo_en  = \mchip.prng_chip_one.counter1.en ;
	assign \mchip.prng_chip_one.sr_sipo1.D  = 8'h00;
	assign \mchip.prng_chip_one.sr_sipo1.clock  = io_in[12];
	assign \mchip.prng_chip_one.sr_sipo1.en  = \mchip.prng_chip_one.counter1.en ;
	assign \mchip.prng_chip_one.sr_sipo1.left  = 1'h1;
	assign \mchip.prng_chip_one.valid  = \mchip.prng_chip_one.ctrl_pth1.curr_state [3];
	assign \mchip.reset  = io_in[13];
endmodule
module d16_bgonzale_pll (
	io_in,
	io_out
);
	wire _000_;
	wire _001_;
	wire _002_;
	wire _003_;
	wire _004_;
	wire _005_;
	wire _006_;
	wire _007_;
	wire _008_;
	wire _009_;
	wire _010_;
	wire _011_;
	wire _012_;
	wire _013_;
	wire _014_;
	wire _015_;
	wire _016_;
	wire _017_;
	wire _018_;
	wire _019_;
	wire _020_;
	wire _021_;
	wire _022_;
	wire _023_;
	wire _024_;
	wire _025_;
	wire _026_;
	wire _027_;
	wire _028_;
	wire _029_;
	wire _030_;
	wire _031_;
	wire _032_;
	wire _033_;
	wire _034_;
	wire _035_;
	wire _036_;
	wire _037_;
	wire _038_;
	wire _039_;
	wire _040_;
	wire _041_;
	wire _042_;
	wire _043_;
	wire _044_;
	wire _045_;
	wire _046_;
	wire _047_;
	wire _048_;
	wire _049_;
	wire _050_;
	wire _051_;
	wire _052_;
	wire _053_;
	wire _054_;
	wire _055_;
	wire _056_;
	wire _057_;
	wire _058_;
	wire _059_;
	wire _060_;
	wire _061_;
	wire _062_;
	wire _063_;
	wire _064_;
	wire _065_;
	wire _066_;
	wire _067_;
	wire _068_;
	wire _069_;
	wire _070_;
	wire _071_;
	wire _072_;
	wire _073_;
	wire _074_;
	wire _075_;
	wire _076_;
	wire _077_;
	wire _078_;
	wire _079_;
	wire _080_;
	wire _081_;
	wire _082_;
	wire _083_;
	wire _084_;
	wire _085_;
	wire _086_;
	wire _087_;
	wire _088_;
	wire _089_;
	wire _090_;
	wire _091_;
	wire _092_;
	wire _093_;
	wire _094_;
	wire _095_;
	wire _096_;
	wire _097_;
	wire _098_;
	wire _099_;
	wire _100_;
	wire _101_;
	wire _102_;
	wire _103_;
	wire _104_;
	wire _105_;
	wire _106_;
	wire _107_;
	wire _108_;
	wire _109_;
	wire _110_;
	wire _111_;
	wire _112_;
	wire _113_;
	wire _114_;
	wire _115_;
	wire _116_;
	wire _117_;
	wire _118_;
	wire _119_;
	wire _120_;
	wire _121_;
	wire _122_;
	wire _123_;
	wire _124_;
	wire _125_;
	wire _126_;
	wire _127_;
	wire _128_;
	wire _129_;
	wire _130_;
	wire _131_;
	wire _132_;
	wire _133_;
	wire _134_;
	wire _135_;
	wire _136_;
	wire _137_;
	wire _138_;
	wire _139_;
	wire _140_;
	wire _141_;
	wire _142_;
	wire _143_;
	wire _144_;
	wire _145_;
	wire _146_;
	wire _147_;
	wire _148_;
	wire _149_;
	wire _150_;
	wire _151_;
	wire _152_;
	wire _153_;
	wire _154_;
	wire _155_;
	wire _156_;
	wire _157_;
	wire _158_;
	wire _159_;
	wire _160_;
	wire _161_;
	wire _162_;
	wire _163_;
	wire _164_;
	wire _165_;
	wire _166_;
	wire _167_;
	wire _168_;
	wire _169_;
	wire _170_;
	wire _171_;
	wire _172_;
	wire _173_;
	wire _174_;
	wire _175_;
	wire _176_;
	wire _177_;
	wire _178_;
	wire _179_;
	wire _180_;
	wire [8:0] _181_;
	wire [8:0] _182_;
	input wire [13:0] io_in;
	output wire [13:0] io_out;
	reg [7:0] \mchip.PLL.dig_osc.ctr ;
	wire [7:0] \mchip.PLL.dig_osc.freq_step ;
	wire \mchip.PLL.dig_osc.i_sys_clk ;
	wire \mchip.PLL.dig_osc.lead_or_lag ;
	wire \mchip.PLL.dig_osc.out_of_phase ;
	wire [7:0] \mchip.PLL.dig_osc.phase_corr ;
	wire \mchip.PLL.dig_osc.rec_clk ;
	wire [7:0] \mchip.PLL.i_freq_step ;
	wire [2:0] \mchip.PLL.i_loop_gain ;
	wire \mchip.PLL.i_ref_clk ;
	wire \mchip.PLL.i_sys_clk ;
	wire \mchip.PLL.lead_or_lag ;
	wire \mchip.PLL.loop_fil.i_sys_clk ;
	wire [2:0] \mchip.PLL.loop_fil.loop_gain ;
	reg [7:0] \mchip.PLL.loop_fil.phase_corr  = 8'h00;
	wire \mchip.PLL.o_lead_or_lag ;
	wire \mchip.PLL.o_phase_error ;
	wire \mchip.PLL.o_rec_clk ;
	wire \mchip.PLL.out_of_phase ;
	wire [7:0] \mchip.PLL.phase_corr ;
	wire \mchip.PLL.phase_det.i_sys_clk ;
	wire \mchip.PLL.phase_det.lead_or_lag ;
	reg \mchip.PLL.phase_det.matched  = 1'h0;
	wire \mchip.PLL.phase_det.out_of_phase ;
	wire \mchip.PLL.phase_det.rec_clk ;
	wire \mchip.PLL.phase_det.ref_clk ;
	wire \mchip.clock ;
	reg [8:0] \mchip.counter ;
	wire [11:0] \mchip.io_in ;
	wire [11:0] \mchip.io_out ;
	reg \mchip.new_clock ;
	wire \mchip.reset ;
	assign _148_ = \mchip.PLL.dig_osc.ctr [5] & io_in[9];
	assign _149_ = \mchip.PLL.dig_osc.ctr [4] & io_in[8];
	assign _150_ = \mchip.PLL.dig_osc.ctr [5] ^ io_in[9];
	assign _151_ = _150_ & _149_;
	assign _152_ = _151_ | _148_;
	assign _153_ = ~(\mchip.PLL.dig_osc.ctr [3] & io_in[7]);
	assign _154_ = \mchip.PLL.dig_osc.ctr [2] & io_in[6];
	assign _155_ = \mchip.PLL.dig_osc.ctr [3] ^ io_in[7];
	assign _156_ = _155_ & _154_;
	assign _157_ = _153_ & ~_156_;
	assign _158_ = \mchip.PLL.dig_osc.ctr [2] ^ io_in[6];
	assign _159_ = _158_ & _155_;
	assign _160_ = ~(io_in[5] & \mchip.PLL.dig_osc.ctr [1]);
	assign _161_ = io_in[4] & \mchip.PLL.dig_osc.ctr [0];
	assign _162_ = io_in[5] ^ \mchip.PLL.dig_osc.ctr [1];
	assign _163_ = _162_ & _161_;
	assign _164_ = _160_ & ~_163_;
	assign _165_ = _159_ & ~_164_;
	assign _166_ = _157_ & ~_165_;
	assign _167_ = \mchip.PLL.dig_osc.ctr [4] ^ io_in[8];
	assign _168_ = ~(_150_ & _167_);
	assign _169_ = ~(_168_ | _166_);
	assign _170_ = _169_ | _152_;
	assign _171_ = ~(io_in[10] ^ \mchip.PLL.dig_osc.ctr [6]);
	assign _172_ = ~(_171_ ^ _170_);
	assign _173_ = ~\mchip.PLL.loop_fil.phase_corr [4];
	assign _174_ = ~(\mchip.PLL.loop_fil.phase_corr [1] | \mchip.PLL.loop_fil.phase_corr [0]);
	assign _175_ = \mchip.PLL.loop_fil.phase_corr [2] | \mchip.PLL.loop_fil.phase_corr [3];
	assign _176_ = _174_ & ~_175_;
	assign _177_ = ~(_176_ & _173_);
	assign _178_ = _177_ ^ \mchip.PLL.loop_fil.phase_corr [5];
	assign _179_ = \mchip.PLL.dig_osc.ctr [7] & ~io_in[0];
	assign _180_ = io_in[0] & ~\mchip.PLL.dig_osc.ctr [7];
	assign \mchip.PLL.dig_osc.lead_or_lag  = (\mchip.PLL.phase_det.matched  ? _180_ : _179_);
	assign _016_ = ~(\mchip.PLL.loop_fil.phase_corr [7] ^ io_in[11]);
	assign _017_ = io_in[10] ^ \mchip.PLL.loop_fil.phase_corr [6];
	assign _018_ = _016_ & ~_017_;
	assign _019_ = \mchip.PLL.loop_fil.phase_corr [4] ^ io_in[8];
	assign _020_ = io_in[9] ^ \mchip.PLL.loop_fil.phase_corr [5];
	assign _021_ = _020_ | _019_;
	assign _022_ = _018_ & ~_021_;
	assign _023_ = \mchip.PLL.loop_fil.phase_corr [0] ^ io_in[4];
	assign _024_ = \mchip.PLL.loop_fil.phase_corr [1] ^ io_in[5];
	assign _025_ = ~(_024_ | _023_);
	assign _026_ = ~(io_in[6] ^ \mchip.PLL.loop_fil.phase_corr [2]);
	assign _027_ = io_in[7] ^ \mchip.PLL.loop_fil.phase_corr [3];
	assign _028_ = _026_ & ~_027_;
	assign _029_ = ~(_028_ & _025_);
	assign _030_ = _022_ & ~_029_;
	assign _031_ = \mchip.PLL.loop_fil.phase_corr [7] | ~io_in[11];
	assign _032_ = \mchip.PLL.loop_fil.phase_corr [6] | ~io_in[10];
	assign _033_ = _016_ & ~_032_;
	assign _034_ = _031_ & ~_033_;
	assign _035_ = \mchip.PLL.loop_fil.phase_corr [5] | ~io_in[9];
	assign _036_ = io_in[8] & ~\mchip.PLL.loop_fil.phase_corr [4];
	assign _037_ = _036_ & ~_020_;
	assign _038_ = _035_ & ~_037_;
	assign _039_ = _018_ & ~_038_;
	assign _040_ = _034_ & ~_039_;
	assign _041_ = \mchip.PLL.loop_fil.phase_corr [3] | ~io_in[7];
	assign _042_ = io_in[6] & ~\mchip.PLL.loop_fil.phase_corr [2];
	assign _043_ = _042_ & ~_027_;
	assign _044_ = _041_ & ~_043_;
	assign _045_ = \mchip.PLL.loop_fil.phase_corr [1] | ~io_in[5];
	assign _046_ = io_in[4] | ~\mchip.PLL.loop_fil.phase_corr [0];
	assign _047_ = _046_ & ~_024_;
	assign _048_ = _045_ & ~_047_;
	assign _049_ = _028_ & ~_048_;
	assign _050_ = _044_ & ~_049_;
	assign _051_ = _022_ & ~_050_;
	assign _052_ = _040_ & ~_051_;
	assign _053_ = _052_ | _030_;
	assign _054_ = \mchip.PLL.dig_osc.lead_or_lag  & ~_053_;
	assign _055_ = (_054_ ? \mchip.PLL.loop_fil.phase_corr [5] : _178_);
	assign _056_ = _167_ & ~_166_;
	assign _057_ = ~(_056_ | _149_);
	assign _058_ = ~(_150_ ^ _057_);
	assign _059_ = _058_ & ~_055_;
	assign _060_ = _176_ ^ _173_;
	assign _061_ = (_054_ ? \mchip.PLL.loop_fil.phase_corr [4] : _060_);
	assign _062_ = ~(_166_ ^ _167_);
	assign _063_ = _062_ & ~_061_;
	assign _064_ = _058_ ^ _055_;
	assign _065_ = _063_ & ~_064_;
	assign _066_ = _065_ | _059_;
	assign _067_ = ~\mchip.PLL.loop_fil.phase_corr [1];
	assign _068_ = \mchip.PLL.loop_fil.phase_corr [1] ^ \mchip.PLL.loop_fil.phase_corr [0];
	assign _069_ = ~_068_;
	assign _070_ = (_054_ ? _067_ : _069_);
	assign _071_ = _162_ ^ _161_;
	assign _072_ = _071_ ^ _070_;
	assign _073_ = io_in[4] ^ \mchip.PLL.dig_osc.ctr [0];
	assign _074_ = \mchip.PLL.loop_fil.phase_corr [0] & ~_073_;
	assign _075_ = _072_ & ~_074_;
	assign _076_ = _071_ & _070_;
	assign _077_ = _076_ | _075_;
	assign _078_ = \mchip.PLL.loop_fil.phase_corr [2] | ~_174_;
	assign _079_ = _078_ ^ \mchip.PLL.loop_fil.phase_corr [3];
	assign _080_ = (_054_ ? \mchip.PLL.loop_fil.phase_corr [3] : _079_);
	assign _081_ = ~_158_;
	assign _082_ = _164_ | _081_;
	assign _083_ = _082_ & ~_154_;
	assign _084_ = ~(_083_ ^ _155_);
	assign _085_ = _084_ ^ _080_;
	assign _086_ = ~(_174_ ^ \mchip.PLL.loop_fil.phase_corr [2]);
	assign _087_ = (_054_ ? \mchip.PLL.loop_fil.phase_corr [2] : _086_);
	assign _088_ = _164_ ^ _081_;
	assign _089_ = _088_ ^ _087_;
	assign _090_ = _089_ | _085_;
	assign _091_ = _077_ & ~_090_;
	assign _092_ = _084_ & ~_080_;
	assign _093_ = _087_ | ~_088_;
	assign _094_ = ~(_093_ | _085_);
	assign _095_ = _094_ | _092_;
	assign _096_ = _095_ | _091_;
	assign _097_ = _062_ ^ _061_;
	assign _098_ = _097_ | _064_;
	assign _099_ = _096_ & ~_098_;
	assign _100_ = _099_ | _066_;
	assign _101_ = ~\mchip.PLL.loop_fil.phase_corr [6];
	assign _102_ = \mchip.PLL.loop_fil.phase_corr [4] | \mchip.PLL.loop_fil.phase_corr [5];
	assign _103_ = _176_ & ~_102_;
	assign _104_ = _103_ ^ \mchip.PLL.loop_fil.phase_corr [6];
	assign _105_ = (_054_ ? _101_ : _104_);
	assign _106_ = _172_ ^ _105_;
	assign _107_ = _106_ ^ _100_;
	assign _108_ = ~(_180_ | _179_);
	assign _008_ = (_108_ ? _172_ : _107_);
	assign _109_ = _170_ & ~_171_;
	assign _110_ = io_in[10] & \mchip.PLL.dig_osc.ctr [6];
	assign _111_ = _110_ | _109_;
	assign _112_ = \mchip.PLL.dig_osc.ctr [7] ^ io_in[11];
	assign _113_ = _112_ ^ _111_;
	assign _114_ = _172_ & _105_;
	assign _115_ = _106_ & _100_;
	assign _116_ = _115_ | _114_;
	assign _117_ = ~\mchip.PLL.loop_fil.phase_corr [7];
	assign _118_ = _103_ & ~\mchip.PLL.loop_fil.phase_corr [6];
	assign _119_ = _118_ ^ \mchip.PLL.loop_fil.phase_corr [7];
	assign _120_ = (_054_ ? _117_ : _119_);
	assign _121_ = _113_ ^ _120_;
	assign _122_ = _121_ ^ _116_;
	assign _009_ = (_108_ ? _113_ : _122_);
	assign _182_[1] = \mchip.counter [0] ^ \mchip.counter [1];
	assign _123_ = \mchip.counter [0] & \mchip.counter [1];
	assign _182_[2] = _123_ ^ \mchip.counter [2];
	assign _124_ = _123_ & \mchip.counter [2];
	assign _182_[3] = _124_ ^ \mchip.counter [3];
	assign _125_ = ~(\mchip.counter [3] & \mchip.counter [2]);
	assign _126_ = _123_ & ~_125_;
	assign _182_[4] = _126_ ^ \mchip.counter [4];
	assign _127_ = _126_ & \mchip.counter [4];
	assign _182_[5] = _127_ ^ \mchip.counter [5];
	assign _128_ = ~(\mchip.counter [5] & \mchip.counter [4]);
	assign _129_ = _126_ & ~_128_;
	assign _182_[6] = _129_ ^ \mchip.counter [6];
	assign _130_ = _129_ & \mchip.counter [6];
	assign _182_[7] = _130_ ^ \mchip.counter [7];
	assign _131_ = ~(\mchip.counter [7] & \mchip.counter [6]);
	assign _132_ = _131_ | _128_;
	assign _133_ = _126_ & ~_132_;
	assign _182_[8] = _133_ ^ \mchip.counter [8];
	assign _012_ = io_in[1] & io_in[2];
	assign _013_ = io_in[2] & ~io_in[1];
	assign _014_ = io_in[1] & ~io_in[2];
	assign _015_ = ~(io_in[1] | io_in[2]);
	assign _181_[0] = ~\mchip.counter [0];
	assign _134_ = \mchip.counter [3] | ~\mchip.counter [2];
	assign _135_ = \mchip.counter [0] | \mchip.counter [1];
	assign _136_ = _135_ | _134_;
	assign _137_ = ~(_136_ | _132_);
	assign _000_ = ~(_137_ & \mchip.counter [8]);
	assign _001_ = ~\mchip.new_clock ;
	assign _011_ = ~(io_in[0] | \mchip.PLL.dig_osc.ctr [7]);
	assign _010_ = io_in[0] & \mchip.PLL.dig_osc.ctr [7];
	assign \mchip.PLL.dig_osc.out_of_phase  = ~_108_;
	assign _138_ = _073_ ^ \mchip.PLL.loop_fil.phase_corr [0];
	assign _002_ = (_108_ ? _073_ : _138_);
	assign _139_ = ~(_074_ ^ _072_);
	assign _003_ = (_108_ ? _071_ : _139_);
	assign _140_ = ~(_089_ ^ _077_);
	assign _004_ = (_108_ ? _088_ : _140_);
	assign _141_ = _077_ & ~_089_;
	assign _142_ = _093_ & ~_141_;
	assign _143_ = _142_ ^ _085_;
	assign _005_ = (_108_ ? _084_ : _143_);
	assign _144_ = ~(_097_ ^ _096_);
	assign _006_ = (_108_ ? _062_ : _144_);
	assign _145_ = _097_ | ~_096_;
	assign _146_ = _145_ & ~_063_;
	assign _147_ = _146_ ^ _064_;
	assign _007_ = (_108_ ? _058_ : _147_);
	always @(posedge \mchip.new_clock )
		if (!io_in[13])
			\mchip.PLL.dig_osc.ctr [0] <= 1'h0;
		else
			\mchip.PLL.dig_osc.ctr [0] <= _002_;
	always @(posedge \mchip.new_clock )
		if (!io_in[13])
			\mchip.PLL.dig_osc.ctr [1] <= 1'h0;
		else
			\mchip.PLL.dig_osc.ctr [1] <= _003_;
	always @(posedge \mchip.new_clock )
		if (!io_in[13])
			\mchip.PLL.dig_osc.ctr [2] <= 1'h0;
		else
			\mchip.PLL.dig_osc.ctr [2] <= _004_;
	always @(posedge \mchip.new_clock )
		if (!io_in[13])
			\mchip.PLL.dig_osc.ctr [3] <= 1'h0;
		else
			\mchip.PLL.dig_osc.ctr [3] <= _005_;
	always @(posedge \mchip.new_clock )
		if (!io_in[13])
			\mchip.PLL.dig_osc.ctr [4] <= 1'h0;
		else
			\mchip.PLL.dig_osc.ctr [4] <= _006_;
	always @(posedge \mchip.new_clock )
		if (!io_in[13])
			\mchip.PLL.dig_osc.ctr [5] <= 1'h0;
		else
			\mchip.PLL.dig_osc.ctr [5] <= _007_;
	always @(posedge \mchip.new_clock )
		if (!io_in[13])
			\mchip.PLL.dig_osc.ctr [6] <= 1'h0;
		else
			\mchip.PLL.dig_osc.ctr [6] <= _008_;
	always @(posedge \mchip.new_clock )
		if (!io_in[13])
			\mchip.PLL.dig_osc.ctr [7] <= 1'h0;
		else
			\mchip.PLL.dig_osc.ctr [7] <= _009_;
	always @(posedge \mchip.new_clock )
		if (_010_)
			\mchip.PLL.phase_det.matched  <= 1'h1;
		else if (_011_)
			\mchip.PLL.phase_det.matched  <= 1'h0;
	always @(posedge io_in[12])
		if (!_000_)
			\mchip.counter [0] <= 1'h0;
		else
			\mchip.counter [0] <= _181_[0];
	always @(posedge io_in[12])
		if (!_000_)
			\mchip.counter [1] <= 1'h0;
		else
			\mchip.counter [1] <= _182_[1];
	always @(posedge io_in[12])
		if (!_000_)
			\mchip.counter [2] <= 1'h0;
		else
			\mchip.counter [2] <= _182_[2];
	always @(posedge io_in[12])
		if (!_000_)
			\mchip.counter [3] <= 1'h0;
		else
			\mchip.counter [3] <= _182_[3];
	always @(posedge io_in[12])
		if (!_000_)
			\mchip.counter [4] <= 1'h0;
		else
			\mchip.counter [4] <= _182_[4];
	always @(posedge io_in[12])
		if (!_000_)
			\mchip.counter [5] <= 1'h0;
		else
			\mchip.counter [5] <= _182_[5];
	always @(posedge io_in[12])
		if (!_000_)
			\mchip.counter [6] <= 1'h0;
		else
			\mchip.counter [6] <= _182_[6];
	always @(posedge io_in[12])
		if (!_000_)
			\mchip.counter [7] <= 1'h0;
		else
			\mchip.counter [7] <= _182_[7];
	always @(posedge io_in[12])
		if (!_000_)
			\mchip.counter [8] <= 1'h0;
		else
			\mchip.counter [8] <= _182_[8];
	always @(posedge io_in[12])
		if (!_000_)
			\mchip.new_clock  <= _001_;
	always @(posedge \mchip.new_clock )
		if (io_in[3])
			\mchip.PLL.loop_fil.phase_corr [7] <= 1'h0;
		else
			\mchip.PLL.loop_fil.phase_corr [7] <= _015_;
	always @(posedge \mchip.new_clock )
		if (!io_in[3])
			\mchip.PLL.loop_fil.phase_corr [0] <= 1'h0;
		else
			\mchip.PLL.loop_fil.phase_corr [0] <= _012_;
	always @(posedge \mchip.new_clock )
		if (!io_in[3])
			\mchip.PLL.loop_fil.phase_corr [1] <= 1'h0;
		else
			\mchip.PLL.loop_fil.phase_corr [1] <= _013_;
	always @(posedge \mchip.new_clock )
		if (!io_in[3])
			\mchip.PLL.loop_fil.phase_corr [2] <= 1'h0;
		else
			\mchip.PLL.loop_fil.phase_corr [2] <= _014_;
	always @(posedge \mchip.new_clock )
		if (!io_in[3])
			\mchip.PLL.loop_fil.phase_corr [3] <= 1'h0;
		else
			\mchip.PLL.loop_fil.phase_corr [3] <= _015_;
	always @(posedge \mchip.new_clock )
		if (io_in[3])
			\mchip.PLL.loop_fil.phase_corr [4] <= 1'h0;
		else
			\mchip.PLL.loop_fil.phase_corr [4] <= _012_;
	always @(posedge \mchip.new_clock )
		if (io_in[3])
			\mchip.PLL.loop_fil.phase_corr [5] <= 1'h0;
		else
			\mchip.PLL.loop_fil.phase_corr [5] <= _013_;
	always @(posedge \mchip.new_clock )
		if (io_in[3])
			\mchip.PLL.loop_fil.phase_corr [6] <= 1'h0;
		else
			\mchip.PLL.loop_fil.phase_corr [6] <= _014_;
	assign _181_[8:1] = \mchip.counter [8:1];
	assign _182_[0] = _181_[0];
	assign io_out = {11'h000, \mchip.PLL.dig_osc.out_of_phase , \mchip.PLL.dig_osc.lead_or_lag , \mchip.PLL.dig_osc.ctr [7]};
	assign \mchip.PLL.dig_osc.freq_step  = io_in[11:4];
	assign \mchip.PLL.dig_osc.i_sys_clk  = \mchip.new_clock ;
	assign \mchip.PLL.dig_osc.phase_corr  = \mchip.PLL.loop_fil.phase_corr ;
	assign \mchip.PLL.dig_osc.rec_clk  = \mchip.PLL.dig_osc.ctr [7];
	assign \mchip.PLL.i_freq_step  = io_in[11:4];
	assign \mchip.PLL.i_loop_gain  = io_in[3:1];
	assign \mchip.PLL.i_ref_clk  = io_in[0];
	assign \mchip.PLL.i_sys_clk  = \mchip.new_clock ;
	assign \mchip.PLL.lead_or_lag  = \mchip.PLL.dig_osc.lead_or_lag ;
	assign \mchip.PLL.loop_fil.i_sys_clk  = \mchip.new_clock ;
	assign \mchip.PLL.loop_fil.loop_gain  = io_in[3:1];
	assign \mchip.PLL.o_lead_or_lag  = \mchip.PLL.dig_osc.lead_or_lag ;
	assign \mchip.PLL.o_phase_error  = \mchip.PLL.dig_osc.out_of_phase ;
	assign \mchip.PLL.o_rec_clk  = \mchip.PLL.dig_osc.ctr [7];
	assign \mchip.PLL.out_of_phase  = \mchip.PLL.dig_osc.out_of_phase ;
	assign \mchip.PLL.phase_corr  = \mchip.PLL.loop_fil.phase_corr ;
	assign \mchip.PLL.phase_det.i_sys_clk  = \mchip.new_clock ;
	assign \mchip.PLL.phase_det.lead_or_lag  = \mchip.PLL.dig_osc.lead_or_lag ;
	assign \mchip.PLL.phase_det.out_of_phase  = \mchip.PLL.dig_osc.out_of_phase ;
	assign \mchip.PLL.phase_det.rec_clk  = \mchip.PLL.dig_osc.ctr [7];
	assign \mchip.PLL.phase_det.ref_clk  = io_in[0];
	assign \mchip.clock  = io_in[12];
	assign \mchip.io_in  = io_in[11:0];
	assign \mchip.io_out  = {9'h000, \mchip.PLL.dig_osc.out_of_phase , \mchip.PLL.dig_osc.lead_or_lag , \mchip.PLL.dig_osc.ctr [7]};
	assign \mchip.reset  = io_in[13];
endmodule
module d17_njayawar_tetris (
	io_in,
	io_out
);
	wire _0000_;
	wire _0001_;
	wire _0002_;
	wire _0003_;
	wire _0004_;
	wire _0005_;
	wire _0006_;
	wire _0007_;
	wire _0008_;
	wire _0009_;
	wire _0010_;
	wire _0011_;
	wire _0012_;
	wire _0013_;
	wire _0014_;
	wire _0015_;
	wire _0016_;
	wire _0017_;
	wire _0018_;
	wire _0019_;
	wire _0020_;
	wire _0021_;
	wire _0022_;
	wire _0023_;
	wire _0024_;
	wire _0025_;
	wire _0026_;
	wire _0027_;
	wire _0028_;
	wire _0029_;
	wire _0030_;
	wire _0031_;
	wire _0032_;
	wire _0033_;
	wire _0034_;
	wire _0035_;
	wire _0036_;
	wire _0037_;
	wire _0038_;
	wire _0039_;
	wire _0040_;
	wire _0041_;
	wire _0042_;
	wire _0043_;
	wire _0044_;
	wire _0045_;
	wire _0046_;
	wire _0047_;
	wire _0048_;
	wire _0049_;
	wire _0050_;
	wire _0051_;
	wire _0052_;
	wire _0053_;
	wire _0054_;
	wire _0055_;
	wire _0056_;
	wire _0057_;
	wire _0058_;
	wire _0059_;
	wire _0060_;
	wire _0061_;
	wire _0062_;
	wire _0063_;
	wire _0064_;
	wire _0065_;
	wire _0066_;
	wire _0067_;
	wire _0068_;
	wire _0069_;
	wire _0070_;
	wire _0071_;
	wire _0072_;
	wire _0073_;
	wire _0074_;
	wire _0075_;
	wire _0076_;
	wire _0077_;
	wire _0078_;
	wire _0079_;
	wire _0080_;
	wire _0081_;
	wire _0082_;
	wire _0083_;
	wire _0084_;
	wire _0085_;
	wire _0086_;
	wire _0087_;
	wire _0088_;
	wire _0089_;
	wire _0090_;
	wire _0091_;
	wire _0092_;
	wire _0093_;
	wire _0094_;
	wire _0095_;
	wire _0096_;
	wire _0097_;
	wire _0098_;
	wire _0099_;
	wire _0100_;
	wire _0101_;
	wire _0102_;
	wire _0103_;
	wire _0104_;
	wire _0105_;
	wire _0106_;
	wire _0107_;
	wire _0108_;
	wire _0109_;
	wire _0110_;
	wire _0111_;
	wire _0112_;
	wire _0113_;
	wire _0114_;
	wire _0115_;
	wire _0116_;
	wire _0117_;
	wire _0118_;
	wire _0119_;
	wire _0120_;
	wire _0121_;
	wire _0122_;
	wire _0123_;
	wire _0124_;
	wire _0125_;
	wire _0126_;
	wire _0127_;
	wire _0128_;
	wire _0129_;
	wire _0130_;
	wire _0131_;
	wire _0132_;
	wire _0133_;
	wire _0134_;
	wire _0135_;
	wire _0136_;
	wire _0137_;
	wire _0138_;
	wire _0139_;
	wire _0140_;
	wire _0141_;
	wire _0142_;
	wire _0143_;
	wire _0144_;
	wire _0145_;
	wire _0146_;
	wire _0147_;
	wire _0148_;
	wire _0149_;
	wire _0150_;
	wire _0151_;
	wire _0152_;
	wire _0153_;
	wire _0154_;
	wire _0155_;
	wire _0156_;
	wire _0157_;
	wire _0158_;
	wire _0159_;
	wire _0160_;
	wire _0161_;
	wire _0162_;
	wire _0163_;
	wire _0164_;
	wire _0165_;
	wire _0166_;
	wire _0167_;
	wire _0168_;
	wire _0169_;
	wire _0170_;
	wire _0171_;
	wire _0172_;
	wire _0173_;
	wire _0174_;
	wire _0175_;
	wire _0176_;
	wire _0177_;
	wire _0178_;
	wire _0179_;
	wire _0180_;
	wire _0181_;
	wire _0182_;
	wire _0183_;
	wire _0184_;
	wire _0185_;
	wire _0186_;
	wire _0187_;
	wire _0188_;
	wire _0189_;
	wire _0190_;
	wire _0191_;
	wire _0192_;
	wire _0193_;
	wire _0194_;
	wire _0195_;
	wire _0196_;
	wire _0197_;
	wire _0198_;
	wire _0199_;
	wire _0200_;
	wire _0201_;
	wire _0202_;
	wire _0203_;
	wire _0204_;
	wire _0205_;
	wire _0206_;
	wire _0207_;
	wire _0208_;
	wire _0209_;
	wire _0210_;
	wire _0211_;
	wire _0212_;
	wire _0213_;
	wire _0214_;
	wire _0215_;
	wire _0216_;
	wire _0217_;
	wire _0218_;
	wire _0219_;
	wire _0220_;
	wire _0221_;
	wire _0222_;
	wire _0223_;
	wire _0224_;
	wire _0225_;
	wire _0226_;
	wire _0227_;
	wire _0228_;
	wire _0229_;
	wire _0230_;
	wire _0231_;
	wire _0232_;
	wire _0233_;
	wire _0234_;
	wire _0235_;
	wire _0236_;
	wire _0237_;
	wire _0238_;
	wire _0239_;
	wire _0240_;
	wire _0241_;
	wire _0242_;
	wire _0243_;
	wire _0244_;
	wire _0245_;
	wire _0246_;
	wire _0247_;
	wire _0248_;
	wire _0249_;
	wire _0250_;
	wire _0251_;
	wire _0252_;
	wire _0253_;
	wire _0254_;
	wire _0255_;
	wire _0256_;
	wire _0257_;
	wire _0258_;
	wire _0259_;
	wire _0260_;
	wire _0261_;
	wire _0262_;
	wire _0263_;
	wire _0264_;
	wire _0265_;
	wire _0266_;
	wire _0267_;
	wire _0268_;
	wire _0269_;
	wire _0270_;
	wire _0271_;
	wire _0272_;
	wire _0273_;
	wire _0274_;
	wire _0275_;
	wire _0276_;
	wire _0277_;
	wire _0278_;
	wire _0279_;
	wire _0280_;
	wire _0281_;
	wire _0282_;
	wire _0283_;
	wire _0284_;
	wire _0285_;
	wire _0286_;
	wire _0287_;
	wire _0288_;
	wire _0289_;
	wire _0290_;
	wire _0291_;
	wire _0292_;
	wire _0293_;
	wire _0294_;
	wire _0295_;
	wire _0296_;
	wire _0297_;
	wire _0298_;
	wire _0299_;
	wire _0300_;
	wire _0301_;
	wire _0302_;
	wire _0303_;
	wire _0304_;
	wire _0305_;
	wire _0306_;
	wire _0307_;
	wire _0308_;
	wire _0309_;
	wire _0310_;
	wire _0311_;
	wire _0312_;
	wire _0313_;
	wire _0314_;
	wire _0315_;
	wire _0316_;
	wire _0317_;
	wire _0318_;
	wire _0319_;
	wire _0320_;
	wire _0321_;
	wire _0322_;
	wire _0323_;
	wire _0324_;
	wire _0325_;
	wire _0326_;
	wire _0327_;
	wire _0328_;
	wire _0329_;
	wire _0330_;
	wire _0331_;
	wire _0332_;
	wire _0333_;
	wire _0334_;
	wire _0335_;
	wire _0336_;
	wire _0337_;
	wire _0338_;
	wire _0339_;
	wire _0340_;
	wire _0341_;
	wire _0342_;
	wire _0343_;
	wire _0344_;
	wire _0345_;
	wire _0346_;
	wire _0347_;
	wire _0348_;
	wire _0349_;
	wire _0350_;
	wire _0351_;
	wire _0352_;
	wire _0353_;
	wire _0354_;
	wire _0355_;
	wire _0356_;
	wire _0357_;
	wire _0358_;
	wire _0359_;
	wire _0360_;
	wire _0361_;
	wire _0362_;
	wire _0363_;
	wire _0364_;
	wire _0365_;
	wire _0366_;
	wire _0367_;
	wire _0368_;
	wire _0369_;
	wire _0370_;
	wire _0371_;
	wire _0372_;
	wire _0373_;
	wire _0374_;
	wire _0375_;
	wire _0376_;
	wire _0377_;
	wire _0378_;
	wire _0379_;
	wire _0380_;
	wire _0381_;
	wire _0382_;
	wire _0383_;
	wire _0384_;
	wire _0385_;
	wire _0386_;
	wire _0387_;
	wire _0388_;
	wire _0389_;
	wire _0390_;
	wire _0391_;
	wire _0392_;
	wire _0393_;
	wire _0394_;
	wire _0395_;
	wire _0396_;
	wire _0397_;
	wire _0398_;
	wire _0399_;
	wire _0400_;
	wire _0401_;
	wire _0402_;
	wire _0403_;
	wire _0404_;
	wire _0405_;
	wire _0406_;
	wire _0407_;
	wire _0408_;
	wire _0409_;
	wire _0410_;
	wire _0411_;
	wire _0412_;
	wire _0413_;
	wire _0414_;
	wire _0415_;
	wire _0416_;
	wire _0417_;
	wire _0418_;
	wire _0419_;
	wire _0420_;
	wire _0421_;
	wire _0422_;
	wire _0423_;
	wire _0424_;
	wire _0425_;
	wire _0426_;
	wire _0427_;
	wire _0428_;
	wire _0429_;
	wire _0430_;
	wire _0431_;
	wire _0432_;
	wire _0433_;
	wire _0434_;
	wire _0435_;
	wire _0436_;
	wire _0437_;
	wire _0438_;
	wire _0439_;
	wire _0440_;
	wire _0441_;
	wire _0442_;
	wire _0443_;
	wire _0444_;
	wire _0445_;
	wire _0446_;
	wire _0447_;
	wire _0448_;
	wire _0449_;
	wire _0450_;
	wire _0451_;
	wire _0452_;
	wire _0453_;
	wire _0454_;
	wire _0455_;
	wire _0456_;
	wire _0457_;
	wire _0458_;
	wire _0459_;
	wire _0460_;
	wire _0461_;
	wire _0462_;
	wire _0463_;
	wire _0464_;
	wire _0465_;
	wire _0466_;
	wire _0467_;
	wire _0468_;
	wire _0469_;
	wire _0470_;
	wire _0471_;
	wire _0472_;
	wire _0473_;
	wire _0474_;
	wire _0475_;
	wire _0476_;
	wire _0477_;
	wire _0478_;
	wire _0479_;
	wire _0480_;
	wire _0481_;
	wire _0482_;
	wire _0483_;
	wire _0484_;
	wire _0485_;
	wire _0486_;
	wire _0487_;
	wire _0488_;
	wire _0489_;
	wire _0490_;
	wire _0491_;
	wire _0492_;
	wire _0493_;
	wire _0494_;
	wire _0495_;
	wire _0496_;
	wire _0497_;
	wire _0498_;
	wire _0499_;
	wire _0500_;
	wire _0501_;
	wire _0502_;
	wire _0503_;
	wire _0504_;
	wire _0505_;
	wire _0506_;
	wire _0507_;
	wire _0508_;
	wire _0509_;
	wire _0510_;
	wire _0511_;
	wire _0512_;
	wire _0513_;
	wire _0514_;
	wire _0515_;
	wire _0516_;
	wire _0517_;
	wire _0518_;
	wire _0519_;
	wire _0520_;
	wire _0521_;
	wire _0522_;
	wire _0523_;
	wire _0524_;
	wire _0525_;
	wire _0526_;
	wire _0527_;
	wire _0528_;
	wire _0529_;
	wire _0530_;
	wire _0531_;
	wire _0532_;
	wire _0533_;
	wire _0534_;
	wire _0535_;
	wire _0536_;
	wire _0537_;
	wire _0538_;
	wire _0539_;
	wire _0540_;
	wire _0541_;
	wire _0542_;
	wire _0543_;
	wire _0544_;
	wire _0545_;
	wire _0546_;
	wire _0547_;
	wire _0548_;
	wire _0549_;
	wire _0550_;
	wire _0551_;
	wire _0552_;
	wire _0553_;
	wire _0554_;
	wire _0555_;
	wire _0556_;
	wire _0557_;
	wire _0558_;
	wire _0559_;
	wire _0560_;
	wire _0561_;
	wire _0562_;
	wire _0563_;
	wire _0564_;
	wire _0565_;
	wire _0566_;
	wire _0567_;
	wire _0568_;
	wire _0569_;
	wire _0570_;
	wire _0571_;
	wire _0572_;
	wire _0573_;
	wire _0574_;
	wire _0575_;
	wire _0576_;
	wire _0577_;
	wire _0578_;
	wire _0579_;
	wire _0580_;
	wire _0581_;
	wire _0582_;
	wire _0583_;
	wire _0584_;
	wire _0585_;
	wire _0586_;
	wire _0587_;
	wire _0588_;
	wire _0589_;
	wire _0590_;
	wire _0591_;
	wire _0592_;
	wire _0593_;
	wire _0594_;
	wire _0595_;
	wire _0596_;
	wire _0597_;
	wire _0598_;
	wire _0599_;
	wire _0600_;
	wire _0601_;
	wire _0602_;
	wire _0603_;
	wire _0604_;
	wire _0605_;
	wire _0606_;
	wire _0607_;
	wire _0608_;
	wire _0609_;
	wire _0610_;
	wire _0611_;
	wire _0612_;
	wire _0613_;
	wire _0614_;
	wire _0615_;
	wire _0616_;
	wire _0617_;
	wire _0618_;
	wire _0619_;
	wire _0620_;
	wire _0621_;
	wire _0622_;
	wire _0623_;
	wire _0624_;
	wire _0625_;
	wire _0626_;
	wire _0627_;
	wire _0628_;
	wire _0629_;
	wire _0630_;
	wire _0631_;
	wire _0632_;
	wire _0633_;
	wire _0634_;
	wire _0635_;
	wire _0636_;
	wire _0637_;
	wire _0638_;
	wire _0639_;
	wire _0640_;
	wire _0641_;
	wire _0642_;
	wire _0643_;
	wire _0644_;
	wire _0645_;
	wire _0646_;
	wire _0647_;
	wire _0648_;
	wire _0649_;
	wire _0650_;
	wire _0651_;
	wire _0652_;
	wire _0653_;
	wire _0654_;
	wire _0655_;
	wire _0656_;
	wire _0657_;
	wire _0658_;
	wire _0659_;
	wire _0660_;
	wire _0661_;
	wire _0662_;
	wire _0663_;
	wire _0664_;
	wire _0665_;
	wire _0666_;
	wire _0667_;
	wire _0668_;
	wire _0669_;
	wire _0670_;
	wire _0671_;
	wire _0672_;
	wire _0673_;
	wire _0674_;
	wire _0675_;
	wire _0676_;
	wire _0677_;
	wire _0678_;
	wire _0679_;
	wire _0680_;
	wire _0681_;
	wire _0682_;
	wire _0683_;
	wire _0684_;
	wire _0685_;
	wire _0686_;
	wire _0687_;
	wire _0688_;
	wire _0689_;
	wire _0690_;
	wire _0691_;
	wire _0692_;
	wire _0693_;
	wire _0694_;
	wire _0695_;
	wire _0696_;
	wire _0697_;
	wire _0698_;
	wire _0699_;
	wire _0700_;
	wire _0701_;
	wire _0702_;
	wire _0703_;
	wire _0704_;
	wire _0705_;
	wire _0706_;
	wire _0707_;
	wire _0708_;
	wire _0709_;
	wire _0710_;
	wire _0711_;
	wire _0712_;
	wire _0713_;
	wire _0714_;
	wire _0715_;
	wire _0716_;
	wire _0717_;
	wire _0718_;
	wire _0719_;
	wire _0720_;
	wire _0721_;
	wire _0722_;
	wire _0723_;
	wire _0724_;
	wire _0725_;
	wire _0726_;
	wire _0727_;
	wire _0728_;
	wire _0729_;
	wire _0730_;
	wire _0731_;
	wire _0732_;
	wire _0733_;
	wire _0734_;
	wire _0735_;
	wire _0736_;
	wire _0737_;
	wire _0738_;
	wire _0739_;
	wire _0740_;
	wire _0741_;
	wire _0742_;
	wire _0743_;
	wire _0744_;
	wire _0745_;
	wire _0746_;
	wire _0747_;
	wire _0748_;
	wire _0749_;
	wire _0750_;
	wire _0751_;
	wire _0752_;
	wire _0753_;
	wire _0754_;
	wire _0755_;
	wire _0756_;
	wire _0757_;
	wire _0758_;
	wire _0759_;
	wire _0760_;
	wire _0761_;
	wire _0762_;
	wire _0763_;
	wire _0764_;
	wire _0765_;
	wire _0766_;
	wire _0767_;
	wire _0768_;
	wire _0769_;
	wire _0770_;
	wire _0771_;
	wire _0772_;
	wire _0773_;
	wire _0774_;
	wire _0775_;
	wire _0776_;
	wire _0777_;
	wire _0778_;
	wire _0779_;
	wire _0780_;
	wire _0781_;
	wire _0782_;
	wire _0783_;
	wire _0784_;
	wire _0785_;
	wire _0786_;
	wire _0787_;
	wire _0788_;
	wire _0789_;
	wire _0790_;
	wire _0791_;
	wire _0792_;
	wire _0793_;
	wire _0794_;
	wire _0795_;
	wire _0796_;
	wire _0797_;
	wire _0798_;
	wire _0799_;
	wire _0800_;
	wire _0801_;
	wire _0802_;
	wire _0803_;
	wire _0804_;
	wire _0805_;
	wire _0806_;
	wire _0807_;
	wire _0808_;
	wire _0809_;
	wire _0810_;
	wire _0811_;
	wire _0812_;
	wire _0813_;
	wire _0814_;
	wire _0815_;
	wire _0816_;
	wire _0817_;
	wire _0818_;
	wire _0819_;
	wire _0820_;
	wire _0821_;
	wire _0822_;
	wire _0823_;
	wire _0824_;
	wire _0825_;
	wire _0826_;
	wire _0827_;
	wire _0828_;
	wire _0829_;
	wire _0830_;
	wire _0831_;
	wire _0832_;
	wire _0833_;
	wire _0834_;
	wire _0835_;
	wire _0836_;
	wire _0837_;
	wire _0838_;
	wire _0839_;
	wire _0840_;
	wire _0841_;
	wire _0842_;
	wire _0843_;
	wire _0844_;
	wire _0845_;
	wire _0846_;
	wire _0847_;
	wire _0848_;
	wire _0849_;
	wire _0850_;
	wire _0851_;
	wire _0852_;
	wire _0853_;
	wire _0854_;
	wire _0855_;
	wire _0856_;
	wire _0857_;
	wire _0858_;
	wire _0859_;
	wire _0860_;
	wire _0861_;
	wire _0862_;
	wire _0863_;
	wire _0864_;
	wire _0865_;
	wire _0866_;
	wire _0867_;
	wire _0868_;
	wire _0869_;
	wire _0870_;
	wire _0871_;
	wire _0872_;
	wire _0873_;
	wire _0874_;
	wire _0875_;
	wire _0876_;
	wire _0877_;
	wire _0878_;
	wire _0879_;
	wire _0880_;
	wire _0881_;
	wire _0882_;
	wire _0883_;
	wire _0884_;
	wire _0885_;
	wire _0886_;
	wire _0887_;
	wire _0888_;
	wire _0889_;
	wire _0890_;
	wire _0891_;
	wire _0892_;
	wire _0893_;
	wire _0894_;
	wire _0895_;
	wire _0896_;
	wire _0897_;
	wire _0898_;
	wire _0899_;
	wire _0900_;
	wire _0901_;
	wire _0902_;
	wire _0903_;
	wire _0904_;
	wire _0905_;
	wire _0906_;
	wire _0907_;
	wire _0908_;
	wire _0909_;
	wire _0910_;
	wire _0911_;
	wire _0912_;
	wire _0913_;
	wire _0914_;
	wire _0915_;
	wire _0916_;
	wire _0917_;
	wire _0918_;
	wire _0919_;
	wire _0920_;
	wire _0921_;
	wire _0922_;
	wire _0923_;
	wire _0924_;
	wire _0925_;
	wire _0926_;
	wire _0927_;
	wire _0928_;
	wire _0929_;
	wire _0930_;
	wire _0931_;
	wire _0932_;
	wire _0933_;
	wire _0934_;
	wire _0935_;
	wire _0936_;
	wire _0937_;
	wire _0938_;
	wire _0939_;
	wire _0940_;
	wire _0941_;
	wire _0942_;
	wire _0943_;
	wire _0944_;
	wire _0945_;
	wire _0946_;
	wire _0947_;
	wire _0948_;
	wire _0949_;
	wire _0950_;
	wire _0951_;
	wire _0952_;
	wire _0953_;
	wire _0954_;
	wire _0955_;
	wire _0956_;
	wire _0957_;
	wire _0958_;
	wire _0959_;
	wire _0960_;
	wire _0961_;
	wire _0962_;
	wire _0963_;
	wire _0964_;
	wire _0965_;
	wire _0966_;
	wire _0967_;
	wire _0968_;
	wire _0969_;
	wire _0970_;
	wire _0971_;
	wire _0972_;
	wire _0973_;
	wire _0974_;
	wire _0975_;
	wire _0976_;
	wire _0977_;
	wire _0978_;
	wire _0979_;
	wire _0980_;
	wire _0981_;
	wire _0982_;
	wire _0983_;
	wire _0984_;
	wire _0985_;
	wire _0986_;
	wire _0987_;
	wire _0988_;
	wire _0989_;
	wire _0990_;
	wire _0991_;
	wire _0992_;
	wire _0993_;
	wire _0994_;
	wire _0995_;
	wire _0996_;
	wire _0997_;
	wire _0998_;
	wire _0999_;
	wire _1000_;
	wire _1001_;
	wire _1002_;
	wire _1003_;
	wire _1004_;
	wire _1005_;
	wire _1006_;
	wire _1007_;
	wire _1008_;
	wire _1009_;
	wire _1010_;
	wire _1011_;
	wire _1012_;
	wire _1013_;
	wire _1014_;
	wire _1015_;
	wire _1016_;
	wire _1017_;
	wire _1018_;
	wire _1019_;
	wire _1020_;
	wire _1021_;
	wire _1022_;
	wire _1023_;
	wire _1024_;
	wire _1025_;
	wire _1026_;
	wire _1027_;
	wire _1028_;
	wire _1029_;
	wire _1030_;
	wire _1031_;
	wire _1032_;
	wire _1033_;
	wire _1034_;
	wire _1035_;
	wire _1036_;
	wire _1037_;
	wire _1038_;
	wire _1039_;
	wire _1040_;
	wire _1041_;
	wire _1042_;
	wire _1043_;
	wire _1044_;
	wire _1045_;
	wire _1046_;
	wire _1047_;
	wire _1048_;
	wire _1049_;
	wire _1050_;
	wire _1051_;
	wire _1052_;
	wire _1053_;
	wire _1054_;
	wire _1055_;
	wire _1056_;
	wire _1057_;
	wire _1058_;
	wire _1059_;
	wire _1060_;
	wire _1061_;
	wire _1062_;
	wire _1063_;
	wire _1064_;
	wire _1065_;
	wire _1066_;
	wire _1067_;
	wire _1068_;
	wire _1069_;
	wire _1070_;
	wire _1071_;
	wire [7:0] _1072_;
	wire [7:0] _1073_;
	wire [31:0] _1074_;
	wire [2:0] _1075_;
	wire [3:0] _1076_;
	wire [3:0] _1077_;
	wire [3:0] _1078_;
	wire [3:0] _1079_;
	wire [3:0] _1080_;
	wire [3:0] _1081_;
	wire [3:0] _1082_;
	wire [3:0] _1083_;
	wire [26:0] _1084_;
	wire [26:0] _1085_;
	wire [26:0] _1086_;
	wire [26:0] _1087_;
	input wire [13:0] io_in;
	output wire [13:0] io_out;
	reg [2:0] \mchip.chip_design.bounce.bounce_pos ;
	wire \mchip.chip_design.bounce.clock ;
	wire \mchip.chip_design.bounce.game_running ;
	wire \mchip.chip_design.bounce.reset ;
	reg \mchip.chip_design.bounce.state ;
	wire [2:0] \mchip.chip_design.bounce_pos ;
	wire \mchip.chip_design.clock ;
	wire \mchip.chip_design.drop_btn ;
	reg \mchip.chip_design.drop_button ;
	reg \mchip.chip_design.drop_int ;
	wire [3:0] \mchip.chip_design.drop_pos[0] ;
	wire [3:0] \mchip.chip_design.drop_pos[1] ;
	wire [3:0] \mchip.chip_design.drop_pos[2] ;
	wire [3:0] \mchip.chip_design.drop_pos[3] ;
	wire [3:0] \mchip.chip_design.drop_pos[4] ;
	wire [3:0] \mchip.chip_design.drop_pos[5] ;
	wire [3:0] \mchip.chip_design.drop_pos[6] ;
	wire [3:0] \mchip.chip_design.drop_pos[7] ;
	wire \mchip.chip_design.game_running ;
	wire \mchip.chip_design.genblk1[0].col.clock ;
	reg [3:0] \mchip.chip_design.genblk1[0].col.drop_pos ;
	wire \mchip.chip_design.genblk1[0].col.nextState ;
	wire \mchip.chip_design.genblk1[0].col.reset ;
	wire \mchip.chip_design.genblk1[0].col.stack_dec ;
	reg [3:0] \mchip.chip_design.genblk1[0].col.stack_pos ;
	reg \mchip.chip_design.genblk1[0].col.state ;
	wire \mchip.chip_design.genblk1[1].col.clock ;
	reg [3:0] \mchip.chip_design.genblk1[1].col.drop_pos ;
	wire \mchip.chip_design.genblk1[1].col.nextState ;
	wire \mchip.chip_design.genblk1[1].col.reset ;
	wire \mchip.chip_design.genblk1[1].col.stack_dec ;
	reg [3:0] \mchip.chip_design.genblk1[1].col.stack_pos ;
	reg \mchip.chip_design.genblk1[1].col.state ;
	wire \mchip.chip_design.genblk1[2].col.clock ;
	reg [3:0] \mchip.chip_design.genblk1[2].col.drop_pos ;
	wire \mchip.chip_design.genblk1[2].col.nextState ;
	wire \mchip.chip_design.genblk1[2].col.reset ;
	wire \mchip.chip_design.genblk1[2].col.stack_dec ;
	reg [3:0] \mchip.chip_design.genblk1[2].col.stack_pos ;
	reg \mchip.chip_design.genblk1[2].col.state ;
	wire \mchip.chip_design.genblk1[3].col.clock ;
	reg [3:0] \mchip.chip_design.genblk1[3].col.drop_pos ;
	wire \mchip.chip_design.genblk1[3].col.nextState ;
	wire \mchip.chip_design.genblk1[3].col.reset ;
	wire \mchip.chip_design.genblk1[3].col.stack_dec ;
	reg [3:0] \mchip.chip_design.genblk1[3].col.stack_pos ;
	reg \mchip.chip_design.genblk1[3].col.state ;
	wire \mchip.chip_design.genblk1[4].col.clock ;
	reg [3:0] \mchip.chip_design.genblk1[4].col.drop_pos ;
	wire \mchip.chip_design.genblk1[4].col.nextState ;
	wire \mchip.chip_design.genblk1[4].col.reset ;
	wire \mchip.chip_design.genblk1[4].col.stack_dec ;
	reg [3:0] \mchip.chip_design.genblk1[4].col.stack_pos ;
	reg \mchip.chip_design.genblk1[4].col.state ;
	wire \mchip.chip_design.genblk1[5].col.clock ;
	reg [3:0] \mchip.chip_design.genblk1[5].col.drop_pos ;
	wire \mchip.chip_design.genblk1[5].col.nextState ;
	wire \mchip.chip_design.genblk1[5].col.reset ;
	wire \mchip.chip_design.genblk1[5].col.stack_dec ;
	reg [3:0] \mchip.chip_design.genblk1[5].col.stack_pos ;
	reg \mchip.chip_design.genblk1[5].col.state ;
	wire \mchip.chip_design.genblk1[6].col.clock ;
	reg [3:0] \mchip.chip_design.genblk1[6].col.drop_pos ;
	wire \mchip.chip_design.genblk1[6].col.nextState ;
	wire \mchip.chip_design.genblk1[6].col.reset ;
	wire \mchip.chip_design.genblk1[6].col.stack_dec ;
	reg [3:0] \mchip.chip_design.genblk1[6].col.stack_pos ;
	reg \mchip.chip_design.genblk1[6].col.state ;
	wire \mchip.chip_design.genblk1[7].col.clock ;
	reg [3:0] \mchip.chip_design.genblk1[7].col.drop_pos ;
	wire \mchip.chip_design.genblk1[7].col.nextState ;
	wire \mchip.chip_design.genblk1[7].col.reset ;
	wire \mchip.chip_design.genblk1[7].col.stack_dec ;
	reg [3:0] \mchip.chip_design.genblk1[7].col.stack_pos ;
	reg \mchip.chip_design.genblk1[7].col.state ;
	wire [5:0] \mchip.chip_design.initial_game_speed ;
	wire [11:0] \mchip.chip_design.inputs ;
	reg \mchip.chip_design.new_game ;
	wire \mchip.chip_design.new_game_btn ;
	reg \mchip.chip_design.new_game_int ;
	wire [11:0] \mchip.chip_design.outputs ;
	reg \mchip.chip_design.prev_drop_button ;
	wire \mchip.chip_design.reset ;
	reg [7:0] \mchip.chip_design.score ;
	wire \mchip.chip_design.stack_dec ;
	wire [3:0] \mchip.chip_design.stack_pos[0] ;
	wire [3:0] \mchip.chip_design.stack_pos[1] ;
	wire [3:0] \mchip.chip_design.stack_pos[2] ;
	wire [3:0] \mchip.chip_design.stack_pos[3] ;
	wire [3:0] \mchip.chip_design.stack_pos[4] ;
	wire [3:0] \mchip.chip_design.stack_pos[5] ;
	wire [3:0] \mchip.chip_design.stack_pos[6] ;
	wire [3:0] \mchip.chip_design.stack_pos[7] ;
	reg [3:0] \mchip.chip_design.state ;
	reg [26:0] \mchip.chip_design.timing.bounce_cnt ;
	wire [26:0] \mchip.chip_design.timing.bounce_max_val ;
	wire \mchip.chip_design.timing.clock ;
	reg [26:0] \mchip.chip_design.timing.drop_cnt ;
	wire [26:0] \mchip.chip_design.timing.drop_max_val ;
	wire [5:0] \mchip.chip_design.timing.initial_game_speed ;
	wire [26:0] \mchip.chip_design.timing.initial_game_speed_base ;
	wire \mchip.chip_design.timing.reset ;
	wire [7:0] \mchip.chip_design.timing.score ;
	wire [26:0] \mchip.chip_design.timing.score_base ;
	wire [3:0] \mchip.chip_design.update_request_location ;
	wire [7:0] \mchip.chip_design.update_value ;
	wire \mchip.clock ;
	wire [11:0] \mchip.io_in ;
	wire [11:0] \mchip.io_out ;
	wire \mchip.reset ;
	assign _1084_[0] = ~\mchip.chip_design.timing.drop_cnt [0];
	assign _1083_[0] = ~\mchip.chip_design.genblk1[7].col.drop_pos [0];
	assign _1082_[0] = ~\mchip.chip_design.genblk1[6].col.drop_pos [0];
	assign _1081_[0] = ~\mchip.chip_design.genblk1[5].col.drop_pos [0];
	assign _1080_[0] = ~\mchip.chip_design.genblk1[4].col.drop_pos [0];
	assign _1079_[0] = ~\mchip.chip_design.genblk1[3].col.drop_pos [0];
	assign _1078_[0] = ~\mchip.chip_design.genblk1[2].col.drop_pos [0];
	assign _1077_[0] = ~\mchip.chip_design.genblk1[1].col.drop_pos [0];
	assign _1076_[0] = ~\mchip.chip_design.genblk1[0].col.drop_pos [0];
	assign _0435_ = ~(\mchip.chip_design.genblk1[1].col.stack_pos [1] | \mchip.chip_design.genblk1[1].col.stack_pos [0]);
	assign _0436_ = \mchip.chip_design.genblk1[1].col.stack_pos [2] | \mchip.chip_design.genblk1[1].col.stack_pos [3];
	assign _0437_ = _0435_ & ~_0436_;
	assign _0438_ = ~(\mchip.chip_design.genblk1[0].col.stack_pos [1] | \mchip.chip_design.genblk1[0].col.stack_pos [0]);
	assign _0439_ = \mchip.chip_design.genblk1[0].col.stack_pos [3] | \mchip.chip_design.genblk1[0].col.stack_pos [2];
	assign _0440_ = _0438_ & ~_0439_;
	assign _0441_ = ~(_0440_ | _0437_);
	assign _0442_ = ~(\mchip.chip_design.genblk1[3].col.stack_pos [1] | \mchip.chip_design.genblk1[3].col.stack_pos [0]);
	assign _0443_ = \mchip.chip_design.genblk1[3].col.stack_pos [3] | \mchip.chip_design.genblk1[3].col.stack_pos [2];
	assign _0444_ = _0442_ & ~_0443_;
	assign _0445_ = ~(\mchip.chip_design.genblk1[2].col.stack_pos [0] | \mchip.chip_design.genblk1[2].col.stack_pos [1]);
	assign _0446_ = \mchip.chip_design.genblk1[2].col.stack_pos [3] | \mchip.chip_design.genblk1[2].col.stack_pos [2];
	assign _0447_ = _0445_ & ~_0446_;
	assign _0448_ = _0447_ | _0444_;
	assign _0449_ = _0441_ & ~_0448_;
	assign _0450_ = ~(\mchip.chip_design.genblk1[7].col.stack_pos [0] | \mchip.chip_design.genblk1[7].col.stack_pos [1]);
	assign _0451_ = \mchip.chip_design.genblk1[7].col.stack_pos [2] | \mchip.chip_design.genblk1[7].col.stack_pos [3];
	assign _0452_ = _0450_ & ~_0451_;
	assign _0453_ = ~(\mchip.chip_design.genblk1[6].col.stack_pos [0] | \mchip.chip_design.genblk1[6].col.stack_pos [1]);
	assign _0454_ = \mchip.chip_design.genblk1[6].col.stack_pos [3] | \mchip.chip_design.genblk1[6].col.stack_pos [2];
	assign _0455_ = _0453_ & ~_0454_;
	assign _0456_ = _0455_ | _0452_;
	assign _0457_ = ~(\mchip.chip_design.genblk1[5].col.stack_pos [0] | \mchip.chip_design.genblk1[5].col.stack_pos [1]);
	assign _0458_ = \mchip.chip_design.genblk1[5].col.stack_pos [3] | \mchip.chip_design.genblk1[5].col.stack_pos [2];
	assign _0459_ = _0457_ & ~_0458_;
	assign _0460_ = ~(\mchip.chip_design.genblk1[4].col.stack_pos [0] | \mchip.chip_design.genblk1[4].col.stack_pos [1]);
	assign _0461_ = \mchip.chip_design.genblk1[4].col.stack_pos [2] | \mchip.chip_design.genblk1[4].col.stack_pos [3];
	assign _0462_ = _0460_ & ~_0461_;
	assign _0463_ = _0462_ | _0459_;
	assign _0464_ = _0463_ | _0456_;
	assign \mchip.chip_design.genblk1[0].col.stack_dec  = _0449_ & ~_0464_;
	assign _0465_ = \mchip.chip_design.prev_drop_button  | ~\mchip.chip_design.drop_button ;
	assign _0466_ = \mchip.chip_design.genblk1[1].col.stack_pos [3] | \mchip.chip_design.genblk1[0].col.stack_pos [3];
	assign _0467_ = _0466_ | \mchip.chip_design.genblk1[2].col.stack_pos [3];
	assign _0468_ = _0467_ | \mchip.chip_design.genblk1[3].col.stack_pos [3];
	assign _0469_ = _0468_ | \mchip.chip_design.genblk1[4].col.stack_pos [3];
	assign _0470_ = _0469_ | \mchip.chip_design.genblk1[5].col.stack_pos [3];
	assign _0471_ = ~(_0470_ | \mchip.chip_design.genblk1[6].col.stack_pos [3]);
	assign _0472_ = _0471_ & ~\mchip.chip_design.genblk1[7].col.stack_pos [3];
	assign _0473_ = _0465_ | ~_0472_;
	assign _0474_ = _0473_ | \mchip.chip_design.new_game ;
	assign _0475_ = ~(_0472_ | \mchip.chip_design.new_game );
	assign _0476_ = _0475_ | io_in[13];
	assign _0477_ = _0476_ | _0474_;
	assign _0478_ = \mchip.chip_design.state [2] & ~_0477_;
	assign _0479_ = ~io_in[13];
	assign _0480_ = ~(\mchip.chip_design.genblk1[1].col.stack_pos [0] ^ \mchip.chip_design.genblk1[1].col.drop_pos [0]);
	assign _0481_ = \mchip.chip_design.genblk1[1].col.stack_pos [1] & \mchip.chip_design.genblk1[1].col.stack_pos [0];
	assign _0482_ = ~(_0481_ | _0435_);
	assign _0483_ = _0482_ ^ \mchip.chip_design.genblk1[1].col.drop_pos [1];
	assign _0484_ = _0483_ | _0480_;
	assign _0485_ = _0481_ & \mchip.chip_design.genblk1[1].col.stack_pos [2];
	assign _0486_ = _0485_ ^ \mchip.chip_design.genblk1[1].col.stack_pos [3];
	assign _0487_ = _0486_ ^ \mchip.chip_design.genblk1[1].col.drop_pos [3];
	assign _0488_ = _0481_ ^ \mchip.chip_design.genblk1[1].col.stack_pos [2];
	assign _0489_ = _0488_ ^ \mchip.chip_design.genblk1[1].col.drop_pos [2];
	assign _0490_ = _0489_ | _0487_;
	assign _0491_ = _0490_ | _0484_;
	assign _0492_ = \mchip.chip_design.genblk1[1].col.state  & ~_0491_;
	assign _0493_ = \mchip.chip_design.genblk1[0].col.stack_pos [1] & \mchip.chip_design.genblk1[0].col.stack_pos [0];
	assign _0494_ = _0493_ & \mchip.chip_design.genblk1[0].col.stack_pos [2];
	assign _0495_ = _0494_ ^ \mchip.chip_design.genblk1[0].col.stack_pos [3];
	assign _0496_ = _0495_ ^ \mchip.chip_design.genblk1[0].col.drop_pos [3];
	assign _0497_ = _0493_ ^ \mchip.chip_design.genblk1[0].col.stack_pos [2];
	assign _0498_ = _0497_ ^ \mchip.chip_design.genblk1[0].col.drop_pos [2];
	assign _0499_ = _0498_ | _0496_;
	assign _0500_ = ~(_0493_ | _0438_);
	assign _0501_ = _0500_ ^ \mchip.chip_design.genblk1[0].col.drop_pos [1];
	assign _0502_ = ~(\mchip.chip_design.genblk1[0].col.stack_pos [0] ^ \mchip.chip_design.genblk1[0].col.drop_pos [0]);
	assign _0503_ = _0502_ | _0501_;
	assign _0504_ = _0503_ | _0499_;
	assign _0505_ = \mchip.chip_design.genblk1[0].col.state  & ~_0504_;
	assign _0506_ = ~(_0505_ | _0492_);
	assign _0507_ = ~(\mchip.chip_design.genblk1[3].col.stack_pos [0] ^ \mchip.chip_design.genblk1[3].col.drop_pos [0]);
	assign _0508_ = \mchip.chip_design.genblk1[3].col.stack_pos [1] & \mchip.chip_design.genblk1[3].col.stack_pos [0];
	assign _0509_ = ~(_0508_ | _0442_);
	assign _0510_ = _0509_ ^ \mchip.chip_design.genblk1[3].col.drop_pos [1];
	assign _0511_ = _0510_ | _0507_;
	assign _0512_ = _0508_ & \mchip.chip_design.genblk1[3].col.stack_pos [2];
	assign _0513_ = _0512_ ^ \mchip.chip_design.genblk1[3].col.stack_pos [3];
	assign _0514_ = _0513_ ^ \mchip.chip_design.genblk1[3].col.drop_pos [3];
	assign _0515_ = _0508_ ^ \mchip.chip_design.genblk1[3].col.stack_pos [2];
	assign _0516_ = _0515_ ^ \mchip.chip_design.genblk1[3].col.drop_pos [2];
	assign _0517_ = _0516_ | _0514_;
	assign _0518_ = _0517_ | _0511_;
	assign _0519_ = \mchip.chip_design.genblk1[3].col.state  & ~_0518_;
	assign _0520_ = ~(\mchip.chip_design.genblk1[2].col.stack_pos [0] ^ \mchip.chip_design.genblk1[2].col.drop_pos [0]);
	assign _0521_ = \mchip.chip_design.genblk1[2].col.stack_pos [0] & \mchip.chip_design.genblk1[2].col.stack_pos [1];
	assign _0522_ = ~(_0521_ | _0445_);
	assign _0523_ = _0522_ ^ \mchip.chip_design.genblk1[2].col.drop_pos [1];
	assign _0524_ = _0523_ | _0520_;
	assign _0525_ = _0521_ & \mchip.chip_design.genblk1[2].col.stack_pos [2];
	assign _0526_ = _0525_ ^ \mchip.chip_design.genblk1[2].col.stack_pos [3];
	assign _0527_ = _0526_ ^ \mchip.chip_design.genblk1[2].col.drop_pos [3];
	assign _0528_ = _0521_ ^ \mchip.chip_design.genblk1[2].col.stack_pos [2];
	assign _0529_ = _0528_ ^ \mchip.chip_design.genblk1[2].col.drop_pos [2];
	assign _0530_ = _0529_ | _0527_;
	assign _0531_ = _0530_ | _0524_;
	assign _0532_ = \mchip.chip_design.genblk1[2].col.state  & ~_0531_;
	assign _0533_ = _0532_ | _0519_;
	assign _0534_ = _0506_ & ~_0533_;
	assign _0535_ = ~(\mchip.chip_design.genblk1[7].col.stack_pos [0] ^ \mchip.chip_design.genblk1[7].col.drop_pos [0]);
	assign _0536_ = \mchip.chip_design.genblk1[7].col.stack_pos [0] & \mchip.chip_design.genblk1[7].col.stack_pos [1];
	assign _0537_ = ~(_0536_ | _0450_);
	assign _0538_ = _0537_ ^ \mchip.chip_design.genblk1[7].col.drop_pos [1];
	assign _0539_ = _0538_ | _0535_;
	assign _0540_ = _0536_ & \mchip.chip_design.genblk1[7].col.stack_pos [2];
	assign _0541_ = _0540_ ^ \mchip.chip_design.genblk1[7].col.stack_pos [3];
	assign _0542_ = _0541_ ^ \mchip.chip_design.genblk1[7].col.drop_pos [3];
	assign _0543_ = _0536_ ^ \mchip.chip_design.genblk1[7].col.stack_pos [2];
	assign _0544_ = _0543_ ^ \mchip.chip_design.genblk1[7].col.drop_pos [2];
	assign _0545_ = _0544_ | _0542_;
	assign _0546_ = _0545_ | _0539_;
	assign _0547_ = \mchip.chip_design.genblk1[7].col.state  & ~_0546_;
	assign _0548_ = ~(\mchip.chip_design.genblk1[6].col.stack_pos [0] ^ \mchip.chip_design.genblk1[6].col.drop_pos [0]);
	assign _0549_ = \mchip.chip_design.genblk1[6].col.stack_pos [0] & \mchip.chip_design.genblk1[6].col.stack_pos [1];
	assign _0550_ = ~(_0549_ | _0453_);
	assign _0551_ = _0550_ ^ \mchip.chip_design.genblk1[6].col.drop_pos [1];
	assign _0552_ = _0551_ | _0548_;
	assign _0553_ = _0549_ & \mchip.chip_design.genblk1[6].col.stack_pos [2];
	assign _0554_ = _0553_ ^ \mchip.chip_design.genblk1[6].col.stack_pos [3];
	assign _0555_ = _0554_ ^ \mchip.chip_design.genblk1[6].col.drop_pos [3];
	assign _0556_ = _0549_ ^ \mchip.chip_design.genblk1[6].col.stack_pos [2];
	assign _0557_ = _0556_ ^ \mchip.chip_design.genblk1[6].col.drop_pos [2];
	assign _0558_ = _0557_ | _0555_;
	assign _0559_ = _0558_ | _0552_;
	assign _0560_ = \mchip.chip_design.genblk1[6].col.state  & ~_0559_;
	assign _0561_ = _0560_ | _0547_;
	assign _0562_ = ~(\mchip.chip_design.genblk1[5].col.stack_pos [0] ^ \mchip.chip_design.genblk1[5].col.drop_pos [0]);
	assign _0563_ = \mchip.chip_design.genblk1[5].col.stack_pos [0] & \mchip.chip_design.genblk1[5].col.stack_pos [1];
	assign _0564_ = ~(_0563_ | _0457_);
	assign _0565_ = _0564_ ^ \mchip.chip_design.genblk1[5].col.drop_pos [1];
	assign _0566_ = _0565_ | _0562_;
	assign _0567_ = _0563_ & \mchip.chip_design.genblk1[5].col.stack_pos [2];
	assign _0568_ = _0567_ ^ \mchip.chip_design.genblk1[5].col.stack_pos [3];
	assign _0569_ = _0568_ ^ \mchip.chip_design.genblk1[5].col.drop_pos [3];
	assign _0570_ = _0563_ ^ \mchip.chip_design.genblk1[5].col.stack_pos [2];
	assign _0571_ = _0570_ ^ \mchip.chip_design.genblk1[5].col.drop_pos [2];
	assign _0572_ = _0571_ | _0569_;
	assign _0573_ = _0572_ | _0566_;
	assign _0574_ = \mchip.chip_design.genblk1[5].col.state  & ~_0573_;
	assign _0575_ = ~(\mchip.chip_design.genblk1[4].col.stack_pos [0] ^ \mchip.chip_design.genblk1[4].col.drop_pos [0]);
	assign _0576_ = \mchip.chip_design.genblk1[4].col.stack_pos [0] & \mchip.chip_design.genblk1[4].col.stack_pos [1];
	assign _0577_ = ~(_0576_ | _0460_);
	assign _0578_ = _0577_ ^ \mchip.chip_design.genblk1[4].col.drop_pos [1];
	assign _0579_ = _0578_ | _0575_;
	assign _0580_ = _0576_ & \mchip.chip_design.genblk1[4].col.stack_pos [2];
	assign _0581_ = _0580_ ^ \mchip.chip_design.genblk1[4].col.stack_pos [3];
	assign _0582_ = _0581_ ^ \mchip.chip_design.genblk1[4].col.drop_pos [3];
	assign _0583_ = _0576_ ^ \mchip.chip_design.genblk1[4].col.stack_pos [2];
	assign _0584_ = _0583_ ^ \mchip.chip_design.genblk1[4].col.drop_pos [2];
	assign _0585_ = _0584_ | _0582_;
	assign _0586_ = _0585_ | _0579_;
	assign _0587_ = \mchip.chip_design.genblk1[4].col.state  & ~_0586_;
	assign _0588_ = _0587_ | _0574_;
	assign _0589_ = _0588_ | _0561_;
	assign _0590_ = _0534_ & ~_0589_;
	assign _0591_ = ~(_0590_ & _0479_);
	assign _0592_ = \mchip.chip_design.state [1] & ~_0591_;
	assign _0001_ = _0592_ | _0478_;
	assign _1086_[0] = ~\mchip.chip_design.timing.bounce_cnt [0];
	assign _0593_ = \mchip.chip_design.new_game  | io_in[13];
	assign _0594_ = \mchip.chip_design.state [0] & ~_0593_;
	assign _0000_ = _0594_ | io_in[13];
	assign _0595_ = ~(\mchip.chip_design.timing.drop_cnt [16] | \mchip.chip_design.timing.drop_cnt [17]);
	assign _0596_ = \mchip.chip_design.timing.drop_cnt [18] | \mchip.chip_design.timing.drop_cnt [19];
	assign _0597_ = _0595_ & ~_0596_;
	assign _0598_ = \mchip.chip_design.timing.drop_cnt [22] | \mchip.chip_design.timing.drop_cnt [23];
	assign _0599_ = \mchip.chip_design.timing.drop_cnt [20] | \mchip.chip_design.timing.drop_cnt [21];
	assign _0600_ = _0599_ | _0598_;
	assign _0601_ = _0597_ & ~_0600_;
	assign _0602_ = \mchip.chip_design.timing.drop_cnt [24] | \mchip.chip_design.timing.drop_cnt [25];
	assign _0603_ = _0602_ | \mchip.chip_design.timing.drop_cnt [26];
	assign _0604_ = _0601_ & ~_0603_;
	assign _0605_ = \mchip.chip_design.timing.drop_cnt [14] | \mchip.chip_design.timing.drop_cnt [15];
	assign _0606_ = \mchip.chip_design.timing.drop_cnt [13] | ~\mchip.chip_design.timing.drop_cnt [12];
	assign _0607_ = _0606_ | _0605_;
	assign _0608_ = \mchip.chip_design.timing.drop_cnt [10] | \mchip.chip_design.timing.drop_cnt [11];
	assign _0609_ = ~(\mchip.chip_design.timing.drop_cnt [8] & \mchip.chip_design.timing.drop_cnt [9]);
	assign _0610_ = _0609_ | _0608_;
	assign _0611_ = _0610_ | _0607_;
	assign _0612_ = \mchip.chip_design.timing.drop_cnt [1] | ~\mchip.chip_design.timing.drop_cnt [0];
	assign _0613_ = \mchip.chip_design.timing.drop_cnt [2] | ~\mchip.chip_design.timing.drop_cnt [3];
	assign _0614_ = _0613_ | _0612_;
	assign _0615_ = \mchip.chip_design.timing.drop_cnt [6] | ~\mchip.chip_design.timing.drop_cnt [7];
	assign _0616_ = \mchip.chip_design.timing.drop_cnt [4] | \mchip.chip_design.timing.drop_cnt [5];
	assign _0617_ = _0616_ | _0615_;
	assign _0618_ = _0617_ | _0614_;
	assign _0619_ = _0618_ | _0611_;
	assign _0620_ = _0604_ & ~_0619_;
	assign _0012_ = _0620_ | io_in[13];
	assign _0621_ = _0590_ | io_in[13];
	assign _0622_ = \mchip.chip_design.state [1] & ~_0621_;
	assign _0623_ = _0476_ | ~_0474_;
	assign _0624_ = \mchip.chip_design.state [2] & ~_0623_;
	assign _0625_ = \mchip.chip_design.new_game  & ~io_in[13];
	assign _0626_ = ~(\mchip.chip_design.state [3] | \mchip.chip_design.state [0]);
	assign _0627_ = _0625_ & ~_0626_;
	assign _0628_ = _0627_ | _0624_;
	assign _0002_ = _0628_ | _0622_;
	assign _0629_ = ~(_0475_ & _0479_);
	assign _0630_ = \mchip.chip_design.state [2] & ~_0629_;
	assign _0631_ = \mchip.chip_design.state [3] & ~_0593_;
	assign _0003_ = _0631_ | _0630_;
	assign _0632_ = ~\mchip.chip_design.score [7];
	assign _0633_ = ~\mchip.chip_design.score [5];
	assign _0634_ = \mchip.chip_design.score [7] & \mchip.chip_design.score [1];
	assign _0635_ = ~(_0634_ & \mchip.chip_design.score [2]);
	assign _0636_ = _0634_ ^ \mchip.chip_design.score [2];
	assign _0637_ = _0636_ & ~_0632_;
	assign _0638_ = _0635_ & ~_0637_;
	assign _0639_ = \mchip.chip_design.score [3] & ~_0638_;
	assign _0640_ = ~(_0639_ & \mchip.chip_design.score [4]);
	assign _0641_ = _0639_ ^ \mchip.chip_design.score [4];
	assign _0642_ = _0641_ & ~_0632_;
	assign _0643_ = _0640_ & ~_0642_;
	assign _0644_ = _0643_ | _0633_;
	assign _0645_ = ~\mchip.chip_design.score [3];
	assign _0646_ = _0638_ ^ _0645_;
	assign _0647_ = _0636_ ^ \mchip.chip_design.score [7];
	assign _0648_ = \mchip.chip_design.score [7] ^ \mchip.chip_design.score [1];
	assign _0649_ = \mchip.chip_design.score [6] & \mchip.chip_design.score [0];
	assign _0650_ = ~(_0649_ & _0648_);
	assign _0651_ = ~\mchip.chip_design.score [6];
	assign _0652_ = _0649_ ^ _0648_;
	assign _0653_ = _0652_ & ~_0651_;
	assign _0654_ = _0650_ & ~_0653_;
	assign _0655_ = _0647_ & ~_0654_;
	assign _0656_ = _0655_ & _0646_;
	assign _0657_ = _0655_ ^ _0646_;
	assign _0658_ = _0657_ & ~_0651_;
	assign _0659_ = ~(_0658_ | _0656_);
	assign _0660_ = _0641_ ^ \mchip.chip_design.score [7];
	assign _0661_ = _0660_ & ~_0659_;
	assign _0662_ = _0643_ ^ _0633_;
	assign _0663_ = _0662_ & _0661_;
	assign _0664_ = _0644_ & ~_0663_;
	assign _0665_ = ~(_0660_ ^ _0659_);
	assign _0666_ = _0665_ & _0662_;
	assign _0667_ = \mchip.chip_design.score [6] ^ \mchip.chip_design.score [0];
	assign _0668_ = _0667_ & ~_0633_;
	assign _0669_ = _0652_ ^ \mchip.chip_design.score [6];
	assign _0670_ = _0669_ & _0668_;
	assign _0671_ = ~(_0654_ ^ _0647_);
	assign _0672_ = ~(_0671_ & _0670_);
	assign _0673_ = _0671_ ^ _0670_;
	assign _0674_ = _0673_ & ~_0633_;
	assign _0675_ = _0672_ & ~_0674_;
	assign _0676_ = _0657_ ^ \mchip.chip_design.score [6];
	assign _0677_ = _0675_ | ~_0676_;
	assign _0678_ = _0669_ ^ _0668_;
	assign _0679_ = \mchip.chip_design.score [5] & \mchip.chip_design.score [4];
	assign _0680_ = ~_0679_;
	assign _0681_ = _0667_ ^ \mchip.chip_design.score [5];
	assign _0682_ = _0681_ & ~_0680_;
	assign _0683_ = _0682_ & _0678_;
	assign _0684_ = ~\mchip.chip_design.score [4];
	assign _0685_ = _0682_ ^ _0678_;
	assign _0686_ = _0685_ & ~_0684_;
	assign _0687_ = ~(_0686_ | _0683_);
	assign _0688_ = _0673_ ^ \mchip.chip_design.score [5];
	assign _0689_ = _0688_ & ~_0687_;
	assign _0690_ = _0676_ ^ _0675_;
	assign _0691_ = _0689_ & ~_0690_;
	assign _0692_ = _0677_ & ~_0691_;
	assign _0693_ = _0666_ & ~_0692_;
	assign _0694_ = _0664_ & ~_0693_;
	assign _0695_ = _0688_ ^ _0687_;
	assign _0696_ = ~(_0695_ | _0690_);
	assign _0697_ = _0696_ & _0666_;
	assign _0698_ = _0681_ ^ _0680_;
	assign _0699_ = \mchip.chip_design.score [4] & \mchip.chip_design.score [3];
	assign _0700_ = \mchip.chip_design.score [5] ^ \mchip.chip_design.score [4];
	assign _0701_ = _0700_ & _0699_;
	assign _0702_ = _0701_ & ~_0698_;
	assign _0703_ = _0701_ ^ _0698_;
	assign _0704_ = \mchip.chip_design.score [3] & ~_0703_;
	assign _0705_ = _0704_ | _0702_;
	assign _0706_ = _0685_ ^ \mchip.chip_design.score [4];
	assign _0707_ = ~(_0706_ & _0705_);
	assign _0708_ = _0700_ ^ _0699_;
	assign _0709_ = ~(\mchip.chip_design.score [3] & \mchip.chip_design.score [2]);
	assign _0710_ = \mchip.chip_design.score [4] ^ \mchip.chip_design.score [3];
	assign _0711_ = _0710_ & ~_0709_;
	assign _0712_ = _0711_ & _0708_;
	assign _0713_ = ~\mchip.chip_design.score [2];
	assign _0714_ = _0711_ ^ _0708_;
	assign _0715_ = _0714_ & ~_0713_;
	assign _0716_ = ~(_0715_ | _0712_);
	assign _0717_ = _0703_ ^ _0645_;
	assign _0718_ = _0717_ & ~_0716_;
	assign _0719_ = _0706_ ^ _0705_;
	assign _0720_ = _0719_ & _0718_;
	assign _0721_ = _0707_ & ~_0720_;
	assign _0722_ = ~(_0717_ ^ _0716_);
	assign _0723_ = ~_0722_;
	assign _0724_ = _0719_ & ~_0723_;
	assign _0725_ = _0710_ ^ _0709_;
	assign _0726_ = \mchip.chip_design.score [2] & \mchip.chip_design.score [1];
	assign _0727_ = ~(\mchip.chip_design.score [3] ^ \mchip.chip_design.score [2]);
	assign _0728_ = _0726_ & ~_0727_;
	assign _0729_ = _0728_ & ~_0725_;
	assign _0730_ = _0728_ ^ _0725_;
	assign _0731_ = \mchip.chip_design.score [1] & ~_0730_;
	assign _0732_ = ~(_0731_ | _0729_);
	assign _0733_ = _0714_ ^ \mchip.chip_design.score [2];
	assign _0734_ = _0732_ | ~_0733_;
	assign _0735_ = _0730_ ^ \mchip.chip_design.score [1];
	assign _0736_ = _0727_ ^ _0726_;
	assign _0737_ = \mchip.chip_design.score [1] & \mchip.chip_design.score [0];
	assign _0738_ = ~(\mchip.chip_design.score [2] ^ \mchip.chip_design.score [1]);
	assign _0739_ = _0737_ & ~_0738_;
	assign _0740_ = _0736_ | ~_0739_;
	assign _0741_ = _0739_ ^ _0736_;
	assign _0742_ = \mchip.chip_design.score [0] & ~_0741_;
	assign _0743_ = _0740_ & ~_0742_;
	assign _0744_ = ~(_0743_ | _0735_);
	assign _0745_ = _0733_ ^ _0732_;
	assign _0746_ = _0744_ & ~_0745_;
	assign _0747_ = _0734_ & ~_0746_;
	assign _0748_ = _0724_ & ~_0747_;
	assign _0749_ = _0721_ & ~_0748_;
	assign _0750_ = _0697_ & ~_0749_;
	assign _0751_ = _0694_ & ~_0750_;
	assign _0752_ = \mchip.chip_design.score [6] & ~_0751_;
	assign _0753_ = _0752_ ^ _0632_;
	assign _0754_ = io_in[10] ^ io_in[9];
	assign _0755_ = ~(_0754_ & io_in[7]);
	assign _0756_ = io_in[11] ^ io_in[8];
	assign _0757_ = _0756_ ^ io_in[10];
	assign _0758_ = _0755_ | ~_0757_;
	assign _0759_ = io_in[10] & io_in[9];
	assign _0760_ = _0757_ ^ _0755_;
	assign _0761_ = _0759_ & ~_0760_;
	assign _0762_ = _0758_ & ~_0761_;
	assign _0763_ = ~io_in[10];
	assign _0764_ = _0756_ & ~_0763_;
	assign _0765_ = io_in[11] & ~io_in[8];
	assign _0766_ = io_in[9] ^ io_in[6];
	assign _0767_ = _0766_ ^ _0765_;
	assign _0768_ = _0767_ ^ _0764_;
	assign _0769_ = _0768_ & ~_0762_;
	assign _0770_ = ~(io_in[8] & io_in[7]);
	assign _0771_ = io_in[7] | ~io_in[8];
	assign _0772_ = _0766_ & ~_0771_;
	assign _0773_ = _0770_ & ~_0772_;
	assign _0774_ = _0754_ ^ io_in[7];
	assign _0775_ = _0773_ | ~_0774_;
	assign _0776_ = io_in[9] & io_in[6];
	assign _0777_ = _0774_ ^ _0773_;
	assign _0778_ = _0776_ & ~_0777_;
	assign _0779_ = _0778_ | ~_0775_;
	assign _0780_ = _0760_ ^ _0759_;
	assign _0781_ = _0779_ & ~_0780_;
	assign _0782_ = _0780_ ^ _0779_;
	assign _0783_ = _0777_ ^ _0776_;
	assign _0784_ = _0783_ | _0782_;
	assign _0785_ = io_in[7] & io_in[6];
	assign _0786_ = io_in[8] ^ io_in[7];
	assign _0787_ = _0786_ & _0785_;
	assign _0788_ = ~(_0771_ ^ _0766_);
	assign _0789_ = _0788_ & _0787_;
	assign _0790_ = _0789_ & ~_0784_;
	assign _0791_ = _0790_ | _0781_;
	assign _0792_ = _0768_ ^ _0762_;
	assign _0793_ = _0791_ & ~_0792_;
	assign _0794_ = ~(_0793_ | _0769_);
	assign _0795_ = ~(_0767_ & _0764_);
	assign _0796_ = ~(io_in[11] & io_in[8]);
	assign _0797_ = _0766_ & _0765_;
	assign _0798_ = _0796_ & ~_0797_;
	assign _0799_ = ~(io_in[10] ^ io_in[7]);
	assign _0800_ = _0799_ ^ _0798_;
	assign _0801_ = ~(_0800_ ^ _0776_);
	assign _0802_ = ~(_0801_ ^ _0795_);
	assign _0803_ = _0802_ ^ _0794_;
	assign _0804_ = ~(_0792_ ^ _0791_);
	assign _0805_ = _0803_ & ~_0804_;
	assign _0806_ = _0789_ & ~_0783_;
	assign _0807_ = ~(_0806_ ^ _0782_);
	assign _0808_ = ~(_0789_ ^ _0783_);
	assign _0809_ = _0808_ | _0807_;
	assign _0810_ = _0805_ & ~_0809_;
	assign _0811_ = _0788_ ^ _0787_;
	assign _0812_ = ~(io_in[7] | io_in[6]);
	assign _0813_ = _0786_ ^ _0785_;
	assign _0814_ = _0813_ | ~_0811_;
	assign _0815_ = _0812_ & ~_0814_;
	assign _0816_ = _0811_ & ~_0815_;
	assign _0817_ = _0810_ & ~_0816_;
	assign _0818_ = _0803_ & ~_0817_;
	assign _0819_ = io_in[10] & io_in[7];
	assign _0820_ = _0819_ & _0756_;
	assign _0821_ = ~(_0796_ ^ io_in[9]);
	assign _0822_ = _0821_ & _0820_;
	assign _0823_ = _0821_ ^ _0820_;
	assign _0824_ = _0799_ | _0798_;
	assign _0825_ = _0800_ & _0776_;
	assign _0826_ = _0824_ & ~_0825_;
	assign _0827_ = _0819_ ^ _0756_;
	assign _0828_ = _0826_ | ~_0827_;
	assign _0829_ = _0823_ & ~_0828_;
	assign _0830_ = _0829_ | _0822_;
	assign _0831_ = _0827_ ^ _0826_;
	assign _0832_ = _0823_ & ~_0831_;
	assign _0833_ = _0801_ | _0795_;
	assign _0834_ = _0769_ & ~_0802_;
	assign _0835_ = _0833_ & ~_0834_;
	assign _0836_ = _0802_ | _0792_;
	assign _0837_ = _0781_ & ~_0836_;
	assign _0838_ = _0835_ & ~_0837_;
	assign _0839_ = _0836_ | _0784_;
	assign _0840_ = _0789_ & ~_0839_;
	assign _0841_ = _0838_ & ~_0840_;
	assign _0842_ = _0832_ & ~_0841_;
	assign _0843_ = ~(_0842_ | _0830_);
	assign _0844_ = io_in[9] & ~_0796_;
	assign _0845_ = _0844_ ^ _0763_;
	assign _0846_ = _0845_ | _0843_;
	assign _0847_ = _0844_ & ~_0763_;
	assign _0848_ = _0847_ ^ io_in[11];
	assign _0849_ = _0848_ ^ _0846_;
	assign _0850_ = ~(_0845_ ^ _0843_);
	assign _0851_ = _0850_ & _0849_;
	assign _0852_ = ~(_0841_ | _0831_);
	assign _0853_ = _0828_ & ~_0852_;
	assign _0854_ = _0853_ ^ _0823_;
	assign _0855_ = ~(_0841_ ^ _0831_);
	assign _0856_ = ~(_0855_ | _0854_);
	assign _0857_ = ~(_0856_ & _0851_);
	assign _0858_ = _0857_ | _0818_;
	assign _0859_ = _0851_ & ~_0856_;
	assign _0860_ = _0859_ | ~_0858_;
	assign _0861_ = ~(_0847_ & io_in[11]);
	assign _0862_ = _0845_ | ~_0848_;
	assign _0863_ = _0830_ & ~_0862_;
	assign _0864_ = _0861_ & ~_0863_;
	assign _0865_ = _0862_ | ~_0832_;
	assign _0866_ = ~(_0865_ | _0841_);
	assign _0867_ = _0864_ & ~_0866_;
	assign _0868_ = ~(_0867_ ^ _0860_);
	assign _0869_ = _0868_ ^ _0753_;
	assign _0870_ = _0751_ ^ _0651_;
	assign _0871_ = _0856_ & _0818_;
	assign _0872_ = _0850_ & ~_0871_;
	assign _0873_ = _0872_ ^ _0849_;
	assign _0874_ = ~(_0873_ ^ _0870_);
	assign _0875_ = ~(_0874_ & _0869_);
	assign _0876_ = _0747_ | _0723_;
	assign _0877_ = _0718_ | ~_0876_;
	assign _0878_ = _0877_ ^ _0719_;
	assign _0879_ = ~(_0816_ | _0809_);
	assign _0880_ = ~(_0879_ ^ _0804_);
	assign _0881_ = _0880_ & ~_0878_;
	assign _0882_ = ~(_0816_ | _0808_);
	assign _0883_ = ~(_0882_ ^ _0807_);
	assign _0884_ = _0747_ ^ _0723_;
	assign _0885_ = _0883_ & ~_0884_;
	assign _0886_ = ~_0885_;
	assign _0887_ = ~(_0880_ ^ _0878_);
	assign _0888_ = _0887_ & ~_0886_;
	assign _0889_ = ~(_0888_ | _0881_);
	assign _0890_ = ~(_0884_ ^ _0883_);
	assign _0891_ = _0890_ & _0887_;
	assign _0892_ = ~(_0745_ ^ _0744_);
	assign _0893_ = _0816_ ^ _0808_;
	assign _0894_ = _0892_ | ~_0893_;
	assign _0895_ = _0812_ & ~_0813_;
	assign _0896_ = _0895_ ^ _0811_;
	assign _0897_ = _0743_ ^ _0735_;
	assign _0898_ = _0896_ & ~_0897_;
	assign _0899_ = ~_0898_;
	assign _0900_ = ~(_0893_ ^ _0892_);
	assign _0901_ = _0900_ & ~_0899_;
	assign _0902_ = _0894_ & ~_0901_;
	assign _0903_ = _0891_ & ~_0902_;
	assign _0904_ = _0889_ & ~_0903_;
	assign _1072_[0] = ~\mchip.chip_design.score [0];
	assign _0905_ = _0741_ ^ _1072_[0];
	assign _0906_ = ~(_0813_ ^ _0812_);
	assign _0907_ = _0906_ & ~_0905_;
	assign _0908_ = ~(_0812_ | _0785_);
	assign _0909_ = _0908_ ^ io_in[6];
	assign _0910_ = ~(_0738_ ^ _0737_);
	assign _0911_ = _0909_ & ~_0910_;
	assign _0912_ = ~_0911_;
	assign _0913_ = ~(_0906_ ^ _0905_);
	assign _0914_ = _0913_ & ~_0912_;
	assign _0915_ = ~(_0914_ | _0907_);
	assign _0916_ = (\mchip.chip_design.score [1] ? io_in[6] : _1072_[0]);
	assign _0917_ = ~(_0910_ ^ _0909_);
	assign _0918_ = ~(_0917_ & _0913_);
	assign _0919_ = _0916_ & ~_0918_;
	assign _0920_ = _0915_ & ~_0919_;
	assign _0921_ = ~_0920_;
	assign _0922_ = ~(_0897_ ^ _0896_);
	assign _0923_ = ~(_0922_ & _0900_);
	assign _0924_ = _0923_ | ~_0891_;
	assign _0925_ = _0921_ & ~_0924_;
	assign _0926_ = _0904_ & ~_0925_;
	assign _0927_ = ~_0926_;
	assign _0928_ = ~_0665_;
	assign _0929_ = _0696_ & ~_0749_;
	assign _0930_ = _0692_ & ~_0929_;
	assign _0931_ = _0930_ | _0928_;
	assign _0932_ = _0931_ & ~_0661_;
	assign _0933_ = _0932_ ^ _0662_;
	assign _0934_ = _0871_ ^ _0850_;
	assign _0935_ = ~(_0934_ ^ _0933_);
	assign _0936_ = _0930_ ^ _0928_;
	assign _0937_ = _0818_ & ~_0855_;
	assign _0938_ = _0937_ ^ _0854_;
	assign _0939_ = _0938_ ^ _0936_;
	assign _0940_ = _0935_ & ~_0939_;
	assign _0941_ = _0749_ | _0695_;
	assign _0942_ = _0941_ & ~_0689_;
	assign _0943_ = _0942_ ^ _0690_;
	assign _0944_ = _0855_ ^ _0818_;
	assign _0945_ = ~(_0944_ ^ _0943_);
	assign _0946_ = _0749_ ^ _0695_;
	assign _0947_ = _0879_ & ~_0804_;
	assign _0948_ = _0947_ ^ _0803_;
	assign _0949_ = ~(_0948_ ^ _0946_);
	assign _0950_ = ~(_0949_ & _0945_);
	assign _0951_ = _0950_ | ~_0940_;
	assign _0952_ = _0951_ | ~_0927_;
	assign _0953_ = _0943_ | ~_0944_;
	assign _0954_ = _0946_ | ~_0948_;
	assign _0955_ = _0945_ & ~_0954_;
	assign _0956_ = _0953_ & ~_0955_;
	assign _0957_ = _0940_ & ~_0956_;
	assign _0958_ = _0933_ & ~_0934_;
	assign _0959_ = _0936_ | ~_0938_;
	assign _0960_ = _0935_ & ~_0959_;
	assign _0961_ = _0960_ | _0958_;
	assign _0962_ = _0961_ | _0957_;
	assign _0963_ = _0952_ & ~_0962_;
	assign _0964_ = ~(_0963_ | _0875_);
	assign _0965_ = _0868_ & _0753_;
	assign _0966_ = _0870_ | ~_0873_;
	assign _0967_ = _0869_ & ~_0966_;
	assign _0968_ = _0967_ | _0965_;
	assign _0969_ = _0968_ | _0964_;
	assign _0970_ = ~(\mchip.chip_design.score [7] & \mchip.chip_design.score [6]);
	assign _0971_ = ~(_0970_ | _0751_);
	assign _0972_ = _0867_ | _0860_;
	assign _0973_ = _0972_ ^ _0971_;
	assign _0974_ = ~(_0973_ ^ _0969_);
	assign _0975_ = _0974_ ^ \mchip.chip_design.timing.bounce_cnt [16];
	assign _0976_ = _0972_ | _0971_;
	assign _0977_ = _0973_ & _0969_;
	assign _0978_ = _0976_ & ~_0977_;
	assign _0979_ = ~(_0978_ ^ _0972_);
	assign _0980_ = _0979_ ^ \mchip.chip_design.timing.bounce_cnt [17];
	assign _0981_ = _0975_ & ~_0980_;
	assign _0982_ = _0971_ | ~_0972_;
	assign _0983_ = _0968_ & ~_0982_;
	assign _0984_ = _0972_ & ~_0983_;
	assign _0985_ = _0982_ | _0875_;
	assign _0986_ = _0962_ & ~_0985_;
	assign _0987_ = _0984_ & ~_0986_;
	assign _0988_ = _0985_ | _0951_;
	assign _0989_ = _0927_ & ~_0988_;
	assign _0990_ = _0987_ & ~_0989_;
	assign _0991_ = _0972_ & ~_0990_;
	assign _0992_ = ~(_0991_ ^ \mchip.chip_design.timing.bounce_cnt [19]);
	assign _0993_ = ~(_0990_ ^ _0972_);
	assign _0994_ = _0993_ ^ \mchip.chip_design.timing.bounce_cnt [18];
	assign _0995_ = _0994_ | _0992_;
	assign _0996_ = _0981_ & ~_0995_;
	assign _0997_ = ~(_0991_ ^ \mchip.chip_design.timing.bounce_cnt [23]);
	assign _0998_ = ~(_0991_ ^ \mchip.chip_design.timing.bounce_cnt [22]);
	assign _0999_ = _0998_ | _0997_;
	assign _1000_ = ~(_0991_ ^ \mchip.chip_design.timing.bounce_cnt [21]);
	assign _1001_ = ~(_0991_ ^ \mchip.chip_design.timing.bounce_cnt [20]);
	assign _1002_ = _1001_ | _1000_;
	assign _1003_ = _1002_ | _0999_;
	assign _1004_ = _0996_ & ~_1003_;
	assign _1005_ = ~(_0991_ ^ \mchip.chip_design.timing.bounce_cnt [26]);
	assign _1006_ = ~(_0991_ ^ \mchip.chip_design.timing.bounce_cnt [25]);
	assign _1007_ = ~\mchip.chip_design.timing.bounce_cnt [24];
	assign _1008_ = _0991_ ^ _1007_;
	assign _1009_ = _1008_ | _1006_;
	assign _1010_ = _1009_ | _1005_;
	assign _1011_ = _1004_ & ~_1010_;
	assign _1012_ = _0874_ & ~_0963_;
	assign _1013_ = _0966_ & ~_1012_;
	assign _1014_ = ~(_1013_ ^ _0869_);
	assign _1015_ = _1014_ ^ \mchip.chip_design.timing.bounce_cnt [15];
	assign _1016_ = ~(_0963_ ^ _0874_);
	assign _1017_ = _1016_ ^ \mchip.chip_design.timing.bounce_cnt [14];
	assign _1018_ = _1017_ | _1015_;
	assign _1019_ = _0927_ & ~_0950_;
	assign _1020_ = _0956_ & ~_1019_;
	assign _1021_ = ~(_1020_ | _0939_);
	assign _1022_ = _0959_ & ~_1021_;
	assign _1023_ = ~(_1022_ ^ _0935_);
	assign _1024_ = _1023_ ^ \mchip.chip_design.timing.bounce_cnt [13];
	assign _1025_ = _1020_ ^ _0939_;
	assign _1026_ = _1025_ ^ \mchip.chip_design.timing.bounce_cnt [12];
	assign _1027_ = _1026_ | _1024_;
	assign _1028_ = _1027_ | _1018_;
	assign _1029_ = _0949_ & ~_0926_;
	assign _1030_ = _0954_ & ~_1029_;
	assign _1031_ = ~(_1030_ ^ _0945_);
	assign _1032_ = _1031_ ^ \mchip.chip_design.timing.bounce_cnt [11];
	assign _1033_ = ~(_0949_ ^ _0926_);
	assign _1034_ = _1033_ ^ \mchip.chip_design.timing.bounce_cnt [10];
	assign _1035_ = _1034_ | _1032_;
	assign _1036_ = _0921_ & ~_0923_;
	assign _1037_ = _0902_ & ~_1036_;
	assign _1038_ = _0890_ & ~_1037_;
	assign _1039_ = _0886_ & ~_1038_;
	assign _1040_ = ~(_1039_ ^ _0887_);
	assign _1041_ = _1040_ ^ \mchip.chip_design.timing.bounce_cnt [9];
	assign _1042_ = ~(_1037_ ^ _0890_);
	assign _1043_ = _1042_ ^ \mchip.chip_design.timing.bounce_cnt [8];
	assign _1044_ = _1043_ | _1041_;
	assign _1045_ = _1044_ | _1035_;
	assign _1046_ = _1045_ | _1028_;
	assign _1047_ = \mchip.chip_design.timing.bounce_cnt [1] | ~\mchip.chip_design.timing.bounce_cnt [0];
	assign \mchip.chip_design.timing.score_base [3] = \mchip.chip_design.score [1] ^ \mchip.chip_design.score [0];
	assign _1048_ = ~(\mchip.chip_design.timing.score_base [3] ^ io_in[6]);
	assign _1049_ = _1048_ ^ _1072_[0];
	assign _1050_ = _1049_ ^ \mchip.chip_design.timing.bounce_cnt [3];
	assign _1051_ = \mchip.chip_design.score [0] ^ \mchip.chip_design.timing.bounce_cnt [2];
	assign _1052_ = _1051_ | _1050_;
	assign _1053_ = _1052_ | _1047_;
	assign _1054_ = _0922_ & ~_0920_;
	assign _1055_ = _0899_ & ~_1054_;
	assign _1056_ = ~(_1055_ ^ _0900_);
	assign _1057_ = _1056_ ^ \mchip.chip_design.timing.bounce_cnt [7];
	assign _1058_ = ~(_0922_ ^ _0920_);
	assign _1059_ = _1058_ ^ \mchip.chip_design.timing.bounce_cnt [6];
	assign _1060_ = _1059_ | _1057_;
	assign _1061_ = _0917_ & _0916_;
	assign _1062_ = _0912_ & ~_1061_;
	assign _1063_ = ~(_1062_ ^ _0913_);
	assign _1064_ = _1063_ ^ \mchip.chip_design.timing.bounce_cnt [5];
	assign _1065_ = _0917_ ^ _0916_;
	assign _1066_ = _1065_ ^ \mchip.chip_design.timing.bounce_cnt [4];
	assign _1067_ = _1066_ | _1064_;
	assign _1068_ = _1067_ | _1060_;
	assign _1069_ = _1068_ | _1053_;
	assign _1070_ = _1069_ | _1046_;
	assign _1071_ = _1011_ & ~_1070_;
	assign _0013_ = _1071_ | io_in[13];
	assign _0004_ = _0547_ | \mchip.chip_design.genblk1[0].col.stack_dec ;
	assign _0005_ = _0560_ | \mchip.chip_design.genblk1[0].col.stack_dec ;
	assign _0006_ = _0574_ | \mchip.chip_design.genblk1[0].col.stack_dec ;
	assign _0007_ = _0587_ | \mchip.chip_design.genblk1[0].col.stack_dec ;
	assign _0008_ = _0519_ | \mchip.chip_design.genblk1[0].col.stack_dec ;
	assign _0009_ = _0532_ | \mchip.chip_design.genblk1[0].col.stack_dec ;
	assign _0010_ = _0492_ | \mchip.chip_design.genblk1[0].col.stack_dec ;
	assign _0011_ = _0505_ | \mchip.chip_design.genblk1[0].col.stack_dec ;
	assign _0066_ = ~(\mchip.chip_design.bounce.bounce_pos [0] | \mchip.chip_design.bounce.bounce_pos [1]);
	assign _0067_ = _0066_ & ~\mchip.chip_design.bounce.bounce_pos [2];
	assign _0068_ = _0067_ & ~\mchip.chip_design.bounce.state ;
	assign _0014_ = _0068_ | io_in[13];
	assign _0069_ = ~\mchip.chip_design.state [1];
	assign _0070_ = ~(\mchip.chip_design.state [3] | \mchip.chip_design.state [2]);
	assign _0071_ = (_0070_ ? _0069_ : \mchip.chip_design.new_game );
	assign _0015_ = _0071_ | io_in[13];
	assign _0072_ = \mchip.chip_design.timing.bounce_cnt [1] | \mchip.chip_design.timing.bounce_cnt [0];
	assign _0073_ = _0072_ | _1052_;
	assign _0074_ = _0073_ | _1068_;
	assign _0075_ = _0074_ | _1046_;
	assign _0076_ = _1011_ & ~_0075_;
	assign _0077_ = \mchip.chip_design.new_game  & ~_0626_;
	assign _0078_ = _0069_ & ~_0077_;
	assign _0079_ = _0626_ & ~\mchip.chip_design.state [1];
	assign _0080_ = (_0079_ ? _0475_ : _0078_);
	assign _0081_ = _0076_ & ~_0080_;
	assign _0082_ = ~(_0475_ | _0474_);
	assign _0083_ = (_0079_ ? _0082_ : \mchip.chip_design.state [1]);
	assign _0017_ = _0081_ & ~_0083_;
	assign \mchip.chip_design.bounce.game_running  = ~_0080_;
	assign _0084_ = ~\mchip.chip_design.bounce.bounce_pos [2];
	assign _0085_ = ~(\mchip.chip_design.bounce.bounce_pos [0] & \mchip.chip_design.bounce.bounce_pos [1]);
	assign _0086_ = _0085_ | _0084_;
	assign _0016_ = \mchip.chip_design.bounce.state  & ~_0086_;
	assign _0087_ = \mchip.chip_design.timing.drop_cnt [1] | \mchip.chip_design.timing.drop_cnt [0];
	assign _0088_ = _0087_ | _0613_;
	assign _0089_ = _0088_ | _0617_;
	assign _0090_ = _0089_ | _0611_;
	assign _0091_ = _0604_ & ~_0090_;
	assign _0092_ = ~(_0504_ & \mchip.chip_design.genblk1[0].col.state );
	assign _0018_ = _0091_ & ~_0092_;
	assign _0019_ = _0092_ | io_in[13];
	assign _0093_ = ~(_0491_ & \mchip.chip_design.genblk1[1].col.state );
	assign _0024_ = _0091_ & ~_0093_;
	assign _0025_ = _0093_ | io_in[13];
	assign _0094_ = ~(_0531_ & \mchip.chip_design.genblk1[2].col.state );
	assign _0030_ = _0091_ & ~_0094_;
	assign _0031_ = _0094_ | io_in[13];
	assign _0095_ = ~(_0518_ & \mchip.chip_design.genblk1[3].col.state );
	assign _0036_ = _0091_ & ~_0095_;
	assign _0037_ = _0095_ | io_in[13];
	assign _0096_ = ~(_0586_ & \mchip.chip_design.genblk1[4].col.state );
	assign _0042_ = _0091_ & ~_0096_;
	assign _0043_ = _0096_ | io_in[13];
	assign _0097_ = ~(_0573_ & \mchip.chip_design.genblk1[5].col.state );
	assign _0048_ = _0091_ & ~_0097_;
	assign _0049_ = _0097_ | io_in[13];
	assign _0098_ = ~(_0559_ & \mchip.chip_design.genblk1[6].col.state );
	assign _0054_ = _0091_ & ~_0098_;
	assign _0055_ = _0098_ | io_in[13];
	assign _0099_ = ~(_0546_ & \mchip.chip_design.genblk1[7].col.state );
	assign _0060_ = _0091_ & ~_0099_;
	assign _0061_ = _0099_ | io_in[13];
	assign _0100_ = io_in[3] | ~io_in[2];
	assign _0101_ = _0100_ | io_in[4];
	assign _0102_ = \mchip.chip_design.genblk1[1].col.stack_pos [0] & ~_0101_;
	assign _0103_ = io_in[2] | ~io_in[3];
	assign _0104_ = _0103_ | io_in[4];
	assign _0105_ = \mchip.chip_design.genblk1[2].col.stack_pos [0] & ~_0104_;
	assign _0106_ = ~(io_in[2] & io_in[3]);
	assign _0107_ = _0106_ | io_in[4];
	assign _0108_ = \mchip.chip_design.genblk1[3].col.stack_pos [0] & ~_0107_;
	assign _0109_ = _0108_ | _0105_;
	assign _0110_ = _0109_ | _0102_;
	assign _0111_ = ~io_in[4];
	assign _0112_ = io_in[2] | io_in[3];
	assign _0113_ = _0112_ | _0111_;
	assign _0114_ = \mchip.chip_design.genblk1[4].col.stack_pos [0] & ~_0113_;
	assign _0115_ = _0100_ | _0111_;
	assign _0116_ = \mchip.chip_design.genblk1[5].col.stack_pos [0] & ~_0115_;
	assign _0117_ = _0116_ | _0114_;
	assign _0118_ = _0103_ | _0111_;
	assign _0119_ = \mchip.chip_design.genblk1[6].col.stack_pos [0] & ~_0118_;
	assign _0120_ = _0106_ | _0111_;
	assign _0121_ = \mchip.chip_design.genblk1[7].col.stack_pos [0] & ~_0120_;
	assign _0122_ = _0121_ | _0119_;
	assign _0123_ = _0122_ | _0117_;
	assign _0124_ = _0123_ | _0110_;
	assign _0125_ = ~(io_in[3] & io_in[4]);
	assign _0126_ = io_in[4] & ~io_in[3];
	assign _0127_ = _0125_ & ~_0126_;
	assign _0128_ = io_in[3] & ~io_in[4];
	assign _0129_ = _0128_ | ~_0101_;
	assign _0130_ = _0127_ & ~_0129_;
	assign _0131_ = (_0130_ ? \mchip.chip_design.genblk1[0].col.stack_pos [0] : _0124_);
	assign io_out[4] = (io_in[5] ? \mchip.chip_design.score [0] : _0131_);
	assign _0132_ = \mchip.chip_design.genblk1[1].col.stack_pos [1] & ~_0101_;
	assign _0133_ = \mchip.chip_design.genblk1[2].col.stack_pos [1] & ~_0104_;
	assign _0134_ = \mchip.chip_design.genblk1[3].col.stack_pos [1] & ~_0107_;
	assign _0135_ = _0134_ | _0133_;
	assign _0136_ = _0135_ | _0132_;
	assign _0137_ = \mchip.chip_design.genblk1[4].col.stack_pos [1] & ~_0113_;
	assign _0138_ = \mchip.chip_design.genblk1[5].col.stack_pos [1] & ~_0115_;
	assign _0139_ = _0138_ | _0137_;
	assign _0140_ = \mchip.chip_design.genblk1[6].col.stack_pos [1] & ~_0118_;
	assign _0141_ = \mchip.chip_design.genblk1[7].col.stack_pos [1] & ~_0120_;
	assign _0142_ = _0141_ | _0140_;
	assign _0143_ = _0142_ | _0139_;
	assign _0144_ = _0143_ | _0136_;
	assign _0145_ = (_0130_ ? \mchip.chip_design.genblk1[0].col.stack_pos [1] : _0144_);
	assign io_out[5] = (io_in[5] ? \mchip.chip_design.score [1] : _0145_);
	assign _0146_ = \mchip.chip_design.genblk1[1].col.stack_pos [2] & ~_0101_;
	assign _0147_ = \mchip.chip_design.genblk1[2].col.stack_pos [2] & ~_0104_;
	assign _0148_ = \mchip.chip_design.genblk1[3].col.stack_pos [2] & ~_0107_;
	assign _0149_ = _0148_ | _0147_;
	assign _0150_ = _0149_ | _0146_;
	assign _0151_ = \mchip.chip_design.genblk1[4].col.stack_pos [2] & ~_0113_;
	assign _0152_ = \mchip.chip_design.genblk1[5].col.stack_pos [2] & ~_0115_;
	assign _0153_ = _0152_ | _0151_;
	assign _0154_ = \mchip.chip_design.genblk1[6].col.stack_pos [2] & ~_0118_;
	assign _0155_ = \mchip.chip_design.genblk1[7].col.stack_pos [2] & ~_0120_;
	assign _0156_ = _0155_ | _0154_;
	assign _0157_ = _0156_ | _0153_;
	assign _0158_ = _0157_ | _0150_;
	assign _0159_ = (_0130_ ? \mchip.chip_design.genblk1[0].col.stack_pos [2] : _0158_);
	assign io_out[6] = (io_in[5] ? \mchip.chip_design.score [2] : _0159_);
	assign _0160_ = \mchip.chip_design.genblk1[1].col.stack_pos [3] & ~_0101_;
	assign _0161_ = \mchip.chip_design.genblk1[2].col.stack_pos [3] & ~_0104_;
	assign _0162_ = \mchip.chip_design.genblk1[3].col.stack_pos [3] & ~_0107_;
	assign _0163_ = _0162_ | _0161_;
	assign _0164_ = _0163_ | _0160_;
	assign _0165_ = \mchip.chip_design.genblk1[4].col.stack_pos [3] & ~_0113_;
	assign _0166_ = \mchip.chip_design.genblk1[5].col.stack_pos [3] & ~_0115_;
	assign _0167_ = _0166_ | _0165_;
	assign _0168_ = \mchip.chip_design.genblk1[6].col.stack_pos [3] & ~_0118_;
	assign _0169_ = \mchip.chip_design.genblk1[7].col.stack_pos [3] & ~_0120_;
	assign _0170_ = _0169_ | _0168_;
	assign _0171_ = _0170_ | _0167_;
	assign _0172_ = _0171_ | _0164_;
	assign _0173_ = (_0130_ ? \mchip.chip_design.genblk1[0].col.stack_pos [3] : _0172_);
	assign io_out[7] = (io_in[5] ? \mchip.chip_design.score [3] : _0173_);
	assign _0174_ = \mchip.chip_design.genblk1[1].col.drop_pos [0] & ~_0101_;
	assign _0175_ = \mchip.chip_design.genblk1[2].col.drop_pos [0] & ~_0104_;
	assign _0176_ = \mchip.chip_design.genblk1[3].col.drop_pos [0] & ~_0107_;
	assign _0177_ = _0176_ | _0175_;
	assign _0178_ = _0177_ | _0174_;
	assign _0179_ = \mchip.chip_design.genblk1[4].col.drop_pos [0] & ~_0113_;
	assign _0180_ = \mchip.chip_design.genblk1[5].col.drop_pos [0] & ~_0115_;
	assign _0181_ = _0180_ | _0179_;
	assign _0182_ = \mchip.chip_design.genblk1[6].col.drop_pos [0] & ~_0118_;
	assign _0183_ = \mchip.chip_design.genblk1[7].col.drop_pos [0] & ~_0120_;
	assign _0184_ = _0183_ | _0182_;
	assign _0185_ = _0184_ | _0181_;
	assign _0186_ = _0185_ | _0178_;
	assign _0187_ = (_0130_ ? \mchip.chip_design.genblk1[0].col.drop_pos [0] : _0186_);
	assign io_out[8] = (io_in[5] ? \mchip.chip_design.score [4] : _0187_);
	assign _0188_ = \mchip.chip_design.genblk1[1].col.drop_pos [1] & ~_0101_;
	assign _0189_ = \mchip.chip_design.genblk1[2].col.drop_pos [1] & ~_0104_;
	assign _0190_ = \mchip.chip_design.genblk1[3].col.drop_pos [1] & ~_0107_;
	assign _0191_ = _0190_ | _0189_;
	assign _0192_ = _0191_ | _0188_;
	assign _0193_ = \mchip.chip_design.genblk1[4].col.drop_pos [1] & ~_0113_;
	assign _0194_ = \mchip.chip_design.genblk1[5].col.drop_pos [1] & ~_0115_;
	assign _0195_ = _0194_ | _0193_;
	assign _0196_ = \mchip.chip_design.genblk1[6].col.drop_pos [1] & ~_0118_;
	assign _0197_ = \mchip.chip_design.genblk1[7].col.drop_pos [1] & ~_0120_;
	assign _0198_ = _0197_ | _0196_;
	assign _0199_ = _0198_ | _0195_;
	assign _0200_ = _0199_ | _0192_;
	assign _0201_ = (_0130_ ? \mchip.chip_design.genblk1[0].col.drop_pos [1] : _0200_);
	assign io_out[9] = (io_in[5] ? \mchip.chip_design.score [5] : _0201_);
	assign _0202_ = \mchip.chip_design.genblk1[1].col.drop_pos [2] & ~_0101_;
	assign _0203_ = \mchip.chip_design.genblk1[2].col.drop_pos [2] & ~_0104_;
	assign _0204_ = \mchip.chip_design.genblk1[3].col.drop_pos [2] & ~_0107_;
	assign _0205_ = _0204_ | _0203_;
	assign _0206_ = _0205_ | _0202_;
	assign _0207_ = \mchip.chip_design.genblk1[4].col.drop_pos [2] & ~_0113_;
	assign _0208_ = \mchip.chip_design.genblk1[5].col.drop_pos [2] & ~_0115_;
	assign _0209_ = _0208_ | _0207_;
	assign _0210_ = \mchip.chip_design.genblk1[6].col.drop_pos [2] & ~_0118_;
	assign _0211_ = \mchip.chip_design.genblk1[7].col.drop_pos [2] & ~_0120_;
	assign _0212_ = _0211_ | _0210_;
	assign _0213_ = _0212_ | _0209_;
	assign _0214_ = _0213_ | _0206_;
	assign _0215_ = (_0130_ ? \mchip.chip_design.genblk1[0].col.drop_pos [2] : _0214_);
	assign io_out[10] = (io_in[5] ? \mchip.chip_design.score [6] : _0215_);
	assign _0216_ = \mchip.chip_design.genblk1[1].col.drop_pos [3] & ~_0101_;
	assign _0217_ = \mchip.chip_design.genblk1[2].col.drop_pos [3] & ~_0104_;
	assign _0218_ = \mchip.chip_design.genblk1[3].col.drop_pos [3] & ~_0107_;
	assign _0219_ = _0218_ | _0217_;
	assign _0220_ = _0219_ | _0216_;
	assign _0221_ = \mchip.chip_design.genblk1[4].col.drop_pos [3] & ~_0113_;
	assign _0222_ = \mchip.chip_design.genblk1[5].col.drop_pos [3] & ~_0115_;
	assign _0223_ = _0222_ | _0221_;
	assign _0224_ = \mchip.chip_design.genblk1[6].col.drop_pos [3] & ~_0118_;
	assign _0225_ = \mchip.chip_design.genblk1[7].col.drop_pos [3] & ~_0120_;
	assign _0226_ = _0225_ | _0224_;
	assign _0227_ = _0226_ | _0223_;
	assign _0228_ = _0227_ | _0220_;
	assign _0229_ = (_0130_ ? \mchip.chip_design.genblk1[0].col.drop_pos [3] : _0228_);
	assign io_out[11] = (io_in[5] ? \mchip.chip_design.score [7] : _0229_);
	assign _1074_[0] = ~\mchip.chip_design.bounce.bounce_pos [0];
	assign _0230_ = ~(\mchip.chip_design.state [0] | \mchip.chip_design.state [1]);
	assign _0231_ = _0230_ & ~\mchip.chip_design.state [3];
	assign _0232_ = _0066_ ^ _0084_;
	assign _0233_ = ~_0232_;
	assign _0234_ = \mchip.chip_design.bounce.bounce_pos [0] | ~\mchip.chip_design.bounce.bounce_pos [1];
	assign _0235_ = \mchip.chip_design.bounce.bounce_pos [1] | ~\mchip.chip_design.bounce.bounce_pos [0];
	assign _0236_ = ~(_0235_ & _0234_);
	assign _0237_ = ~(_0067_ & _1074_[0]);
	assign _0238_ = _0237_ | _0236_;
	assign _0239_ = _0233_ & ~_0238_;
	assign _0240_ = ~(_0239_ & _0067_);
	assign _0241_ = _0240_ | _0474_;
	assign _0242_ = _0241_ | _0475_;
	assign _0243_ = _0231_ & ~_0242_;
	assign \mchip.chip_design.genblk1[0].col.nextState  = (\mchip.chip_design.genblk1[0].col.state  ? _0504_ : _0243_);
	assign _0244_ = \mchip.chip_design.genblk1[0].col.stack_dec  & ~\mchip.chip_design.genblk1[0].col.stack_pos [0];
	assign _0245_ = ~(\mchip.chip_design.genblk1[0].col.stack_dec  | \mchip.chip_design.genblk1[0].col.stack_pos [0]);
	assign _0020_ = _0245_ | _0244_;
	assign _0021_ = _0500_ ^ \mchip.chip_design.genblk1[0].col.stack_dec ;
	assign _0246_ = _0438_ ^ \mchip.chip_design.genblk1[0].col.stack_pos [2];
	assign _0022_ = (\mchip.chip_design.genblk1[0].col.stack_dec  ? _0246_ : _0497_);
	assign _0247_ = _0438_ & ~\mchip.chip_design.genblk1[0].col.stack_pos [2];
	assign _0248_ = _0247_ ^ \mchip.chip_design.genblk1[0].col.stack_pos [3];
	assign _0023_ = (\mchip.chip_design.genblk1[0].col.stack_dec  ? _0248_ : _0495_);
	assign _0249_ = _0235_ | ~_0232_;
	assign _0250_ = _0249_ | _0067_;
	assign _0251_ = _0250_ | _0474_;
	assign _0252_ = _0251_ | _0475_;
	assign _0253_ = _0231_ & ~_0252_;
	assign \mchip.chip_design.genblk1[1].col.nextState  = (\mchip.chip_design.genblk1[1].col.state  ? _0491_ : _0253_);
	assign _0254_ = \mchip.chip_design.genblk1[0].col.stack_dec  & ~\mchip.chip_design.genblk1[1].col.stack_pos [0];
	assign _0255_ = ~(\mchip.chip_design.genblk1[0].col.stack_dec  | \mchip.chip_design.genblk1[1].col.stack_pos [0]);
	assign _0026_ = _0255_ | _0254_;
	assign _0027_ = _0482_ ^ \mchip.chip_design.genblk1[0].col.stack_dec ;
	assign _0256_ = _0435_ ^ \mchip.chip_design.genblk1[1].col.stack_pos [2];
	assign _0028_ = (\mchip.chip_design.genblk1[0].col.stack_dec  ? _0256_ : _0488_);
	assign _0257_ = _0435_ & ~\mchip.chip_design.genblk1[1].col.stack_pos [2];
	assign _0258_ = _0257_ ^ \mchip.chip_design.genblk1[1].col.stack_pos [3];
	assign _0029_ = (\mchip.chip_design.genblk1[0].col.stack_dec  ? _0258_ : _0486_);
	assign _0259_ = _0234_ | ~_0232_;
	assign _0260_ = _0259_ | _0067_;
	assign _0261_ = _0260_ | _0474_;
	assign _0262_ = _0261_ | _0475_;
	assign _0263_ = _0231_ & ~_0262_;
	assign \mchip.chip_design.genblk1[2].col.nextState  = (\mchip.chip_design.genblk1[2].col.state  ? _0531_ : _0263_);
	assign _0264_ = \mchip.chip_design.genblk1[0].col.stack_dec  & ~\mchip.chip_design.genblk1[2].col.stack_pos [0];
	assign _0265_ = ~(\mchip.chip_design.genblk1[0].col.stack_dec  | \mchip.chip_design.genblk1[2].col.stack_pos [0]);
	assign _0032_ = _0265_ | _0264_;
	assign _0033_ = _0522_ ^ \mchip.chip_design.genblk1[0].col.stack_dec ;
	assign _0266_ = _0445_ ^ \mchip.chip_design.genblk1[2].col.stack_pos [2];
	assign _0034_ = (\mchip.chip_design.genblk1[0].col.stack_dec  ? _0266_ : _0528_);
	assign _0267_ = _0445_ & ~\mchip.chip_design.genblk1[2].col.stack_pos [2];
	assign _0268_ = _0267_ ^ \mchip.chip_design.genblk1[2].col.stack_pos [3];
	assign _0035_ = (\mchip.chip_design.genblk1[0].col.stack_dec  ? _0268_ : _0526_);
	assign _0269_ = _0085_ | ~_0232_;
	assign _0270_ = _0269_ | _0067_;
	assign _0271_ = _0270_ | _0474_;
	assign _0272_ = _0271_ | _0475_;
	assign _0273_ = _0231_ & ~_0272_;
	assign \mchip.chip_design.genblk1[3].col.nextState  = (\mchip.chip_design.genblk1[3].col.state  ? _0518_ : _0273_);
	assign _0274_ = \mchip.chip_design.genblk1[0].col.stack_dec  & ~\mchip.chip_design.genblk1[3].col.stack_pos [0];
	assign _0275_ = ~(\mchip.chip_design.genblk1[0].col.stack_dec  | \mchip.chip_design.genblk1[3].col.stack_pos [0]);
	assign _0038_ = _0275_ | _0274_;
	assign _0039_ = _0509_ ^ \mchip.chip_design.genblk1[0].col.stack_dec ;
	assign _0276_ = _0442_ ^ \mchip.chip_design.genblk1[3].col.stack_pos [2];
	assign _0040_ = (\mchip.chip_design.genblk1[0].col.stack_dec  ? _0276_ : _0515_);
	assign _0277_ = _0442_ & ~\mchip.chip_design.genblk1[3].col.stack_pos [2];
	assign _0278_ = _0277_ ^ \mchip.chip_design.genblk1[3].col.stack_pos [3];
	assign _0041_ = (\mchip.chip_design.genblk1[0].col.stack_dec  ? _0278_ : _0513_);
	assign _0279_ = _0067_ | \mchip.chip_design.bounce.bounce_pos [0];
	assign _0280_ = _0279_ | _0236_;
	assign _0281_ = _0280_ | _0233_;
	assign _0282_ = _0281_ | _0067_;
	assign _0283_ = _0282_ | _0474_;
	assign _0284_ = _0283_ | _0475_;
	assign _0285_ = _0231_ & ~_0284_;
	assign \mchip.chip_design.genblk1[4].col.nextState  = (\mchip.chip_design.genblk1[4].col.state  ? _0586_ : _0285_);
	assign _0286_ = \mchip.chip_design.genblk1[0].col.stack_dec  & ~\mchip.chip_design.genblk1[4].col.stack_pos [0];
	assign _0287_ = ~(\mchip.chip_design.genblk1[0].col.stack_dec  | \mchip.chip_design.genblk1[4].col.stack_pos [0]);
	assign _0044_ = _0287_ | _0286_;
	assign _0045_ = _0577_ ^ \mchip.chip_design.genblk1[0].col.stack_dec ;
	assign _0288_ = _0460_ ^ \mchip.chip_design.genblk1[4].col.stack_pos [2];
	assign _0046_ = (\mchip.chip_design.genblk1[0].col.stack_dec  ? _0288_ : _0583_);
	assign _0289_ = _0460_ & ~\mchip.chip_design.genblk1[4].col.stack_pos [2];
	assign _0290_ = _0289_ ^ \mchip.chip_design.genblk1[4].col.stack_pos [3];
	assign _0047_ = (\mchip.chip_design.genblk1[0].col.stack_dec  ? _0290_ : _0581_);
	assign _0291_ = _0235_ | _0232_;
	assign _0292_ = _0291_ | _0067_;
	assign _0293_ = _0292_ | _0474_;
	assign _0294_ = _0293_ | _0475_;
	assign _0295_ = _0231_ & ~_0294_;
	assign \mchip.chip_design.genblk1[5].col.nextState  = (\mchip.chip_design.genblk1[5].col.state  ? _0573_ : _0295_);
	assign _0296_ = \mchip.chip_design.genblk1[0].col.stack_dec  & ~\mchip.chip_design.genblk1[5].col.stack_pos [0];
	assign _0297_ = ~(\mchip.chip_design.genblk1[0].col.stack_dec  | \mchip.chip_design.genblk1[5].col.stack_pos [0]);
	assign _0050_ = _0297_ | _0296_;
	assign _0051_ = _0564_ ^ \mchip.chip_design.genblk1[0].col.stack_dec ;
	assign _0298_ = _0457_ ^ \mchip.chip_design.genblk1[5].col.stack_pos [2];
	assign _0052_ = (\mchip.chip_design.genblk1[0].col.stack_dec  ? _0298_ : _0570_);
	assign _0299_ = _0457_ & ~\mchip.chip_design.genblk1[5].col.stack_pos [2];
	assign _0300_ = _0299_ ^ \mchip.chip_design.genblk1[5].col.stack_pos [3];
	assign _0053_ = (\mchip.chip_design.genblk1[0].col.stack_dec  ? _0300_ : _0568_);
	assign _0301_ = _0234_ | _0232_;
	assign _0302_ = _0301_ | _0067_;
	assign _0303_ = _0302_ | _0474_;
	assign _0304_ = _0303_ | _0475_;
	assign _0305_ = _0231_ & ~_0304_;
	assign \mchip.chip_design.genblk1[6].col.nextState  = (\mchip.chip_design.genblk1[6].col.state  ? _0559_ : _0305_);
	assign _0306_ = \mchip.chip_design.genblk1[0].col.stack_dec  & ~\mchip.chip_design.genblk1[6].col.stack_pos [0];
	assign _0307_ = ~(\mchip.chip_design.genblk1[0].col.stack_dec  | \mchip.chip_design.genblk1[6].col.stack_pos [0]);
	assign _0056_ = _0307_ | _0306_;
	assign _0057_ = _0550_ ^ \mchip.chip_design.genblk1[0].col.stack_dec ;
	assign _0308_ = _0453_ ^ \mchip.chip_design.genblk1[6].col.stack_pos [2];
	assign _0058_ = (\mchip.chip_design.genblk1[0].col.stack_dec  ? _0308_ : _0556_);
	assign _0309_ = _0453_ & ~\mchip.chip_design.genblk1[6].col.stack_pos [2];
	assign _0310_ = _0309_ ^ \mchip.chip_design.genblk1[6].col.stack_pos [3];
	assign _0059_ = (\mchip.chip_design.genblk1[0].col.stack_dec  ? _0310_ : _0554_);
	assign _0311_ = _0232_ | _0085_;
	assign _0312_ = _0311_ | _0067_;
	assign _0313_ = _0312_ | _0474_;
	assign _0314_ = _0313_ | _0475_;
	assign _0315_ = _0231_ & ~_0314_;
	assign \mchip.chip_design.genblk1[7].col.nextState  = (\mchip.chip_design.genblk1[7].col.state  ? _0546_ : _0315_);
	assign _0316_ = \mchip.chip_design.genblk1[0].col.stack_dec  & ~\mchip.chip_design.genblk1[7].col.stack_pos [0];
	assign _0317_ = ~(\mchip.chip_design.genblk1[0].col.stack_dec  | \mchip.chip_design.genblk1[7].col.stack_pos [0]);
	assign _0062_ = _0317_ | _0316_;
	assign _0063_ = _0537_ ^ \mchip.chip_design.genblk1[0].col.stack_dec ;
	assign _0318_ = _0450_ ^ \mchip.chip_design.genblk1[7].col.stack_pos [2];
	assign _0064_ = (\mchip.chip_design.genblk1[0].col.stack_dec  ? _0318_ : _0543_);
	assign _0319_ = _0450_ & ~\mchip.chip_design.genblk1[7].col.stack_pos [2];
	assign _0320_ = _0319_ ^ \mchip.chip_design.genblk1[7].col.stack_pos [3];
	assign _0065_ = (\mchip.chip_design.genblk1[0].col.stack_dec  ? _0320_ : _0541_);
	assign _1087_[1] = \mchip.chip_design.timing.bounce_cnt [1] ^ \mchip.chip_design.timing.bounce_cnt [0];
	assign _0321_ = \mchip.chip_design.timing.bounce_cnt [1] & \mchip.chip_design.timing.bounce_cnt [0];
	assign _1087_[2] = _0321_ ^ \mchip.chip_design.timing.bounce_cnt [2];
	assign _0322_ = _0321_ & \mchip.chip_design.timing.bounce_cnt [2];
	assign _1087_[3] = _0322_ ^ \mchip.chip_design.timing.bounce_cnt [3];
	assign _0323_ = ~(\mchip.chip_design.timing.bounce_cnt [3] & \mchip.chip_design.timing.bounce_cnt [2]);
	assign _0324_ = _0321_ & ~_0323_;
	assign _1087_[4] = _0324_ ^ \mchip.chip_design.timing.bounce_cnt [4];
	assign _0325_ = _0324_ & \mchip.chip_design.timing.bounce_cnt [4];
	assign _1087_[5] = _0325_ ^ \mchip.chip_design.timing.bounce_cnt [5];
	assign _0326_ = ~(\mchip.chip_design.timing.bounce_cnt [5] & \mchip.chip_design.timing.bounce_cnt [4]);
	assign _0327_ = _0324_ & ~_0326_;
	assign _1087_[6] = _0327_ ^ \mchip.chip_design.timing.bounce_cnt [6];
	assign _0328_ = _0327_ & \mchip.chip_design.timing.bounce_cnt [6];
	assign _1087_[7] = _0328_ ^ \mchip.chip_design.timing.bounce_cnt [7];
	assign _0329_ = ~(\mchip.chip_design.timing.bounce_cnt [7] & \mchip.chip_design.timing.bounce_cnt [6]);
	assign _0330_ = _0329_ | _0326_;
	assign _0331_ = _0324_ & ~_0330_;
	assign _1087_[8] = _0331_ ^ \mchip.chip_design.timing.bounce_cnt [8];
	assign _0332_ = _0331_ & \mchip.chip_design.timing.bounce_cnt [8];
	assign _1087_[9] = _0332_ ^ \mchip.chip_design.timing.bounce_cnt [9];
	assign _0333_ = ~(\mchip.chip_design.timing.bounce_cnt [9] & \mchip.chip_design.timing.bounce_cnt [8]);
	assign _0334_ = _0331_ & ~_0333_;
	assign _1087_[10] = _0334_ ^ \mchip.chip_design.timing.bounce_cnt [10];
	assign _0335_ = _0334_ & \mchip.chip_design.timing.bounce_cnt [10];
	assign _1087_[11] = _0335_ ^ \mchip.chip_design.timing.bounce_cnt [11];
	assign _0336_ = ~(\mchip.chip_design.timing.bounce_cnt [11] & \mchip.chip_design.timing.bounce_cnt [10]);
	assign _0337_ = _0336_ | _0333_;
	assign _0338_ = _0331_ & ~_0337_;
	assign _1087_[12] = _0338_ ^ \mchip.chip_design.timing.bounce_cnt [12];
	assign _0339_ = _0338_ & \mchip.chip_design.timing.bounce_cnt [12];
	assign _1087_[13] = _0339_ ^ \mchip.chip_design.timing.bounce_cnt [13];
	assign _0340_ = ~(\mchip.chip_design.timing.bounce_cnt [13] & \mchip.chip_design.timing.bounce_cnt [12]);
	assign _0341_ = _0338_ & ~_0340_;
	assign _1087_[14] = _0341_ ^ \mchip.chip_design.timing.bounce_cnt [14];
	assign _0342_ = _0341_ & \mchip.chip_design.timing.bounce_cnt [14];
	assign _1087_[15] = _0342_ ^ \mchip.chip_design.timing.bounce_cnt [15];
	assign _0343_ = ~(\mchip.chip_design.timing.bounce_cnt [15] & \mchip.chip_design.timing.bounce_cnt [14]);
	assign _0344_ = _0343_ | _0340_;
	assign _0345_ = _0344_ | _0337_;
	assign _0346_ = _0331_ & ~_0345_;
	assign _1087_[16] = _0346_ ^ \mchip.chip_design.timing.bounce_cnt [16];
	assign _0347_ = _0346_ & \mchip.chip_design.timing.bounce_cnt [16];
	assign _1087_[17] = _0347_ ^ \mchip.chip_design.timing.bounce_cnt [17];
	assign _0348_ = ~(\mchip.chip_design.timing.bounce_cnt [17] & \mchip.chip_design.timing.bounce_cnt [16]);
	assign _0349_ = _0346_ & ~_0348_;
	assign _1087_[18] = _0349_ ^ \mchip.chip_design.timing.bounce_cnt [18];
	assign _0350_ = _0349_ & \mchip.chip_design.timing.bounce_cnt [18];
	assign _1087_[19] = _0350_ ^ \mchip.chip_design.timing.bounce_cnt [19];
	assign _0351_ = ~(\mchip.chip_design.timing.bounce_cnt [19] & \mchip.chip_design.timing.bounce_cnt [18]);
	assign _0352_ = _0351_ | _0348_;
	assign _0353_ = _0346_ & ~_0352_;
	assign _1087_[20] = _0353_ ^ \mchip.chip_design.timing.bounce_cnt [20];
	assign _0354_ = _0353_ & \mchip.chip_design.timing.bounce_cnt [20];
	assign _1087_[21] = _0354_ ^ \mchip.chip_design.timing.bounce_cnt [21];
	assign _0355_ = ~(\mchip.chip_design.timing.bounce_cnt [21] & \mchip.chip_design.timing.bounce_cnt [20]);
	assign _0356_ = _0353_ & ~_0355_;
	assign _1087_[22] = _0356_ ^ \mchip.chip_design.timing.bounce_cnt [22];
	assign _0357_ = _0356_ & \mchip.chip_design.timing.bounce_cnt [22];
	assign _1087_[23] = _0357_ ^ \mchip.chip_design.timing.bounce_cnt [23];
	assign _0358_ = ~(\mchip.chip_design.timing.bounce_cnt [23] & \mchip.chip_design.timing.bounce_cnt [22]);
	assign _0359_ = _0358_ | _0355_;
	assign _0360_ = _0359_ | _0352_;
	assign _0361_ = _0346_ & ~_0360_;
	assign _1087_[24] = _0361_ ^ \mchip.chip_design.timing.bounce_cnt [24];
	assign _0362_ = _0361_ & ~_1007_;
	assign _1087_[25] = _0362_ ^ \mchip.chip_design.timing.bounce_cnt [25];
	assign _0363_ = ~(\mchip.chip_design.timing.bounce_cnt [25] & \mchip.chip_design.timing.bounce_cnt [24]);
	assign _0364_ = _0361_ & ~_0363_;
	assign _1087_[26] = _0364_ ^ \mchip.chip_design.timing.bounce_cnt [26];
	assign _1073_[2] = _0737_ ^ \mchip.chip_design.score [2];
	assign _0365_ = _0737_ & ~_0713_;
	assign _1073_[3] = _0365_ ^ \mchip.chip_design.score [3];
	assign _0366_ = _0737_ & ~_0709_;
	assign _1073_[4] = _0366_ ^ \mchip.chip_design.score [4];
	assign _0367_ = _0366_ & ~_0684_;
	assign _1073_[5] = _0367_ ^ \mchip.chip_design.score [5];
	assign _0368_ = _0366_ & ~_0680_;
	assign _1073_[6] = _0368_ ^ \mchip.chip_design.score [6];
	assign _0369_ = _0368_ & ~_0651_;
	assign _1073_[7] = _0369_ ^ \mchip.chip_design.score [7];
	assign _1085_[1] = \mchip.chip_design.timing.drop_cnt [1] ^ \mchip.chip_design.timing.drop_cnt [0];
	assign _0370_ = \mchip.chip_design.timing.drop_cnt [1] & \mchip.chip_design.timing.drop_cnt [0];
	assign _1085_[2] = _0370_ ^ \mchip.chip_design.timing.drop_cnt [2];
	assign _0371_ = _0370_ & \mchip.chip_design.timing.drop_cnt [2];
	assign _1085_[3] = _0371_ ^ \mchip.chip_design.timing.drop_cnt [3];
	assign _0372_ = ~(\mchip.chip_design.timing.drop_cnt [3] & \mchip.chip_design.timing.drop_cnt [2]);
	assign _0373_ = _0370_ & ~_0372_;
	assign _1085_[4] = _0373_ ^ \mchip.chip_design.timing.drop_cnt [4];
	assign _0374_ = _0373_ & \mchip.chip_design.timing.drop_cnt [4];
	assign _1085_[5] = _0374_ ^ \mchip.chip_design.timing.drop_cnt [5];
	assign _0375_ = ~(\mchip.chip_design.timing.drop_cnt [4] & \mchip.chip_design.timing.drop_cnt [5]);
	assign _0376_ = _0373_ & ~_0375_;
	assign _1085_[6] = _0376_ ^ \mchip.chip_design.timing.drop_cnt [6];
	assign _0377_ = _0376_ & \mchip.chip_design.timing.drop_cnt [6];
	assign _1085_[7] = _0377_ ^ \mchip.chip_design.timing.drop_cnt [7];
	assign _0378_ = ~(\mchip.chip_design.timing.drop_cnt [7] & \mchip.chip_design.timing.drop_cnt [6]);
	assign _0379_ = ~(_0378_ | _0375_);
	assign _0380_ = ~(_0379_ & _0373_);
	assign _1085_[8] = ~(_0380_ ^ \mchip.chip_design.timing.drop_cnt [8]);
	assign _0381_ = \mchip.chip_design.timing.drop_cnt [8] & ~_0380_;
	assign _1085_[9] = _0381_ ^ \mchip.chip_design.timing.drop_cnt [9];
	assign _0382_ = ~(_0380_ | _0609_);
	assign _1085_[10] = _0382_ ^ \mchip.chip_design.timing.drop_cnt [10];
	assign _0383_ = _0382_ & \mchip.chip_design.timing.drop_cnt [10];
	assign _1085_[11] = _0383_ ^ \mchip.chip_design.timing.drop_cnt [11];
	assign _0384_ = ~(\mchip.chip_design.timing.drop_cnt [10] & \mchip.chip_design.timing.drop_cnt [11]);
	assign _0385_ = _0384_ | _0609_;
	assign _0386_ = ~(_0385_ | _0380_);
	assign _1085_[12] = _0386_ ^ \mchip.chip_design.timing.drop_cnt [12];
	assign _0387_ = _0386_ & \mchip.chip_design.timing.drop_cnt [12];
	assign _1085_[13] = _0387_ ^ \mchip.chip_design.timing.drop_cnt [13];
	assign _0388_ = ~(\mchip.chip_design.timing.drop_cnt [12] & \mchip.chip_design.timing.drop_cnt [13]);
	assign _0389_ = _0386_ & ~_0388_;
	assign _1085_[14] = _0389_ ^ \mchip.chip_design.timing.drop_cnt [14];
	assign _0390_ = _0389_ & \mchip.chip_design.timing.drop_cnt [14];
	assign _1085_[15] = _0390_ ^ \mchip.chip_design.timing.drop_cnt [15];
	assign _0391_ = ~(\mchip.chip_design.timing.drop_cnt [14] & \mchip.chip_design.timing.drop_cnt [15]);
	assign _0392_ = _0391_ | _0388_;
	assign _0393_ = _0392_ | _0385_;
	assign _0394_ = ~(_0393_ | _0380_);
	assign _1085_[16] = _0394_ ^ \mchip.chip_design.timing.drop_cnt [16];
	assign _0395_ = _0394_ & \mchip.chip_design.timing.drop_cnt [16];
	assign _1085_[17] = _0395_ ^ \mchip.chip_design.timing.drop_cnt [17];
	assign _0396_ = ~(\mchip.chip_design.timing.drop_cnt [16] & \mchip.chip_design.timing.drop_cnt [17]);
	assign _0397_ = _0394_ & ~_0396_;
	assign _1085_[18] = _0397_ ^ \mchip.chip_design.timing.drop_cnt [18];
	assign _0398_ = _0397_ & \mchip.chip_design.timing.drop_cnt [18];
	assign _1085_[19] = _0398_ ^ \mchip.chip_design.timing.drop_cnt [19];
	assign _0399_ = ~(\mchip.chip_design.timing.drop_cnt [18] & \mchip.chip_design.timing.drop_cnt [19]);
	assign _0400_ = _0399_ | _0396_;
	assign _0401_ = _0394_ & ~_0400_;
	assign _1085_[20] = _0401_ ^ \mchip.chip_design.timing.drop_cnt [20];
	assign _0402_ = _0401_ & \mchip.chip_design.timing.drop_cnt [20];
	assign _1085_[21] = _0402_ ^ \mchip.chip_design.timing.drop_cnt [21];
	assign _0403_ = ~(\mchip.chip_design.timing.drop_cnt [20] & \mchip.chip_design.timing.drop_cnt [21]);
	assign _0404_ = _0401_ & ~_0403_;
	assign _1085_[22] = _0404_ ^ \mchip.chip_design.timing.drop_cnt [22];
	assign _0405_ = _0404_ & \mchip.chip_design.timing.drop_cnt [22];
	assign _1085_[23] = _0405_ ^ \mchip.chip_design.timing.drop_cnt [23];
	assign _0406_ = ~(\mchip.chip_design.timing.drop_cnt [22] & \mchip.chip_design.timing.drop_cnt [23]);
	assign _0407_ = _0406_ | _0403_;
	assign _0408_ = _0407_ | _0400_;
	assign _0409_ = _0394_ & ~_0408_;
	assign _1085_[24] = _0409_ ^ \mchip.chip_design.timing.drop_cnt [24];
	assign _0410_ = _0409_ & \mchip.chip_design.timing.drop_cnt [24];
	assign _1085_[25] = _0410_ ^ \mchip.chip_design.timing.drop_cnt [25];
	assign _0411_ = ~(\mchip.chip_design.timing.drop_cnt [24] & \mchip.chip_design.timing.drop_cnt [25]);
	assign _0412_ = _0409_ & ~_0411_;
	assign _1085_[26] = _0412_ ^ \mchip.chip_design.timing.drop_cnt [26];
	assign _1083_[1] = ~(\mchip.chip_design.genblk1[7].col.drop_pos [1] ^ \mchip.chip_design.genblk1[7].col.drop_pos [0]);
	assign _0413_ = ~(\mchip.chip_design.genblk1[7].col.drop_pos [1] | \mchip.chip_design.genblk1[7].col.drop_pos [0]);
	assign _1083_[2] = _0413_ ^ \mchip.chip_design.genblk1[7].col.drop_pos [2];
	assign _0414_ = _0413_ & ~\mchip.chip_design.genblk1[7].col.drop_pos [2];
	assign _1083_[3] = _0414_ ^ \mchip.chip_design.genblk1[7].col.drop_pos [3];
	assign _1082_[1] = ~(\mchip.chip_design.genblk1[6].col.drop_pos [1] ^ \mchip.chip_design.genblk1[6].col.drop_pos [0]);
	assign _0415_ = ~(\mchip.chip_design.genblk1[6].col.drop_pos [1] | \mchip.chip_design.genblk1[6].col.drop_pos [0]);
	assign _1082_[2] = _0415_ ^ \mchip.chip_design.genblk1[6].col.drop_pos [2];
	assign _0416_ = _0415_ & ~\mchip.chip_design.genblk1[6].col.drop_pos [2];
	assign _1082_[3] = _0416_ ^ \mchip.chip_design.genblk1[6].col.drop_pos [3];
	assign _1081_[1] = ~(\mchip.chip_design.genblk1[5].col.drop_pos [1] ^ \mchip.chip_design.genblk1[5].col.drop_pos [0]);
	assign _0417_ = ~(\mchip.chip_design.genblk1[5].col.drop_pos [1] | \mchip.chip_design.genblk1[5].col.drop_pos [0]);
	assign _1081_[2] = _0417_ ^ \mchip.chip_design.genblk1[5].col.drop_pos [2];
	assign _0418_ = _0417_ & ~\mchip.chip_design.genblk1[5].col.drop_pos [2];
	assign _1081_[3] = _0418_ ^ \mchip.chip_design.genblk1[5].col.drop_pos [3];
	assign _1080_[1] = ~(\mchip.chip_design.genblk1[4].col.drop_pos [1] ^ \mchip.chip_design.genblk1[4].col.drop_pos [0]);
	assign _0419_ = ~(\mchip.chip_design.genblk1[4].col.drop_pos [1] | \mchip.chip_design.genblk1[4].col.drop_pos [0]);
	assign _1080_[2] = _0419_ ^ \mchip.chip_design.genblk1[4].col.drop_pos [2];
	assign _0420_ = _0419_ & ~\mchip.chip_design.genblk1[4].col.drop_pos [2];
	assign _1080_[3] = _0420_ ^ \mchip.chip_design.genblk1[4].col.drop_pos [3];
	assign _1079_[1] = ~(\mchip.chip_design.genblk1[3].col.drop_pos [1] ^ \mchip.chip_design.genblk1[3].col.drop_pos [0]);
	assign _0421_ = ~(\mchip.chip_design.genblk1[3].col.drop_pos [1] | \mchip.chip_design.genblk1[3].col.drop_pos [0]);
	assign _1079_[2] = _0421_ ^ \mchip.chip_design.genblk1[3].col.drop_pos [2];
	assign _0422_ = _0421_ & ~\mchip.chip_design.genblk1[3].col.drop_pos [2];
	assign _1079_[3] = _0422_ ^ \mchip.chip_design.genblk1[3].col.drop_pos [3];
	assign _1078_[1] = ~(\mchip.chip_design.genblk1[2].col.drop_pos [1] ^ \mchip.chip_design.genblk1[2].col.drop_pos [0]);
	assign _0423_ = ~(\mchip.chip_design.genblk1[2].col.drop_pos [1] | \mchip.chip_design.genblk1[2].col.drop_pos [0]);
	assign _1078_[2] = _0423_ ^ \mchip.chip_design.genblk1[2].col.drop_pos [2];
	assign _0424_ = _0423_ & ~\mchip.chip_design.genblk1[2].col.drop_pos [2];
	assign _1078_[3] = _0424_ ^ \mchip.chip_design.genblk1[2].col.drop_pos [3];
	assign _1077_[1] = ~(\mchip.chip_design.genblk1[1].col.drop_pos [1] ^ \mchip.chip_design.genblk1[1].col.drop_pos [0]);
	assign _0425_ = ~(\mchip.chip_design.genblk1[1].col.drop_pos [1] | \mchip.chip_design.genblk1[1].col.drop_pos [0]);
	assign _1077_[2] = _0425_ ^ \mchip.chip_design.genblk1[1].col.drop_pos [2];
	assign _0426_ = _0425_ & ~\mchip.chip_design.genblk1[1].col.drop_pos [2];
	assign _1077_[3] = _0426_ ^ \mchip.chip_design.genblk1[1].col.drop_pos [3];
	assign _1076_[1] = ~(\mchip.chip_design.genblk1[0].col.drop_pos [1] ^ \mchip.chip_design.genblk1[0].col.drop_pos [0]);
	assign _0427_ = ~(\mchip.chip_design.genblk1[0].col.drop_pos [1] | \mchip.chip_design.genblk1[0].col.drop_pos [0]);
	assign _1076_[2] = _0427_ ^ \mchip.chip_design.genblk1[0].col.drop_pos [2];
	assign _0428_ = _0427_ & ~\mchip.chip_design.genblk1[0].col.drop_pos [2];
	assign _1076_[3] = _0428_ ^ \mchip.chip_design.genblk1[0].col.drop_pos [3];
	assign _0429_ = (\mchip.chip_design.bounce.state  ? _0086_ : _0067_);
	assign _0430_ = ~(_0429_ ^ \mchip.chip_design.bounce.bounce_pos [1]);
	assign _1075_[1] = _0430_ ^ \mchip.chip_design.bounce.bounce_pos [0];
	assign _0431_ = \mchip.chip_design.bounce.bounce_pos [1] & ~_0429_;
	assign _0432_ = _0430_ & ~_1074_[0];
	assign _0433_ = _0432_ | _0431_;
	assign _0434_ = _0429_ ^ _0084_;
	assign _1075_[2] = _0434_ ^ _0433_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.chip_design.bounce.bounce_pos [0] <= 1'h0;
		else if (_0017_)
			\mchip.chip_design.bounce.bounce_pos [0] <= _1074_[0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.chip_design.bounce.bounce_pos [1] <= 1'h0;
		else if (_0017_)
			\mchip.chip_design.bounce.bounce_pos [1] <= _1075_[1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.chip_design.bounce.bounce_pos [2] <= 1'h0;
		else if (_0017_)
			\mchip.chip_design.bounce.bounce_pos [2] <= _1075_[2];
	always @(posedge io_in[12]) \mchip.chip_design.prev_drop_button  <= \mchip.chip_design.drop_button ;
	always @(posedge io_in[12]) \mchip.chip_design.drop_button  <= \mchip.chip_design.drop_int ;
	always @(posedge io_in[12])
		if (_0012_)
			\mchip.chip_design.timing.drop_cnt [0] <= 1'h0;
		else
			\mchip.chip_design.timing.drop_cnt [0] <= _1084_[0];
	always @(posedge io_in[12])
		if (_0012_)
			\mchip.chip_design.timing.drop_cnt [1] <= 1'h0;
		else
			\mchip.chip_design.timing.drop_cnt [1] <= _1085_[1];
	always @(posedge io_in[12])
		if (_0012_)
			\mchip.chip_design.timing.drop_cnt [2] <= 1'h0;
		else
			\mchip.chip_design.timing.drop_cnt [2] <= _1085_[2];
	always @(posedge io_in[12])
		if (_0012_)
			\mchip.chip_design.timing.drop_cnt [3] <= 1'h0;
		else
			\mchip.chip_design.timing.drop_cnt [3] <= _1085_[3];
	always @(posedge io_in[12])
		if (_0012_)
			\mchip.chip_design.timing.drop_cnt [4] <= 1'h0;
		else
			\mchip.chip_design.timing.drop_cnt [4] <= _1085_[4];
	always @(posedge io_in[12])
		if (_0012_)
			\mchip.chip_design.timing.drop_cnt [5] <= 1'h0;
		else
			\mchip.chip_design.timing.drop_cnt [5] <= _1085_[5];
	always @(posedge io_in[12])
		if (_0012_)
			\mchip.chip_design.timing.drop_cnt [6] <= 1'h0;
		else
			\mchip.chip_design.timing.drop_cnt [6] <= _1085_[6];
	always @(posedge io_in[12])
		if (_0012_)
			\mchip.chip_design.timing.drop_cnt [7] <= 1'h0;
		else
			\mchip.chip_design.timing.drop_cnt [7] <= _1085_[7];
	always @(posedge io_in[12])
		if (_0012_)
			\mchip.chip_design.timing.drop_cnt [8] <= 1'h0;
		else
			\mchip.chip_design.timing.drop_cnt [8] <= _1085_[8];
	always @(posedge io_in[12])
		if (_0012_)
			\mchip.chip_design.timing.drop_cnt [9] <= 1'h0;
		else
			\mchip.chip_design.timing.drop_cnt [9] <= _1085_[9];
	always @(posedge io_in[12])
		if (_0012_)
			\mchip.chip_design.timing.drop_cnt [10] <= 1'h0;
		else
			\mchip.chip_design.timing.drop_cnt [10] <= _1085_[10];
	always @(posedge io_in[12])
		if (_0012_)
			\mchip.chip_design.timing.drop_cnt [11] <= 1'h0;
		else
			\mchip.chip_design.timing.drop_cnt [11] <= _1085_[11];
	always @(posedge io_in[12])
		if (_0012_)
			\mchip.chip_design.timing.drop_cnt [12] <= 1'h0;
		else
			\mchip.chip_design.timing.drop_cnt [12] <= _1085_[12];
	always @(posedge io_in[12])
		if (_0012_)
			\mchip.chip_design.timing.drop_cnt [13] <= 1'h0;
		else
			\mchip.chip_design.timing.drop_cnt [13] <= _1085_[13];
	always @(posedge io_in[12])
		if (_0012_)
			\mchip.chip_design.timing.drop_cnt [14] <= 1'h0;
		else
			\mchip.chip_design.timing.drop_cnt [14] <= _1085_[14];
	always @(posedge io_in[12])
		if (_0012_)
			\mchip.chip_design.timing.drop_cnt [15] <= 1'h0;
		else
			\mchip.chip_design.timing.drop_cnt [15] <= _1085_[15];
	always @(posedge io_in[12])
		if (_0012_)
			\mchip.chip_design.timing.drop_cnt [16] <= 1'h0;
		else
			\mchip.chip_design.timing.drop_cnt [16] <= _1085_[16];
	always @(posedge io_in[12])
		if (_0012_)
			\mchip.chip_design.timing.drop_cnt [17] <= 1'h0;
		else
			\mchip.chip_design.timing.drop_cnt [17] <= _1085_[17];
	always @(posedge io_in[12])
		if (_0012_)
			\mchip.chip_design.timing.drop_cnt [18] <= 1'h0;
		else
			\mchip.chip_design.timing.drop_cnt [18] <= _1085_[18];
	always @(posedge io_in[12])
		if (_0012_)
			\mchip.chip_design.timing.drop_cnt [19] <= 1'h0;
		else
			\mchip.chip_design.timing.drop_cnt [19] <= _1085_[19];
	always @(posedge io_in[12])
		if (_0012_)
			\mchip.chip_design.timing.drop_cnt [20] <= 1'h0;
		else
			\mchip.chip_design.timing.drop_cnt [20] <= _1085_[20];
	always @(posedge io_in[12])
		if (_0012_)
			\mchip.chip_design.timing.drop_cnt [21] <= 1'h0;
		else
			\mchip.chip_design.timing.drop_cnt [21] <= _1085_[21];
	always @(posedge io_in[12])
		if (_0012_)
			\mchip.chip_design.timing.drop_cnt [22] <= 1'h0;
		else
			\mchip.chip_design.timing.drop_cnt [22] <= _1085_[22];
	always @(posedge io_in[12])
		if (_0012_)
			\mchip.chip_design.timing.drop_cnt [23] <= 1'h0;
		else
			\mchip.chip_design.timing.drop_cnt [23] <= _1085_[23];
	always @(posedge io_in[12])
		if (_0012_)
			\mchip.chip_design.timing.drop_cnt [24] <= 1'h0;
		else
			\mchip.chip_design.timing.drop_cnt [24] <= _1085_[24];
	always @(posedge io_in[12])
		if (_0012_)
			\mchip.chip_design.timing.drop_cnt [25] <= 1'h0;
		else
			\mchip.chip_design.timing.drop_cnt [25] <= _1085_[25];
	always @(posedge io_in[12])
		if (_0012_)
			\mchip.chip_design.timing.drop_cnt [26] <= 1'h0;
		else
			\mchip.chip_design.timing.drop_cnt [26] <= _1085_[26];
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.chip_design.score [0] <= 1'h0;
		else if (\mchip.chip_design.genblk1[0].col.stack_dec )
			\mchip.chip_design.score [0] <= _1072_[0];
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.chip_design.score [1] <= 1'h0;
		else if (\mchip.chip_design.genblk1[0].col.stack_dec )
			\mchip.chip_design.score [1] <= \mchip.chip_design.timing.score_base [3];
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.chip_design.score [2] <= 1'h0;
		else if (\mchip.chip_design.genblk1[0].col.stack_dec )
			\mchip.chip_design.score [2] <= _1073_[2];
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.chip_design.score [3] <= 1'h0;
		else if (\mchip.chip_design.genblk1[0].col.stack_dec )
			\mchip.chip_design.score [3] <= _1073_[3];
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.chip_design.score [4] <= 1'h0;
		else if (\mchip.chip_design.genblk1[0].col.stack_dec )
			\mchip.chip_design.score [4] <= _1073_[4];
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.chip_design.score [5] <= 1'h0;
		else if (\mchip.chip_design.genblk1[0].col.stack_dec )
			\mchip.chip_design.score [5] <= _1073_[5];
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.chip_design.score [6] <= 1'h0;
		else if (\mchip.chip_design.genblk1[0].col.stack_dec )
			\mchip.chip_design.score [6] <= _1073_[6];
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.chip_design.score [7] <= 1'h0;
		else if (\mchip.chip_design.genblk1[0].col.stack_dec )
			\mchip.chip_design.score [7] <= _1073_[7];
	always @(posedge io_in[12]) \mchip.chip_design.new_game_int  <= io_in[1];
	always @(posedge io_in[12]) \mchip.chip_design.new_game  <= \mchip.chip_design.new_game_int ;
	always @(posedge io_in[12]) \mchip.chip_design.drop_int  <= io_in[0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.chip_design.genblk1[7].col.state  <= 1'h0;
		else
			\mchip.chip_design.genblk1[7].col.state  <= \mchip.chip_design.genblk1[7].col.nextState ;
	always @(posedge io_in[12])
		if (_0013_)
			\mchip.chip_design.timing.bounce_cnt [0] <= 1'h0;
		else
			\mchip.chip_design.timing.bounce_cnt [0] <= _1086_[0];
	always @(posedge io_in[12])
		if (_0013_)
			\mchip.chip_design.timing.bounce_cnt [1] <= 1'h0;
		else
			\mchip.chip_design.timing.bounce_cnt [1] <= _1087_[1];
	always @(posedge io_in[12])
		if (_0013_)
			\mchip.chip_design.timing.bounce_cnt [2] <= 1'h0;
		else
			\mchip.chip_design.timing.bounce_cnt [2] <= _1087_[2];
	always @(posedge io_in[12])
		if (_0013_)
			\mchip.chip_design.timing.bounce_cnt [3] <= 1'h0;
		else
			\mchip.chip_design.timing.bounce_cnt [3] <= _1087_[3];
	always @(posedge io_in[12])
		if (_0013_)
			\mchip.chip_design.timing.bounce_cnt [4] <= 1'h0;
		else
			\mchip.chip_design.timing.bounce_cnt [4] <= _1087_[4];
	always @(posedge io_in[12])
		if (_0013_)
			\mchip.chip_design.timing.bounce_cnt [5] <= 1'h0;
		else
			\mchip.chip_design.timing.bounce_cnt [5] <= _1087_[5];
	always @(posedge io_in[12])
		if (_0013_)
			\mchip.chip_design.timing.bounce_cnt [6] <= 1'h0;
		else
			\mchip.chip_design.timing.bounce_cnt [6] <= _1087_[6];
	always @(posedge io_in[12])
		if (_0013_)
			\mchip.chip_design.timing.bounce_cnt [7] <= 1'h0;
		else
			\mchip.chip_design.timing.bounce_cnt [7] <= _1087_[7];
	always @(posedge io_in[12])
		if (_0013_)
			\mchip.chip_design.timing.bounce_cnt [8] <= 1'h0;
		else
			\mchip.chip_design.timing.bounce_cnt [8] <= _1087_[8];
	always @(posedge io_in[12])
		if (_0013_)
			\mchip.chip_design.timing.bounce_cnt [9] <= 1'h0;
		else
			\mchip.chip_design.timing.bounce_cnt [9] <= _1087_[9];
	always @(posedge io_in[12])
		if (_0013_)
			\mchip.chip_design.timing.bounce_cnt [10] <= 1'h0;
		else
			\mchip.chip_design.timing.bounce_cnt [10] <= _1087_[10];
	always @(posedge io_in[12])
		if (_0013_)
			\mchip.chip_design.timing.bounce_cnt [11] <= 1'h0;
		else
			\mchip.chip_design.timing.bounce_cnt [11] <= _1087_[11];
	always @(posedge io_in[12])
		if (_0013_)
			\mchip.chip_design.timing.bounce_cnt [12] <= 1'h0;
		else
			\mchip.chip_design.timing.bounce_cnt [12] <= _1087_[12];
	always @(posedge io_in[12])
		if (_0013_)
			\mchip.chip_design.timing.bounce_cnt [13] <= 1'h0;
		else
			\mchip.chip_design.timing.bounce_cnt [13] <= _1087_[13];
	always @(posedge io_in[12])
		if (_0013_)
			\mchip.chip_design.timing.bounce_cnt [14] <= 1'h0;
		else
			\mchip.chip_design.timing.bounce_cnt [14] <= _1087_[14];
	always @(posedge io_in[12])
		if (_0013_)
			\mchip.chip_design.timing.bounce_cnt [15] <= 1'h0;
		else
			\mchip.chip_design.timing.bounce_cnt [15] <= _1087_[15];
	always @(posedge io_in[12])
		if (_0013_)
			\mchip.chip_design.timing.bounce_cnt [16] <= 1'h0;
		else
			\mchip.chip_design.timing.bounce_cnt [16] <= _1087_[16];
	always @(posedge io_in[12])
		if (_0013_)
			\mchip.chip_design.timing.bounce_cnt [17] <= 1'h0;
		else
			\mchip.chip_design.timing.bounce_cnt [17] <= _1087_[17];
	always @(posedge io_in[12])
		if (_0013_)
			\mchip.chip_design.timing.bounce_cnt [18] <= 1'h0;
		else
			\mchip.chip_design.timing.bounce_cnt [18] <= _1087_[18];
	always @(posedge io_in[12])
		if (_0013_)
			\mchip.chip_design.timing.bounce_cnt [19] <= 1'h0;
		else
			\mchip.chip_design.timing.bounce_cnt [19] <= _1087_[19];
	always @(posedge io_in[12])
		if (_0013_)
			\mchip.chip_design.timing.bounce_cnt [20] <= 1'h0;
		else
			\mchip.chip_design.timing.bounce_cnt [20] <= _1087_[20];
	always @(posedge io_in[12])
		if (_0013_)
			\mchip.chip_design.timing.bounce_cnt [21] <= 1'h0;
		else
			\mchip.chip_design.timing.bounce_cnt [21] <= _1087_[21];
	always @(posedge io_in[12])
		if (_0013_)
			\mchip.chip_design.timing.bounce_cnt [22] <= 1'h0;
		else
			\mchip.chip_design.timing.bounce_cnt [22] <= _1087_[22];
	always @(posedge io_in[12])
		if (_0013_)
			\mchip.chip_design.timing.bounce_cnt [23] <= 1'h0;
		else
			\mchip.chip_design.timing.bounce_cnt [23] <= _1087_[23];
	always @(posedge io_in[12])
		if (_0013_)
			\mchip.chip_design.timing.bounce_cnt [24] <= 1'h0;
		else
			\mchip.chip_design.timing.bounce_cnt [24] <= _1087_[24];
	always @(posedge io_in[12])
		if (_0013_)
			\mchip.chip_design.timing.bounce_cnt [25] <= 1'h0;
		else
			\mchip.chip_design.timing.bounce_cnt [25] <= _1087_[25];
	always @(posedge io_in[12])
		if (_0013_)
			\mchip.chip_design.timing.bounce_cnt [26] <= 1'h0;
		else
			\mchip.chip_design.timing.bounce_cnt [26] <= _1087_[26];
	always @(posedge io_in[12])
		if (_0014_)
			\mchip.chip_design.bounce.state  <= 1'h1;
		else if (_0016_)
			\mchip.chip_design.bounce.state  <= 1'h0;
	always @(posedge io_in[12])
		if (_0019_)
			\mchip.chip_design.genblk1[0].col.drop_pos [0] <= 1'h1;
		else if (_0018_)
			\mchip.chip_design.genblk1[0].col.drop_pos [0] <= _1076_[0];
	always @(posedge io_in[12])
		if (_0019_)
			\mchip.chip_design.genblk1[0].col.drop_pos [1] <= 1'h0;
		else if (_0018_)
			\mchip.chip_design.genblk1[0].col.drop_pos [1] <= _1076_[1];
	always @(posedge io_in[12])
		if (_0019_)
			\mchip.chip_design.genblk1[0].col.drop_pos [2] <= 1'h0;
		else if (_0018_)
			\mchip.chip_design.genblk1[0].col.drop_pos [2] <= _1076_[2];
	always @(posedge io_in[12])
		if (_0019_)
			\mchip.chip_design.genblk1[0].col.drop_pos [3] <= 1'h1;
		else if (_0018_)
			\mchip.chip_design.genblk1[0].col.drop_pos [3] <= _1076_[3];
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.chip_design.genblk1[0].col.stack_pos [0] <= 1'h0;
		else if (_0011_)
			\mchip.chip_design.genblk1[0].col.stack_pos [0] <= _0020_;
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.chip_design.genblk1[0].col.stack_pos [1] <= 1'h0;
		else if (_0011_)
			\mchip.chip_design.genblk1[0].col.stack_pos [1] <= _0021_;
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.chip_design.genblk1[0].col.stack_pos [2] <= 1'h0;
		else if (_0011_)
			\mchip.chip_design.genblk1[0].col.stack_pos [2] <= _0022_;
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.chip_design.genblk1[0].col.stack_pos [3] <= 1'h0;
		else if (_0011_)
			\mchip.chip_design.genblk1[0].col.stack_pos [3] <= _0023_;
	always @(posedge io_in[12])
		if (_0025_)
			\mchip.chip_design.genblk1[1].col.drop_pos [0] <= 1'h1;
		else if (_0024_)
			\mchip.chip_design.genblk1[1].col.drop_pos [0] <= _1077_[0];
	always @(posedge io_in[12])
		if (_0025_)
			\mchip.chip_design.genblk1[1].col.drop_pos [1] <= 1'h0;
		else if (_0024_)
			\mchip.chip_design.genblk1[1].col.drop_pos [1] <= _1077_[1];
	always @(posedge io_in[12])
		if (_0025_)
			\mchip.chip_design.genblk1[1].col.drop_pos [2] <= 1'h0;
		else if (_0024_)
			\mchip.chip_design.genblk1[1].col.drop_pos [2] <= _1077_[2];
	always @(posedge io_in[12])
		if (_0025_)
			\mchip.chip_design.genblk1[1].col.drop_pos [3] <= 1'h1;
		else if (_0024_)
			\mchip.chip_design.genblk1[1].col.drop_pos [3] <= _1077_[3];
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.chip_design.genblk1[1].col.stack_pos [0] <= 1'h0;
		else if (_0010_)
			\mchip.chip_design.genblk1[1].col.stack_pos [0] <= _0026_;
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.chip_design.genblk1[1].col.stack_pos [1] <= 1'h0;
		else if (_0010_)
			\mchip.chip_design.genblk1[1].col.stack_pos [1] <= _0027_;
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.chip_design.genblk1[1].col.stack_pos [2] <= 1'h0;
		else if (_0010_)
			\mchip.chip_design.genblk1[1].col.stack_pos [2] <= _0028_;
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.chip_design.genblk1[1].col.stack_pos [3] <= 1'h0;
		else if (_0010_)
			\mchip.chip_design.genblk1[1].col.stack_pos [3] <= _0029_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.chip_design.genblk1[0].col.state  <= 1'h0;
		else
			\mchip.chip_design.genblk1[0].col.state  <= \mchip.chip_design.genblk1[0].col.nextState ;
	always @(posedge io_in[12])
		if (_0031_)
			\mchip.chip_design.genblk1[2].col.drop_pos [0] <= 1'h1;
		else if (_0030_)
			\mchip.chip_design.genblk1[2].col.drop_pos [0] <= _1078_[0];
	always @(posedge io_in[12])
		if (_0031_)
			\mchip.chip_design.genblk1[2].col.drop_pos [1] <= 1'h0;
		else if (_0030_)
			\mchip.chip_design.genblk1[2].col.drop_pos [1] <= _1078_[1];
	always @(posedge io_in[12])
		if (_0031_)
			\mchip.chip_design.genblk1[2].col.drop_pos [2] <= 1'h0;
		else if (_0030_)
			\mchip.chip_design.genblk1[2].col.drop_pos [2] <= _1078_[2];
	always @(posedge io_in[12])
		if (_0031_)
			\mchip.chip_design.genblk1[2].col.drop_pos [3] <= 1'h1;
		else if (_0030_)
			\mchip.chip_design.genblk1[2].col.drop_pos [3] <= _1078_[3];
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.chip_design.genblk1[2].col.stack_pos [0] <= 1'h0;
		else if (_0009_)
			\mchip.chip_design.genblk1[2].col.stack_pos [0] <= _0032_;
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.chip_design.genblk1[2].col.stack_pos [1] <= 1'h0;
		else if (_0009_)
			\mchip.chip_design.genblk1[2].col.stack_pos [1] <= _0033_;
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.chip_design.genblk1[2].col.stack_pos [2] <= 1'h0;
		else if (_0009_)
			\mchip.chip_design.genblk1[2].col.stack_pos [2] <= _0034_;
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.chip_design.genblk1[2].col.stack_pos [3] <= 1'h0;
		else if (_0009_)
			\mchip.chip_design.genblk1[2].col.stack_pos [3] <= _0035_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.chip_design.genblk1[1].col.state  <= 1'h0;
		else
			\mchip.chip_design.genblk1[1].col.state  <= \mchip.chip_design.genblk1[1].col.nextState ;
	always @(posedge io_in[12])
		if (_0037_)
			\mchip.chip_design.genblk1[3].col.drop_pos [0] <= 1'h1;
		else if (_0036_)
			\mchip.chip_design.genblk1[3].col.drop_pos [0] <= _1079_[0];
	always @(posedge io_in[12])
		if (_0037_)
			\mchip.chip_design.genblk1[3].col.drop_pos [1] <= 1'h0;
		else if (_0036_)
			\mchip.chip_design.genblk1[3].col.drop_pos [1] <= _1079_[1];
	always @(posedge io_in[12])
		if (_0037_)
			\mchip.chip_design.genblk1[3].col.drop_pos [2] <= 1'h0;
		else if (_0036_)
			\mchip.chip_design.genblk1[3].col.drop_pos [2] <= _1079_[2];
	always @(posedge io_in[12])
		if (_0037_)
			\mchip.chip_design.genblk1[3].col.drop_pos [3] <= 1'h1;
		else if (_0036_)
			\mchip.chip_design.genblk1[3].col.drop_pos [3] <= _1079_[3];
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.chip_design.genblk1[3].col.stack_pos [0] <= 1'h0;
		else if (_0008_)
			\mchip.chip_design.genblk1[3].col.stack_pos [0] <= _0038_;
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.chip_design.genblk1[3].col.stack_pos [1] <= 1'h0;
		else if (_0008_)
			\mchip.chip_design.genblk1[3].col.stack_pos [1] <= _0039_;
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.chip_design.genblk1[3].col.stack_pos [2] <= 1'h0;
		else if (_0008_)
			\mchip.chip_design.genblk1[3].col.stack_pos [2] <= _0040_;
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.chip_design.genblk1[3].col.stack_pos [3] <= 1'h0;
		else if (_0008_)
			\mchip.chip_design.genblk1[3].col.stack_pos [3] <= _0041_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.chip_design.genblk1[2].col.state  <= 1'h0;
		else
			\mchip.chip_design.genblk1[2].col.state  <= \mchip.chip_design.genblk1[2].col.nextState ;
	always @(posedge io_in[12])
		if (_0043_)
			\mchip.chip_design.genblk1[4].col.drop_pos [0] <= 1'h1;
		else if (_0042_)
			\mchip.chip_design.genblk1[4].col.drop_pos [0] <= _1080_[0];
	always @(posedge io_in[12])
		if (_0043_)
			\mchip.chip_design.genblk1[4].col.drop_pos [1] <= 1'h0;
		else if (_0042_)
			\mchip.chip_design.genblk1[4].col.drop_pos [1] <= _1080_[1];
	always @(posedge io_in[12])
		if (_0043_)
			\mchip.chip_design.genblk1[4].col.drop_pos [2] <= 1'h0;
		else if (_0042_)
			\mchip.chip_design.genblk1[4].col.drop_pos [2] <= _1080_[2];
	always @(posedge io_in[12])
		if (_0043_)
			\mchip.chip_design.genblk1[4].col.drop_pos [3] <= 1'h1;
		else if (_0042_)
			\mchip.chip_design.genblk1[4].col.drop_pos [3] <= _1080_[3];
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.chip_design.genblk1[4].col.stack_pos [0] <= 1'h0;
		else if (_0007_)
			\mchip.chip_design.genblk1[4].col.stack_pos [0] <= _0044_;
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.chip_design.genblk1[4].col.stack_pos [1] <= 1'h0;
		else if (_0007_)
			\mchip.chip_design.genblk1[4].col.stack_pos [1] <= _0045_;
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.chip_design.genblk1[4].col.stack_pos [2] <= 1'h0;
		else if (_0007_)
			\mchip.chip_design.genblk1[4].col.stack_pos [2] <= _0046_;
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.chip_design.genblk1[4].col.stack_pos [3] <= 1'h0;
		else if (_0007_)
			\mchip.chip_design.genblk1[4].col.stack_pos [3] <= _0047_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.chip_design.genblk1[3].col.state  <= 1'h0;
		else
			\mchip.chip_design.genblk1[3].col.state  <= \mchip.chip_design.genblk1[3].col.nextState ;
	always @(posedge io_in[12])
		if (_0049_)
			\mchip.chip_design.genblk1[5].col.drop_pos [0] <= 1'h1;
		else if (_0048_)
			\mchip.chip_design.genblk1[5].col.drop_pos [0] <= _1081_[0];
	always @(posedge io_in[12])
		if (_0049_)
			\mchip.chip_design.genblk1[5].col.drop_pos [1] <= 1'h0;
		else if (_0048_)
			\mchip.chip_design.genblk1[5].col.drop_pos [1] <= _1081_[1];
	always @(posedge io_in[12])
		if (_0049_)
			\mchip.chip_design.genblk1[5].col.drop_pos [2] <= 1'h0;
		else if (_0048_)
			\mchip.chip_design.genblk1[5].col.drop_pos [2] <= _1081_[2];
	always @(posedge io_in[12])
		if (_0049_)
			\mchip.chip_design.genblk1[5].col.drop_pos [3] <= 1'h1;
		else if (_0048_)
			\mchip.chip_design.genblk1[5].col.drop_pos [3] <= _1081_[3];
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.chip_design.genblk1[5].col.stack_pos [0] <= 1'h0;
		else if (_0006_)
			\mchip.chip_design.genblk1[5].col.stack_pos [0] <= _0050_;
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.chip_design.genblk1[5].col.stack_pos [1] <= 1'h0;
		else if (_0006_)
			\mchip.chip_design.genblk1[5].col.stack_pos [1] <= _0051_;
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.chip_design.genblk1[5].col.stack_pos [2] <= 1'h0;
		else if (_0006_)
			\mchip.chip_design.genblk1[5].col.stack_pos [2] <= _0052_;
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.chip_design.genblk1[5].col.stack_pos [3] <= 1'h0;
		else if (_0006_)
			\mchip.chip_design.genblk1[5].col.stack_pos [3] <= _0053_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.chip_design.genblk1[4].col.state  <= 1'h0;
		else
			\mchip.chip_design.genblk1[4].col.state  <= \mchip.chip_design.genblk1[4].col.nextState ;
	always @(posedge io_in[12])
		if (_0055_)
			\mchip.chip_design.genblk1[6].col.drop_pos [0] <= 1'h1;
		else if (_0054_)
			\mchip.chip_design.genblk1[6].col.drop_pos [0] <= _1082_[0];
	always @(posedge io_in[12])
		if (_0055_)
			\mchip.chip_design.genblk1[6].col.drop_pos [1] <= 1'h0;
		else if (_0054_)
			\mchip.chip_design.genblk1[6].col.drop_pos [1] <= _1082_[1];
	always @(posedge io_in[12])
		if (_0055_)
			\mchip.chip_design.genblk1[6].col.drop_pos [2] <= 1'h0;
		else if (_0054_)
			\mchip.chip_design.genblk1[6].col.drop_pos [2] <= _1082_[2];
	always @(posedge io_in[12])
		if (_0055_)
			\mchip.chip_design.genblk1[6].col.drop_pos [3] <= 1'h1;
		else if (_0054_)
			\mchip.chip_design.genblk1[6].col.drop_pos [3] <= _1082_[3];
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.chip_design.genblk1[6].col.stack_pos [0] <= 1'h0;
		else if (_0005_)
			\mchip.chip_design.genblk1[6].col.stack_pos [0] <= _0056_;
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.chip_design.genblk1[6].col.stack_pos [1] <= 1'h0;
		else if (_0005_)
			\mchip.chip_design.genblk1[6].col.stack_pos [1] <= _0057_;
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.chip_design.genblk1[6].col.stack_pos [2] <= 1'h0;
		else if (_0005_)
			\mchip.chip_design.genblk1[6].col.stack_pos [2] <= _0058_;
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.chip_design.genblk1[6].col.stack_pos [3] <= 1'h0;
		else if (_0005_)
			\mchip.chip_design.genblk1[6].col.stack_pos [3] <= _0059_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.chip_design.genblk1[5].col.state  <= 1'h0;
		else
			\mchip.chip_design.genblk1[5].col.state  <= \mchip.chip_design.genblk1[5].col.nextState ;
	always @(posedge io_in[12])
		if (_0061_)
			\mchip.chip_design.genblk1[7].col.drop_pos [0] <= 1'h1;
		else if (_0060_)
			\mchip.chip_design.genblk1[7].col.drop_pos [0] <= _1083_[0];
	always @(posedge io_in[12])
		if (_0061_)
			\mchip.chip_design.genblk1[7].col.drop_pos [1] <= 1'h0;
		else if (_0060_)
			\mchip.chip_design.genblk1[7].col.drop_pos [1] <= _1083_[1];
	always @(posedge io_in[12])
		if (_0061_)
			\mchip.chip_design.genblk1[7].col.drop_pos [2] <= 1'h0;
		else if (_0060_)
			\mchip.chip_design.genblk1[7].col.drop_pos [2] <= _1083_[2];
	always @(posedge io_in[12])
		if (_0061_)
			\mchip.chip_design.genblk1[7].col.drop_pos [3] <= 1'h1;
		else if (_0060_)
			\mchip.chip_design.genblk1[7].col.drop_pos [3] <= _1083_[3];
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.chip_design.genblk1[7].col.stack_pos [0] <= 1'h0;
		else if (_0004_)
			\mchip.chip_design.genblk1[7].col.stack_pos [0] <= _0062_;
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.chip_design.genblk1[7].col.stack_pos [1] <= 1'h0;
		else if (_0004_)
			\mchip.chip_design.genblk1[7].col.stack_pos [1] <= _0063_;
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.chip_design.genblk1[7].col.stack_pos [2] <= 1'h0;
		else if (_0004_)
			\mchip.chip_design.genblk1[7].col.stack_pos [2] <= _0064_;
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.chip_design.genblk1[7].col.stack_pos [3] <= 1'h0;
		else if (_0004_)
			\mchip.chip_design.genblk1[7].col.stack_pos [3] <= _0065_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.chip_design.genblk1[6].col.state  <= 1'h0;
		else
			\mchip.chip_design.genblk1[6].col.state  <= \mchip.chip_design.genblk1[6].col.nextState ;
	always @(posedge io_in[12]) \mchip.chip_design.state [0] <= _0000_;
	always @(posedge io_in[12]) \mchip.chip_design.state [1] <= _0001_;
	always @(posedge io_in[12]) \mchip.chip_design.state [2] <= _0002_;
	always @(posedge io_in[12]) \mchip.chip_design.state [3] <= _0003_;
	assign _1072_[7:1] = \mchip.chip_design.score [7:1];
	assign _1073_[1:0] = {\mchip.chip_design.timing.score_base [3], _1072_[0]};
	assign _1074_[31:1] = 31'h7ffffffc;
	assign _1075_[0] = _1074_[0];
	assign _1084_[26:1] = \mchip.chip_design.timing.drop_cnt [26:1];
	assign _1085_[0] = _1084_[0];
	assign _1086_[26:1] = \mchip.chip_design.timing.bounce_cnt [26:1];
	assign _1087_[0] = _1086_[0];
	assign {io_out[13:12], io_out[3:0]} = {2'h0, \mchip.chip_design.bounce.bounce_pos , \mchip.chip_design.bounce.game_running };
	assign \mchip.chip_design.bounce.clock  = io_in[12];
	assign \mchip.chip_design.bounce.reset  = io_in[13];
	assign \mchip.chip_design.bounce_pos  = \mchip.chip_design.bounce.bounce_pos ;
	assign \mchip.chip_design.clock  = io_in[12];
	assign \mchip.chip_design.drop_btn  = io_in[0];
	assign \mchip.chip_design.drop_pos[0]  = \mchip.chip_design.genblk1[0].col.drop_pos ;
	assign \mchip.chip_design.drop_pos[1]  = \mchip.chip_design.genblk1[1].col.drop_pos ;
	assign \mchip.chip_design.drop_pos[2]  = \mchip.chip_design.genblk1[2].col.drop_pos ;
	assign \mchip.chip_design.drop_pos[3]  = \mchip.chip_design.genblk1[3].col.drop_pos ;
	assign \mchip.chip_design.drop_pos[4]  = \mchip.chip_design.genblk1[4].col.drop_pos ;
	assign \mchip.chip_design.drop_pos[5]  = \mchip.chip_design.genblk1[5].col.drop_pos ;
	assign \mchip.chip_design.drop_pos[6]  = \mchip.chip_design.genblk1[6].col.drop_pos ;
	assign \mchip.chip_design.drop_pos[7]  = \mchip.chip_design.genblk1[7].col.drop_pos ;
	assign \mchip.chip_design.game_running  = \mchip.chip_design.bounce.game_running ;
	assign \mchip.chip_design.genblk1[0].col.clock  = io_in[12];
	assign \mchip.chip_design.genblk1[0].col.reset  = io_in[13];
	assign \mchip.chip_design.genblk1[1].col.clock  = io_in[12];
	assign \mchip.chip_design.genblk1[1].col.reset  = io_in[13];
	assign \mchip.chip_design.genblk1[1].col.stack_dec  = \mchip.chip_design.genblk1[0].col.stack_dec ;
	assign \mchip.chip_design.genblk1[2].col.clock  = io_in[12];
	assign \mchip.chip_design.genblk1[2].col.reset  = io_in[13];
	assign \mchip.chip_design.genblk1[2].col.stack_dec  = \mchip.chip_design.genblk1[0].col.stack_dec ;
	assign \mchip.chip_design.genblk1[3].col.clock  = io_in[12];
	assign \mchip.chip_design.genblk1[3].col.reset  = io_in[13];
	assign \mchip.chip_design.genblk1[3].col.stack_dec  = \mchip.chip_design.genblk1[0].col.stack_dec ;
	assign \mchip.chip_design.genblk1[4].col.clock  = io_in[12];
	assign \mchip.chip_design.genblk1[4].col.reset  = io_in[13];
	assign \mchip.chip_design.genblk1[4].col.stack_dec  = \mchip.chip_design.genblk1[0].col.stack_dec ;
	assign \mchip.chip_design.genblk1[5].col.clock  = io_in[12];
	assign \mchip.chip_design.genblk1[5].col.reset  = io_in[13];
	assign \mchip.chip_design.genblk1[5].col.stack_dec  = \mchip.chip_design.genblk1[0].col.stack_dec ;
	assign \mchip.chip_design.genblk1[6].col.clock  = io_in[12];
	assign \mchip.chip_design.genblk1[6].col.reset  = io_in[13];
	assign \mchip.chip_design.genblk1[6].col.stack_dec  = \mchip.chip_design.genblk1[0].col.stack_dec ;
	assign \mchip.chip_design.genblk1[7].col.clock  = io_in[12];
	assign \mchip.chip_design.genblk1[7].col.reset  = io_in[13];
	assign \mchip.chip_design.genblk1[7].col.stack_dec  = \mchip.chip_design.genblk1[0].col.stack_dec ;
	assign \mchip.chip_design.initial_game_speed  = io_in[11:6];
	assign \mchip.chip_design.inputs  = io_in[11:0];
	assign \mchip.chip_design.new_game_btn  = io_in[1];
	assign \mchip.chip_design.outputs  = {io_out[11:4], \mchip.chip_design.bounce.bounce_pos , \mchip.chip_design.bounce.game_running };
	assign \mchip.chip_design.reset  = io_in[13];
	assign \mchip.chip_design.stack_dec  = \mchip.chip_design.genblk1[0].col.stack_dec ;
	assign \mchip.chip_design.stack_pos[0]  = \mchip.chip_design.genblk1[0].col.stack_pos ;
	assign \mchip.chip_design.stack_pos[1]  = \mchip.chip_design.genblk1[1].col.stack_pos ;
	assign \mchip.chip_design.stack_pos[2]  = \mchip.chip_design.genblk1[2].col.stack_pos ;
	assign \mchip.chip_design.stack_pos[3]  = \mchip.chip_design.genblk1[3].col.stack_pos ;
	assign \mchip.chip_design.stack_pos[4]  = \mchip.chip_design.genblk1[4].col.stack_pos ;
	assign \mchip.chip_design.stack_pos[5]  = \mchip.chip_design.genblk1[5].col.stack_pos ;
	assign \mchip.chip_design.stack_pos[6]  = \mchip.chip_design.genblk1[6].col.stack_pos ;
	assign \mchip.chip_design.stack_pos[7]  = \mchip.chip_design.genblk1[7].col.stack_pos ;
	assign \mchip.chip_design.timing.bounce_max_val  = {24'h000000, \mchip.chip_design.score [0], 2'h0};
	assign \mchip.chip_design.timing.clock  = io_in[12];
	assign \mchip.chip_design.timing.drop_max_val  = 27'h0001388;
	assign \mchip.chip_design.timing.initial_game_speed  = io_in[11:6];
	assign \mchip.chip_design.timing.initial_game_speed_base  = {23'h000000, io_in[6], 3'h0};
	assign \mchip.chip_design.timing.reset  = io_in[13];
	assign \mchip.chip_design.timing.score  = \mchip.chip_design.score ;
	assign {\mchip.chip_design.timing.score_base [26:4], \mchip.chip_design.timing.score_base [2:0]} = {23'h000000, \mchip.chip_design.score [0], 2'h0};
	assign \mchip.chip_design.update_request_location  = io_in[5:2];
	assign \mchip.chip_design.update_value  = io_out[11:4];
	assign \mchip.clock  = io_in[12];
	assign \mchip.io_in  = io_in[11:0];
	assign \mchip.io_out  = {io_out[11:4], \mchip.chip_design.bounce.bounce_pos , \mchip.chip_design.bounce.game_running };
	assign \mchip.reset  = io_in[13];
endmodule
module d18_nikhildj_mac (
	io_in,
	io_out
);
	wire _000_;
	wire _001_;
	wire _002_;
	wire _003_;
	wire _004_;
	wire _005_;
	wire _006_;
	wire _007_;
	wire _008_;
	wire _009_;
	wire _010_;
	wire _011_;
	wire _012_;
	wire _013_;
	wire _014_;
	wire _015_;
	wire _016_;
	wire _017_;
	wire _018_;
	wire _019_;
	wire _020_;
	wire _021_;
	wire _022_;
	wire _023_;
	wire _024_;
	wire _025_;
	wire _026_;
	wire _027_;
	wire _028_;
	wire _029_;
	wire _030_;
	wire _031_;
	wire _032_;
	wire _033_;
	wire _034_;
	wire _035_;
	wire _036_;
	wire _037_;
	wire _038_;
	wire _039_;
	wire _040_;
	wire _041_;
	wire _042_;
	wire _043_;
	wire _044_;
	wire _045_;
	wire _046_;
	wire _047_;
	wire _048_;
	wire _049_;
	wire _050_;
	wire _051_;
	wire _052_;
	wire _053_;
	wire _054_;
	wire _055_;
	wire _056_;
	wire _057_;
	wire _058_;
	wire _059_;
	wire _060_;
	wire _061_;
	wire _062_;
	wire _063_;
	wire _064_;
	wire _065_;
	wire _066_;
	wire _067_;
	wire _068_;
	wire _069_;
	wire _070_;
	wire _071_;
	wire _072_;
	wire _073_;
	wire _074_;
	wire _075_;
	wire _076_;
	wire _077_;
	wire _078_;
	wire _079_;
	wire _080_;
	wire _081_;
	wire _082_;
	wire _083_;
	wire _084_;
	wire _085_;
	wire _086_;
	wire _087_;
	wire _088_;
	wire _089_;
	wire _090_;
	wire _091_;
	wire _092_;
	wire _093_;
	wire _094_;
	wire _095_;
	wire _096_;
	wire _097_;
	wire _098_;
	wire _099_;
	wire _100_;
	wire _101_;
	wire _102_;
	wire _103_;
	wire _104_;
	wire _105_;
	wire _106_;
	wire _107_;
	wire _108_;
	wire _109_;
	wire _110_;
	wire _111_;
	wire _112_;
	wire _113_;
	wire _114_;
	wire _115_;
	wire _116_;
	wire _117_;
	wire _118_;
	wire _119_;
	wire _120_;
	wire _121_;
	wire _122_;
	wire _123_;
	wire _124_;
	wire _125_;
	wire _126_;
	wire _127_;
	wire _128_;
	wire _129_;
	wire _130_;
	wire _131_;
	wire _132_;
	wire _133_;
	wire _134_;
	wire _135_;
	wire _136_;
	wire _137_;
	wire _138_;
	wire _139_;
	wire _140_;
	wire _141_;
	wire _142_;
	wire _143_;
	wire _144_;
	wire _145_;
	wire _146_;
	wire _147_;
	wire _148_;
	wire _149_;
	wire _150_;
	wire _151_;
	wire _152_;
	wire _153_;
	wire _154_;
	wire _155_;
	wire _156_;
	wire _157_;
	wire _158_;
	wire _159_;
	wire _160_;
	wire _161_;
	wire _162_;
	wire _163_;
	wire _164_;
	wire _165_;
	wire _166_;
	wire _167_;
	wire _168_;
	wire _169_;
	wire _170_;
	wire _171_;
	wire _172_;
	wire _173_;
	wire _174_;
	wire _175_;
	wire _176_;
	wire _177_;
	wire _178_;
	wire _179_;
	wire _180_;
	wire _181_;
	wire _182_;
	wire _183_;
	wire _184_;
	wire _185_;
	wire _186_;
	wire _187_;
	wire _188_;
	wire _189_;
	wire _190_;
	wire _191_;
	wire _192_;
	wire _193_;
	wire _194_;
	wire _195_;
	wire _196_;
	wire _197_;
	wire _198_;
	wire _199_;
	wire _200_;
	wire _201_;
	wire _202_;
	wire _203_;
	wire _204_;
	wire _205_;
	wire _206_;
	wire _207_;
	wire _208_;
	wire _209_;
	wire _210_;
	wire _211_;
	wire _212_;
	wire _213_;
	wire _214_;
	wire _215_;
	wire _216_;
	wire _217_;
	wire _218_;
	wire _219_;
	wire _220_;
	wire _221_;
	wire _222_;
	wire _223_;
	wire _224_;
	wire _225_;
	wire _226_;
	wire _227_;
	wire _228_;
	wire _229_;
	wire _230_;
	wire _231_;
	wire _232_;
	wire _233_;
	wire _234_;
	wire _235_;
	wire _236_;
	wire _237_;
	wire _238_;
	wire _239_;
	wire _240_;
	wire _241_;
	wire _242_;
	wire _243_;
	wire _244_;
	wire _245_;
	wire _246_;
	wire _247_;
	wire _248_;
	wire _249_;
	wire _250_;
	wire _251_;
	wire _252_;
	input wire [13:0] io_in;
	output wire [13:0] io_out;
	wire \mchip.Begin_mul ;
	wire \mchip.End_mul ;
	wire \mchip.Finish ;
	wire \mchip.Load_op ;
	wire \mchip.START ;
	reg \mchip._Finish ;
	wire \mchip.aa.accmulate.dff_gen[0].d2.D ;
	reg \mchip.aa.accmulate.dff_gen[0].d2.Q ;
	wire \mchip.aa.accmulate.dff_gen[10].d2.D ;
	reg \mchip.aa.accmulate.dff_gen[10].d2.Q ;
	wire \mchip.aa.accmulate.dff_gen[11].d2.D ;
	reg \mchip.aa.accmulate.dff_gen[11].d2.Q ;
	wire \mchip.aa.accmulate.dff_gen[12].d2.D ;
	reg \mchip.aa.accmulate.dff_gen[12].d2.Q ;
	wire \mchip.aa.accmulate.dff_gen[13].d2.D ;
	reg \mchip.aa.accmulate.dff_gen[13].d2.Q ;
	wire \mchip.aa.accmulate.dff_gen[14].d2.D ;
	reg \mchip.aa.accmulate.dff_gen[14].d2.Q ;
	wire \mchip.aa.accmulate.dff_gen[15].d2.D ;
	reg \mchip.aa.accmulate.dff_gen[15].d2.Q ;
	reg \mchip.aa.accmulate.dff_gen[16].d2.Q ;
	reg \mchip.aa.accmulate.dff_gen[17].d2.Q ;
	reg \mchip.aa.accmulate.dff_gen[18].d2.Q ;
	reg \mchip.aa.accmulate.dff_gen[19].d2.Q ;
	wire \mchip.aa.accmulate.dff_gen[1].d2.D ;
	reg \mchip.aa.accmulate.dff_gen[1].d2.Q ;
	wire \mchip.aa.accmulate.dff_gen[2].d2.D ;
	reg \mchip.aa.accmulate.dff_gen[2].d2.Q ;
	wire \mchip.aa.accmulate.dff_gen[3].d2.D ;
	reg \mchip.aa.accmulate.dff_gen[3].d2.Q ;
	wire \mchip.aa.accmulate.dff_gen[4].d2.D ;
	reg \mchip.aa.accmulate.dff_gen[4].d2.Q ;
	wire \mchip.aa.accmulate.dff_gen[5].d2.D ;
	reg \mchip.aa.accmulate.dff_gen[5].d2.Q ;
	wire \mchip.aa.accmulate.dff_gen[6].d2.D ;
	reg \mchip.aa.accmulate.dff_gen[6].d2.Q ;
	wire \mchip.aa.accmulate.dff_gen[7].d2.D ;
	reg \mchip.aa.accmulate.dff_gen[7].d2.Q ;
	wire \mchip.aa.accmulate.dff_gen[8].d2.D ;
	reg \mchip.aa.accmulate.dff_gen[8].d2.Q ;
	wire \mchip.aa.accmulate.dff_gen[9].d2.D ;
	reg \mchip.aa.accmulate.dff_gen[9].d2.Q ;
	wire [19:0] \mchip.aa.accmulate.in ;
	wire [19:0] \mchip.aa.accmulate.out ;
	wire [19:0] \mchip.aa.accmulate.temp_out ;
	wire \mchip.aa.add ;
	wire [19:0] \mchip.aa.add_in ;
	wire [19:0] \mchip.aa.add_out ;
	wire [3:0] \mchip.aa.adder.S0.S0.a ;
	wire [3:0] \mchip.aa.adder.S0.S0.b ;
	wire \mchip.aa.adder.S0.S0.carry_in ;
	wire \mchip.aa.adder.S0.S0.fa0.a ;
	wire \mchip.aa.adder.S0.S0.fa0.b ;
	wire \mchip.aa.adder.S0.S0.fa0.carry_in ;
	wire \mchip.aa.adder.S0.S0.fa0.sum ;
	wire \mchip.aa.adder.S0.S0.fa0.w1 ;
	wire \mchip.aa.adder.S0.S0.fa0.w3 ;
	wire \mchip.aa.adder.S0.S0.fa1.a ;
	wire \mchip.aa.adder.S0.S0.fa1.b ;
	wire \mchip.aa.adder.S0.S0.fa1.sum ;
	wire \mchip.aa.adder.S0.S0.fa2.a ;
	wire \mchip.aa.adder.S0.S0.fa2.b ;
	wire \mchip.aa.adder.S0.S0.fa2.sum ;
	wire \mchip.aa.adder.S0.S0.fa3.a ;
	wire \mchip.aa.adder.S0.S0.fa3.b ;
	wire \mchip.aa.adder.S0.S0.fa3.sum ;
	wire [3:0] \mchip.aa.adder.S0.S0.sum ;
	wire [3:0] \mchip.aa.adder.S0.S1.a ;
	wire [3:0] \mchip.aa.adder.S0.S1.b ;
	wire \mchip.aa.adder.S0.S1.carry_in ;
	wire \mchip.aa.adder.S0.S1.fa0.a ;
	wire \mchip.aa.adder.S0.S1.fa0.b ;
	wire \mchip.aa.adder.S0.S1.fa0.carry_in ;
	wire \mchip.aa.adder.S0.S1.fa1.a ;
	wire \mchip.aa.adder.S0.S1.fa1.b ;
	wire \mchip.aa.adder.S0.S1.fa2.a ;
	wire \mchip.aa.adder.S0.S1.fa2.b ;
	wire \mchip.aa.adder.S0.S1.fa3.a ;
	wire \mchip.aa.adder.S0.S1.fa3.b ;
	wire [3:0] \mchip.aa.adder.S0.SUM0 ;
	wire [3:0] \mchip.aa.adder.S0.a ;
	wire [3:0] \mchip.aa.adder.S0.b ;
	wire \mchip.aa.adder.S0.carry_in ;
	wire [3:0] \mchip.aa.adder.S0.sum ;
	wire [3:0] \mchip.aa.adder.S1.S0.a ;
	wire [3:0] \mchip.aa.adder.S1.S0.b ;
	wire \mchip.aa.adder.S1.S0.carry_in ;
	wire \mchip.aa.adder.S1.S0.fa0.a ;
	wire \mchip.aa.adder.S1.S0.fa0.b ;
	wire \mchip.aa.adder.S1.S0.fa0.carry_in ;
	wire \mchip.aa.adder.S1.S0.fa0.w3 ;
	wire \mchip.aa.adder.S1.S0.fa1.a ;
	wire \mchip.aa.adder.S1.S0.fa1.b ;
	wire \mchip.aa.adder.S1.S0.fa2.a ;
	wire \mchip.aa.adder.S1.S0.fa2.b ;
	wire \mchip.aa.adder.S1.S0.fa3.a ;
	wire \mchip.aa.adder.S1.S0.fa3.b ;
	wire [3:0] \mchip.aa.adder.S1.S0.sum ;
	wire [3:0] \mchip.aa.adder.S1.S1.a ;
	wire [3:0] \mchip.aa.adder.S1.S1.b ;
	wire \mchip.aa.adder.S1.S1.carry_in ;
	wire \mchip.aa.adder.S1.S1.fa0.a ;
	wire \mchip.aa.adder.S1.S1.fa0.b ;
	wire \mchip.aa.adder.S1.S1.fa0.carry_in ;
	wire \mchip.aa.adder.S1.S1.fa1.a ;
	wire \mchip.aa.adder.S1.S1.fa1.b ;
	wire \mchip.aa.adder.S1.S1.fa2.a ;
	wire \mchip.aa.adder.S1.S1.fa2.b ;
	wire \mchip.aa.adder.S1.S1.fa3.a ;
	wire \mchip.aa.adder.S1.S1.fa3.b ;
	wire [3:0] \mchip.aa.adder.S1.S1.sum ;
	wire [3:0] \mchip.aa.adder.S1.SUM0 ;
	wire [3:0] \mchip.aa.adder.S1.SUM1 ;
	wire [3:0] \mchip.aa.adder.S1.a ;
	wire [3:0] \mchip.aa.adder.S1.b ;
	wire [3:0] \mchip.aa.adder.S1.sum ;
	wire [3:0] \mchip.aa.adder.S2.S0.a ;
	wire [3:0] \mchip.aa.adder.S2.S0.b ;
	wire \mchip.aa.adder.S2.S0.carry_in ;
	wire \mchip.aa.adder.S2.S0.fa0.a ;
	wire \mchip.aa.adder.S2.S0.fa0.b ;
	wire \mchip.aa.adder.S2.S0.fa0.carry_in ;
	wire \mchip.aa.adder.S2.S0.fa0.w3 ;
	wire \mchip.aa.adder.S2.S0.fa1.a ;
	wire \mchip.aa.adder.S2.S0.fa1.b ;
	wire \mchip.aa.adder.S2.S0.fa2.a ;
	wire \mchip.aa.adder.S2.S0.fa2.b ;
	wire \mchip.aa.adder.S2.S0.fa3.a ;
	wire \mchip.aa.adder.S2.S0.fa3.b ;
	wire [3:0] \mchip.aa.adder.S2.S0.sum ;
	wire [3:0] \mchip.aa.adder.S2.S1.a ;
	wire [3:0] \mchip.aa.adder.S2.S1.b ;
	wire \mchip.aa.adder.S2.S1.carry_in ;
	wire \mchip.aa.adder.S2.S1.fa0.a ;
	wire \mchip.aa.adder.S2.S1.fa0.b ;
	wire \mchip.aa.adder.S2.S1.fa0.carry_in ;
	wire \mchip.aa.adder.S2.S1.fa1.a ;
	wire \mchip.aa.adder.S2.S1.fa1.b ;
	wire \mchip.aa.adder.S2.S1.fa2.a ;
	wire \mchip.aa.adder.S2.S1.fa2.b ;
	wire \mchip.aa.adder.S2.S1.fa3.a ;
	wire \mchip.aa.adder.S2.S1.fa3.b ;
	wire [3:0] \mchip.aa.adder.S2.S1.sum ;
	wire [3:0] \mchip.aa.adder.S2.SUM0 ;
	wire [3:0] \mchip.aa.adder.S2.SUM1 ;
	wire [3:0] \mchip.aa.adder.S2.a ;
	wire [3:0] \mchip.aa.adder.S2.b ;
	wire [3:0] \mchip.aa.adder.S2.sum ;
	wire [3:0] \mchip.aa.adder.S3.S0.a ;
	wire [3:0] \mchip.aa.adder.S3.S0.b ;
	wire \mchip.aa.adder.S3.S0.carry_in ;
	wire \mchip.aa.adder.S3.S0.fa0.a ;
	wire \mchip.aa.adder.S3.S0.fa0.b ;
	wire \mchip.aa.adder.S3.S0.fa0.carry_in ;
	wire \mchip.aa.adder.S3.S0.fa0.w3 ;
	wire \mchip.aa.adder.S3.S0.fa1.a ;
	wire \mchip.aa.adder.S3.S0.fa1.b ;
	wire \mchip.aa.adder.S3.S0.fa2.a ;
	wire \mchip.aa.adder.S3.S0.fa2.b ;
	wire \mchip.aa.adder.S3.S0.fa3.a ;
	wire \mchip.aa.adder.S3.S0.fa3.b ;
	wire [3:0] \mchip.aa.adder.S3.S0.sum ;
	wire [3:0] \mchip.aa.adder.S3.S1.a ;
	wire [3:0] \mchip.aa.adder.S3.S1.b ;
	wire \mchip.aa.adder.S3.S1.carry_in ;
	wire \mchip.aa.adder.S3.S1.fa0.a ;
	wire \mchip.aa.adder.S3.S1.fa0.b ;
	wire \mchip.aa.adder.S3.S1.fa0.carry_in ;
	wire \mchip.aa.adder.S3.S1.fa1.a ;
	wire \mchip.aa.adder.S3.S1.fa1.b ;
	wire \mchip.aa.adder.S3.S1.fa2.a ;
	wire \mchip.aa.adder.S3.S1.fa2.b ;
	wire \mchip.aa.adder.S3.S1.fa3.a ;
	wire \mchip.aa.adder.S3.S1.fa3.b ;
	wire [3:0] \mchip.aa.adder.S3.S1.sum ;
	wire [3:0] \mchip.aa.adder.S3.SUM0 ;
	wire [3:0] \mchip.aa.adder.S3.SUM1 ;
	wire [3:0] \mchip.aa.adder.S3.a ;
	wire [3:0] \mchip.aa.adder.S3.b ;
	wire \mchip.aa.adder.S3.carry_out ;
	wire [3:0] \mchip.aa.adder.S3.sum ;
	wire [3:0] \mchip.aa.adder.S4.S0.a ;
	wire [3:0] \mchip.aa.adder.S4.S0.b ;
	wire \mchip.aa.adder.S4.S0.carry_in ;
	wire \mchip.aa.adder.S4.S0.carry_out ;
	wire \mchip.aa.adder.S4.S0.fa0.a ;
	wire \mchip.aa.adder.S4.S0.fa0.b ;
	wire \mchip.aa.adder.S4.S0.fa0.carry_in ;
	wire \mchip.aa.adder.S4.S0.fa0.carry_out ;
	wire \mchip.aa.adder.S4.S0.fa0.sum ;
	wire \mchip.aa.adder.S4.S0.fa0.w1 ;
	wire \mchip.aa.adder.S4.S0.fa0.w2 ;
	wire \mchip.aa.adder.S4.S0.fa0.w3 ;
	wire \mchip.aa.adder.S4.S0.fa1.a ;
	wire \mchip.aa.adder.S4.S0.fa1.b ;
	wire \mchip.aa.adder.S4.S0.fa1.carry_in ;
	wire \mchip.aa.adder.S4.S0.fa1.carry_out ;
	wire \mchip.aa.adder.S4.S0.fa1.sum ;
	wire \mchip.aa.adder.S4.S0.fa1.w1 ;
	wire \mchip.aa.adder.S4.S0.fa1.w2 ;
	wire \mchip.aa.adder.S4.S0.fa1.w3 ;
	wire \mchip.aa.adder.S4.S0.fa2.a ;
	wire \mchip.aa.adder.S4.S0.fa2.b ;
	wire \mchip.aa.adder.S4.S0.fa2.carry_in ;
	wire \mchip.aa.adder.S4.S0.fa2.carry_out ;
	wire \mchip.aa.adder.S4.S0.fa2.sum ;
	wire \mchip.aa.adder.S4.S0.fa2.w1 ;
	wire \mchip.aa.adder.S4.S0.fa2.w2 ;
	wire \mchip.aa.adder.S4.S0.fa2.w3 ;
	wire \mchip.aa.adder.S4.S0.fa3.a ;
	wire \mchip.aa.adder.S4.S0.fa3.b ;
	wire \mchip.aa.adder.S4.S0.fa3.carry_in ;
	wire \mchip.aa.adder.S4.S0.fa3.carry_out ;
	wire \mchip.aa.adder.S4.S0.fa3.sum ;
	wire \mchip.aa.adder.S4.S0.fa3.w1 ;
	wire \mchip.aa.adder.S4.S0.fa3.w2 ;
	wire \mchip.aa.adder.S4.S0.fa3.w3 ;
	wire [3:0] \mchip.aa.adder.S4.S0.sum ;
	wire \mchip.aa.adder.S4.S0.w1 ;
	wire \mchip.aa.adder.S4.S0.w2 ;
	wire \mchip.aa.adder.S4.S0.w3 ;
	wire [3:0] \mchip.aa.adder.S4.S1.a ;
	wire [3:0] \mchip.aa.adder.S4.S1.b ;
	wire \mchip.aa.adder.S4.S1.carry_in ;
	wire \mchip.aa.adder.S4.S1.fa0.a ;
	wire \mchip.aa.adder.S4.S1.fa0.b ;
	wire \mchip.aa.adder.S4.S1.fa0.carry_in ;
	wire \mchip.aa.adder.S4.S1.fa0.carry_out ;
	wire \mchip.aa.adder.S4.S1.fa0.sum ;
	wire \mchip.aa.adder.S4.S1.fa0.w1 ;
	wire \mchip.aa.adder.S4.S1.fa0.w2 ;
	wire \mchip.aa.adder.S4.S1.fa0.w3 ;
	wire \mchip.aa.adder.S4.S1.fa1.a ;
	wire \mchip.aa.adder.S4.S1.fa1.b ;
	wire \mchip.aa.adder.S4.S1.fa1.carry_in ;
	wire \mchip.aa.adder.S4.S1.fa1.sum ;
	wire \mchip.aa.adder.S4.S1.fa1.w1 ;
	wire \mchip.aa.adder.S4.S1.fa1.w2 ;
	wire \mchip.aa.adder.S4.S1.fa2.a ;
	wire \mchip.aa.adder.S4.S1.fa2.b ;
	wire \mchip.aa.adder.S4.S1.fa2.sum ;
	wire \mchip.aa.adder.S4.S1.fa2.w1 ;
	wire \mchip.aa.adder.S4.S1.fa2.w2 ;
	wire \mchip.aa.adder.S4.S1.fa3.a ;
	wire \mchip.aa.adder.S4.S1.fa3.b ;
	wire \mchip.aa.adder.S4.S1.fa3.sum ;
	wire \mchip.aa.adder.S4.S1.fa3.w1 ;
	wire \mchip.aa.adder.S4.S1.fa3.w2 ;
	wire [3:0] \mchip.aa.adder.S4.S1.sum ;
	wire \mchip.aa.adder.S4.S1.w1 ;
	wire [3:0] \mchip.aa.adder.S4.SUM0 ;
	wire [3:0] \mchip.aa.adder.S4.SUM1 ;
	wire [3:0] \mchip.aa.adder.S4.a ;
	wire [3:0] \mchip.aa.adder.S4.b ;
	wire \mchip.aa.adder.S4.carry0 ;
	wire \mchip.aa.adder.S4.carry_in ;
	wire \mchip.aa.adder.S4.carry_out ;
	wire [19:0] \mchip.aa.adder.a ;
	wire [19:0] \mchip.aa.adder.b ;
	wire \mchip.aa.adder.carry_in ;
	wire \mchip.aa.adder.carry_out ;
	wire [19:0] \mchip.aa.adder.sum ;
	wire \mchip.aa.adder.temp_carry4 ;
	wire \mchip.aa.i0.add ;
	wire \mchip.aa.i0.dff_gen[0].d2.D ;
	reg \mchip.aa.i0.dff_gen[0].d2.Q ;
	wire \mchip.aa.i0.dff_gen[0].d2.clk ;
	wire \mchip.aa.i0.dff_gen[10].d2.D ;
	reg \mchip.aa.i0.dff_gen[10].d2.Q ;
	wire \mchip.aa.i0.dff_gen[10].d2.clk ;
	wire \mchip.aa.i0.dff_gen[11].d2.D ;
	reg \mchip.aa.i0.dff_gen[11].d2.Q ;
	wire \mchip.aa.i0.dff_gen[11].d2.clk ;
	wire \mchip.aa.i0.dff_gen[12].d2.D ;
	reg \mchip.aa.i0.dff_gen[12].d2.Q ;
	wire \mchip.aa.i0.dff_gen[12].d2.clk ;
	wire \mchip.aa.i0.dff_gen[13].d2.D ;
	reg \mchip.aa.i0.dff_gen[13].d2.Q ;
	wire \mchip.aa.i0.dff_gen[13].d2.clk ;
	wire \mchip.aa.i0.dff_gen[14].d2.D ;
	reg \mchip.aa.i0.dff_gen[14].d2.Q ;
	wire \mchip.aa.i0.dff_gen[14].d2.clk ;
	wire \mchip.aa.i0.dff_gen[15].d2.D ;
	reg \mchip.aa.i0.dff_gen[15].d2.Q ;
	wire \mchip.aa.i0.dff_gen[15].d2.clk ;
	wire \mchip.aa.i0.dff_gen[16].d2.D ;
	wire \mchip.aa.i0.dff_gen[16].d2.Q ;
	wire \mchip.aa.i0.dff_gen[16].d2.clk ;
	wire \mchip.aa.i0.dff_gen[17].d2.D ;
	wire \mchip.aa.i0.dff_gen[17].d2.Q ;
	wire \mchip.aa.i0.dff_gen[17].d2.clk ;
	wire \mchip.aa.i0.dff_gen[18].d2.D ;
	wire \mchip.aa.i0.dff_gen[18].d2.Q ;
	wire \mchip.aa.i0.dff_gen[18].d2.clk ;
	wire \mchip.aa.i0.dff_gen[19].d2.D ;
	wire \mchip.aa.i0.dff_gen[19].d2.Q ;
	wire \mchip.aa.i0.dff_gen[19].d2.clk ;
	wire \mchip.aa.i0.dff_gen[1].d2.D ;
	reg \mchip.aa.i0.dff_gen[1].d2.Q ;
	wire \mchip.aa.i0.dff_gen[1].d2.clk ;
	wire \mchip.aa.i0.dff_gen[2].d2.D ;
	reg \mchip.aa.i0.dff_gen[2].d2.Q ;
	wire \mchip.aa.i0.dff_gen[2].d2.clk ;
	wire \mchip.aa.i0.dff_gen[3].d2.D ;
	reg \mchip.aa.i0.dff_gen[3].d2.Q ;
	wire \mchip.aa.i0.dff_gen[3].d2.clk ;
	wire \mchip.aa.i0.dff_gen[4].d2.D ;
	reg \mchip.aa.i0.dff_gen[4].d2.Q ;
	wire \mchip.aa.i0.dff_gen[4].d2.clk ;
	wire \mchip.aa.i0.dff_gen[5].d2.D ;
	reg \mchip.aa.i0.dff_gen[5].d2.Q ;
	wire \mchip.aa.i0.dff_gen[5].d2.clk ;
	wire \mchip.aa.i0.dff_gen[6].d2.D ;
	reg \mchip.aa.i0.dff_gen[6].d2.Q ;
	wire \mchip.aa.i0.dff_gen[6].d2.clk ;
	wire \mchip.aa.i0.dff_gen[7].d2.D ;
	reg \mchip.aa.i0.dff_gen[7].d2.Q ;
	wire \mchip.aa.i0.dff_gen[7].d2.clk ;
	wire \mchip.aa.i0.dff_gen[8].d2.D ;
	reg \mchip.aa.i0.dff_gen[8].d2.Q ;
	wire \mchip.aa.i0.dff_gen[8].d2.clk ;
	wire \mchip.aa.i0.dff_gen[9].d2.D ;
	reg \mchip.aa.i0.dff_gen[9].d2.Q ;
	wire \mchip.aa.i0.dff_gen[9].d2.clk ;
	wire [19:0] \mchip.aa.i0.in ;
	wire [19:0] \mchip.aa.i0.out ;
	wire [19:0] \mchip.aa.i0.temp_out ;
	wire [15:0] \mchip.aa.mult_res_in ;
	wire [19:0] \mchip.aa.mult_res_out ;
	wire [19:0] \mchip.aa.result ;
	wire \mchip.aa.result_carry_out ;
	wire [19:0] \mchip.aa.temp_mult_res_in ;
	wire [19:0] \mchip.aa.temp_result ;
	wire \mchip.add ;
	wire \mchip.clock ;
	wire \mchip.control.Begin_mul ;
	wire \mchip.control.End_mul ;
	wire \mchip.control.Finish ;
	wire \mchip.control.Load_op ;
	wire \mchip.control.START ;
	reg \mchip.control._do_next ;
	wire \mchip.control.add ;
	wire \mchip.control.clk ;
	wire \mchip.control.do_next ;
	reg [6:0] \mchip.control.state ;
	reg [3:0] \mchip.control.temp_count ;
	wire \mchip.do_next ;
	wire [11:0] \mchip.io_in ;
	wire [11:0] \mchip.io_out ;
	wire \mchip.mac_carry_out ;
	wire [19:0] \mchip.mac_res ;
	wire \mchip.mult.Begin_mul ;
	wire \mchip.mult.End_mul ;
	wire \mchip.mult.LSB ;
	wire \mchip.mult.Load_mul ;
	wire [7:0] \mchip.mult.a_in ;
	wire [7:0] \mchip.mult.a_out ;
	wire [7:0] \mchip.mult.b_in ;
	wire [7:0] \mchip.mult.b_out ;
	wire \mchip.mult.clk ;
	wire \mchip.mult.do_add ;
	wire \mchip.mult.do_shift ;
	wire \mchip.mult.i0.Begin_mul ;
	wire \mchip.mult.i0.End_mul ;
	wire \mchip.mult.i0.LSB ;
	wire \mchip.mult.i0.Load_mul ;
	wire \mchip.mult.i0.clk ;
	wire \mchip.mult.i0.do_add ;
	wire \mchip.mult.i0.do_shift ;
	reg [4:0] \mchip.mult.i0.state ;
	reg [2:0] \mchip.mult.i0.temp_count ;
	wire \mchip.mult.i1.Load_mul ;
	wire [7:0] \mchip.mult.i1.a_in ;
	wire [7:0] \mchip.mult.i1.a_out ;
	wire \mchip.mult.i1.r1.Load_op ;
	wire \mchip.mult.i1.r1.dff_gen[0].d1.D ;
	reg \mchip.mult.i1.r1.dff_gen[0].d1.Q ;
	wire \mchip.mult.i1.r1.dff_gen[0].d1.clk ;
	wire \mchip.mult.i1.r1.dff_gen[1].d1.D ;
	reg \mchip.mult.i1.r1.dff_gen[1].d1.Q ;
	wire \mchip.mult.i1.r1.dff_gen[1].d1.clk ;
	wire \mchip.mult.i1.r1.dff_gen[2].d1.D ;
	reg \mchip.mult.i1.r1.dff_gen[2].d1.Q ;
	wire \mchip.mult.i1.r1.dff_gen[2].d1.clk ;
	wire \mchip.mult.i1.r1.dff_gen[3].d1.D ;
	reg \mchip.mult.i1.r1.dff_gen[3].d1.Q ;
	wire \mchip.mult.i1.r1.dff_gen[3].d1.clk ;
	wire \mchip.mult.i1.r1.dff_gen[4].d1.D ;
	reg \mchip.mult.i1.r1.dff_gen[4].d1.Q ;
	wire \mchip.mult.i1.r1.dff_gen[4].d1.clk ;
	wire \mchip.mult.i1.r1.dff_gen[5].d1.D ;
	reg \mchip.mult.i1.r1.dff_gen[5].d1.Q ;
	wire \mchip.mult.i1.r1.dff_gen[5].d1.clk ;
	wire \mchip.mult.i1.r1.dff_gen[6].d1.D ;
	reg \mchip.mult.i1.r1.dff_gen[6].d1.Q ;
	wire \mchip.mult.i1.r1.dff_gen[6].d1.clk ;
	wire \mchip.mult.i1.r1.dff_gen[7].d1.D ;
	reg \mchip.mult.i1.r1.dff_gen[7].d1.Q ;
	wire \mchip.mult.i1.r1.dff_gen[7].d1.clk ;
	wire [7:0] \mchip.mult.i1.r1.in ;
	wire [7:0] \mchip.mult.i1.r1.out ;
	wire [7:0] \mchip.mult.i1.r1.temp_out ;
	wire [3:0] \mchip.mult.i2.S0.S0.a ;
	wire [3:0] \mchip.mult.i2.S0.S0.b ;
	wire \mchip.mult.i2.S0.S0.carry_in ;
	wire \mchip.mult.i2.S0.S0.fa0.a ;
	wire \mchip.mult.i2.S0.S0.fa0.b ;
	wire \mchip.mult.i2.S0.S0.fa0.carry_in ;
	wire \mchip.mult.i2.S0.S0.fa0.w3 ;
	wire \mchip.mult.i2.S0.S0.fa1.a ;
	wire \mchip.mult.i2.S0.S0.fa1.b ;
	wire \mchip.mult.i2.S0.S0.fa2.a ;
	wire \mchip.mult.i2.S0.S0.fa2.b ;
	wire \mchip.mult.i2.S0.S0.fa3.a ;
	wire \mchip.mult.i2.S0.S0.fa3.b ;
	wire [3:0] \mchip.mult.i2.S0.S1.a ;
	wire [3:0] \mchip.mult.i2.S0.S1.b ;
	wire \mchip.mult.i2.S0.S1.carry_in ;
	wire \mchip.mult.i2.S0.S1.fa0.a ;
	wire \mchip.mult.i2.S0.S1.fa0.b ;
	wire \mchip.mult.i2.S0.S1.fa0.carry_in ;
	wire \mchip.mult.i2.S0.S1.fa1.a ;
	wire \mchip.mult.i2.S0.S1.fa1.b ;
	wire \mchip.mult.i2.S0.S1.fa2.a ;
	wire \mchip.mult.i2.S0.S1.fa2.b ;
	wire \mchip.mult.i2.S0.S1.fa3.a ;
	wire \mchip.mult.i2.S0.S1.fa3.b ;
	wire [3:0] \mchip.mult.i2.S0.a ;
	wire [3:0] \mchip.mult.i2.S0.b ;
	wire \mchip.mult.i2.S0.carry_in ;
	wire [3:0] \mchip.mult.i2.S1.S0.a ;
	wire [3:0] \mchip.mult.i2.S1.S0.b ;
	wire \mchip.mult.i2.S1.S0.carry_in ;
	wire \mchip.mult.i2.S1.S0.fa0.a ;
	wire \mchip.mult.i2.S1.S0.fa0.b ;
	wire \mchip.mult.i2.S1.S0.fa0.carry_in ;
	wire \mchip.mult.i2.S1.S0.fa0.w3 ;
	wire \mchip.mult.i2.S1.S0.fa1.a ;
	wire \mchip.mult.i2.S1.S0.fa1.b ;
	wire \mchip.mult.i2.S1.S0.fa2.a ;
	wire \mchip.mult.i2.S1.S0.fa2.b ;
	wire \mchip.mult.i2.S1.S0.fa3.a ;
	wire \mchip.mult.i2.S1.S0.fa3.b ;
	wire [3:0] \mchip.mult.i2.S1.S0.sum ;
	wire [3:0] \mchip.mult.i2.S1.S1.a ;
	wire [3:0] \mchip.mult.i2.S1.S1.b ;
	wire \mchip.mult.i2.S1.S1.carry_in ;
	wire \mchip.mult.i2.S1.S1.fa0.a ;
	wire \mchip.mult.i2.S1.S1.fa0.b ;
	wire \mchip.mult.i2.S1.S1.fa0.carry_in ;
	wire \mchip.mult.i2.S1.S1.fa1.a ;
	wire \mchip.mult.i2.S1.S1.fa1.b ;
	wire \mchip.mult.i2.S1.S1.fa2.a ;
	wire \mchip.mult.i2.S1.S1.fa2.b ;
	wire \mchip.mult.i2.S1.S1.fa3.a ;
	wire \mchip.mult.i2.S1.S1.fa3.b ;
	wire [3:0] \mchip.mult.i2.S1.S1.sum ;
	wire [3:0] \mchip.mult.i2.S1.SUM0 ;
	wire [3:0] \mchip.mult.i2.S1.SUM1 ;
	wire [3:0] \mchip.mult.i2.S1.a ;
	wire [3:0] \mchip.mult.i2.S1.b ;
	wire [7:0] \mchip.mult.i2.a ;
	wire [7:0] \mchip.mult.i2.b ;
	wire \mchip.mult.i2.carry_in ;
	wire \mchip.mult.i3.LSB ;
	wire \mchip.mult.i3.Load_mul ;
	wire [7:0] \mchip.mult.i3.b_in ;
	wire [7:0] \mchip.mult.i3.b_out ;
	wire \mchip.mult.i3.clk ;
	wire \mchip.mult.i3.do_add ;
	wire \mchip.mult.i3.do_shift ;
	wire [15:0] \mchip.mult.i3.mult_out ;
	reg \mchip.mult.i3.temp_Add ;
	wire [16:0] \mchip.mult.i3.temp_register ;
	wire [15:0] \mchip.mult.mult_out ;
	wire [15:0] \mchip.mult_res ;
	reg [7:0] \mchip.op_a_in ;
	wire [7:0] \mchip.op_a_out ;
	reg [7:0] \mchip.op_b_in ;
	wire [7:0] \mchip.op_b_out ;
	wire \mchip.opa.Load_op ;
	wire \mchip.opa.dff_gen[0].d1.D ;
	reg \mchip.opa.dff_gen[0].d1.Q ;
	wire \mchip.opa.dff_gen[0].d1.clk ;
	wire \mchip.opa.dff_gen[1].d1.D ;
	reg \mchip.opa.dff_gen[1].d1.Q ;
	wire \mchip.opa.dff_gen[1].d1.clk ;
	wire \mchip.opa.dff_gen[2].d1.D ;
	reg \mchip.opa.dff_gen[2].d1.Q ;
	wire \mchip.opa.dff_gen[2].d1.clk ;
	wire \mchip.opa.dff_gen[3].d1.D ;
	reg \mchip.opa.dff_gen[3].d1.Q ;
	wire \mchip.opa.dff_gen[3].d1.clk ;
	wire \mchip.opa.dff_gen[4].d1.D ;
	reg \mchip.opa.dff_gen[4].d1.Q ;
	wire \mchip.opa.dff_gen[4].d1.clk ;
	wire \mchip.opa.dff_gen[5].d1.D ;
	reg \mchip.opa.dff_gen[5].d1.Q ;
	wire \mchip.opa.dff_gen[5].d1.clk ;
	wire \mchip.opa.dff_gen[6].d1.D ;
	reg \mchip.opa.dff_gen[6].d1.Q ;
	wire \mchip.opa.dff_gen[6].d1.clk ;
	wire \mchip.opa.dff_gen[7].d1.D ;
	reg \mchip.opa.dff_gen[7].d1.Q ;
	wire \mchip.opa.dff_gen[7].d1.clk ;
	wire [7:0] \mchip.opa.in ;
	wire [7:0] \mchip.opa.out ;
	wire [7:0] \mchip.opa.temp_out ;
	wire \mchip.opb.Load_op ;
	wire \mchip.opb.dff_gen[0].d1.D ;
	reg \mchip.opb.dff_gen[0].d1.Q ;
	wire \mchip.opb.dff_gen[0].d1.clk ;
	wire \mchip.opb.dff_gen[1].d1.D ;
	reg \mchip.opb.dff_gen[1].d1.Q ;
	wire \mchip.opb.dff_gen[1].d1.clk ;
	wire \mchip.opb.dff_gen[2].d1.D ;
	reg \mchip.opb.dff_gen[2].d1.Q ;
	wire \mchip.opb.dff_gen[2].d1.clk ;
	wire \mchip.opb.dff_gen[3].d1.D ;
	reg \mchip.opb.dff_gen[3].d1.Q ;
	wire \mchip.opb.dff_gen[3].d1.clk ;
	wire \mchip.opb.dff_gen[4].d1.D ;
	reg \mchip.opb.dff_gen[4].d1.Q ;
	wire \mchip.opb.dff_gen[4].d1.clk ;
	wire \mchip.opb.dff_gen[5].d1.D ;
	reg \mchip.opb.dff_gen[5].d1.Q ;
	wire \mchip.opb.dff_gen[5].d1.clk ;
	wire \mchip.opb.dff_gen[6].d1.D ;
	reg \mchip.opb.dff_gen[6].d1.Q ;
	wire \mchip.opb.dff_gen[6].d1.clk ;
	wire \mchip.opb.dff_gen[7].d1.D ;
	reg \mchip.opb.dff_gen[7].d1.Q ;
	wire \mchip.opb.dff_gen[7].d1.clk ;
	wire [7:0] \mchip.opb.in ;
	wire [7:0] \mchip.opb.out ;
	wire [7:0] \mchip.opb.temp_out ;
	wire \mchip.reset ;
	reg \mchip.shiftin ;
	reg [19:0] \mchip.shiftout ;
	assign _012_ = io_in[13] | \mchip.control.state [4];
	assign _062_ = \mchip.mult.i0.temp_count [0] & \mchip.mult.i0.temp_count [1];
	assign _063_ = _062_ & \mchip.mult.i0.temp_count [2];
	assign _064_ = _063_ | _012_;
	assign _065_ = \mchip.mult.i0.state [1] & ~_064_;
	assign _066_ = \mchip.mult.i0.state [3] & ~_012_;
	assign _011_ = _066_ | _065_;
	assign _048_ = \mchip.control.state [0] & ~\mchip._Finish ;
	assign _047_ = io_in[8] & ~\mchip.shiftin ;
	assign _014_ = _047_ | _048_;
	assign _067_ = ~(\mchip.control.temp_count [1] | \mchip.control.temp_count [0]);
	assign _068_ = \mchip.control.temp_count [3] | \mchip.control.temp_count [2];
	assign _069_ = _067_ & ~_068_;
	assign _070_ = (\mchip.control.state [5] ? _069_ : \mchip.control.state [3]);
	assign _071_ = io_in[7] & ~\mchip.control._do_next ;
	assign _072_ = \mchip.control.state [3] & ~_071_;
	assign _015_ = _070_ & ~_072_;
	assign _073_ = \mchip.mult.i0.state [4] & ~_012_;
	assign _074_ = _012_ | \mchip.mult.i3.temp_register [0];
	assign _075_ = \mchip.mult.i0.state [2] & ~_074_;
	assign _010_ = _075_ | _073_;
	assign _076_ = _012_ | ~_063_;
	assign _077_ = \mchip.mult.i0.state [1] & ~_076_;
	assign _078_ = _012_ | \mchip.control.state [6];
	assign _079_ = \mchip.mult.i0.state [0] & ~_078_;
	assign _080_ = _079_ | _077_;
	assign _009_ = _080_ | _012_;
	assign _081_ = io_in[11] | io_in[13];
	assign _082_ = \mchip.control.state [0] & ~_081_;
	assign _083_ = io_in[13] | ~_069_;
	assign _084_ = \mchip.control.state [5] & ~_083_;
	assign _085_ = _084_ | io_in[13];
	assign _005_ = _085_ | _082_;
	assign _086_ = \mchip.mult.i0.state [0] | io_in[13];
	assign _087_ = \mchip.control.state [1] & ~_086_;
	assign _088_ = \mchip.control.state [6] & ~io_in[13];
	assign _006_ = _088_ | _087_;
	assign _016_ = _012_ | \mchip.mult.i0.state [3];
	assign _013_ = \mchip.mult.i0.state [1] | \mchip.mult.i0.state [3];
	assign _089_ = _069_ | io_in[13];
	assign _090_ = \mchip.control.state [5] & ~_089_;
	assign _091_ = _071_ | io_in[13];
	assign _092_ = \mchip.control.state [3] & ~_091_;
	assign _008_ = _092_ | _090_;
	assign _093_ = io_in[13] | ~_071_;
	assign _094_ = \mchip.control.state [3] & ~_093_;
	assign _095_ = \mchip.control.state [4] & ~io_in[13];
	assign _007_ = _095_ | _094_;
	assign _096_ = \mchip.control.temp_count [1] ^ \mchip.control.temp_count [0];
	assign _050_ = \mchip.control.state [3] & ~_096_;
	assign _097_ = ~(_067_ ^ \mchip.control.temp_count [2]);
	assign _051_ = \mchip.control.state [3] & ~_097_;
	assign _098_ = _067_ & ~\mchip.control.temp_count [2];
	assign _099_ = ~(_098_ ^ \mchip.control.temp_count [3]);
	assign _052_ = ~(_099_ & \mchip.control.state [3]);
	assign _028_ = (_048_ ? \mchip.aa.accmulate.dff_gen[0].d2.Q  : \mchip.shiftout [1]);
	assign _038_ = (_048_ ? \mchip.aa.accmulate.dff_gen[1].d2.Q  : \mchip.shiftout [2]);
	assign _039_ = (_048_ ? \mchip.aa.accmulate.dff_gen[2].d2.Q  : \mchip.shiftout [3]);
	assign _040_ = (_048_ ? \mchip.aa.accmulate.dff_gen[3].d2.Q  : \mchip.shiftout [4]);
	assign _041_ = (_048_ ? \mchip.aa.accmulate.dff_gen[4].d2.Q  : \mchip.shiftout [5]);
	assign _042_ = (_048_ ? \mchip.aa.accmulate.dff_gen[5].d2.Q  : \mchip.shiftout [6]);
	assign _043_ = (_048_ ? \mchip.aa.accmulate.dff_gen[6].d2.Q  : \mchip.shiftout [7]);
	assign _044_ = (_048_ ? \mchip.aa.accmulate.dff_gen[7].d2.Q  : \mchip.shiftout [8]);
	assign _045_ = (_048_ ? \mchip.aa.accmulate.dff_gen[8].d2.Q  : \mchip.shiftout [9]);
	assign _046_ = (_048_ ? \mchip.aa.accmulate.dff_gen[9].d2.Q  : \mchip.shiftout [10]);
	assign _029_ = (_048_ ? \mchip.aa.accmulate.dff_gen[10].d2.Q  : \mchip.shiftout [11]);
	assign _030_ = (_048_ ? \mchip.aa.accmulate.dff_gen[11].d2.Q  : \mchip.shiftout [12]);
	assign _031_ = (_048_ ? \mchip.aa.accmulate.dff_gen[12].d2.Q  : \mchip.shiftout [13]);
	assign _032_ = (_048_ ? \mchip.aa.accmulate.dff_gen[13].d2.Q  : \mchip.shiftout [14]);
	assign _033_ = (_048_ ? \mchip.aa.accmulate.dff_gen[14].d2.Q  : \mchip.shiftout [15]);
	assign _034_ = (_048_ ? \mchip.aa.accmulate.dff_gen[15].d2.Q  : \mchip.shiftout [16]);
	assign _035_ = (_048_ ? \mchip.aa.accmulate.dff_gen[16].d2.Q  : \mchip.shiftout [17]);
	assign _036_ = (_048_ ? \mchip.aa.accmulate.dff_gen[17].d2.Q  : \mchip.shiftout [18]);
	assign _037_ = (_048_ ? \mchip.aa.accmulate.dff_gen[18].d2.Q  : \mchip.shiftout [19]);
	assign _100_ = \mchip.aa.i0.dff_gen[11].d2.Q  & \mchip.aa.accmulate.dff_gen[11].d2.Q ;
	assign _101_ = \mchip.aa.i0.dff_gen[10].d2.Q  & \mchip.aa.accmulate.dff_gen[10].d2.Q ;
	assign _102_ = \mchip.aa.i0.dff_gen[10].d2.Q  ^ \mchip.aa.accmulate.dff_gen[10].d2.Q ;
	assign _103_ = ~(\mchip.aa.i0.dff_gen[9].d2.Q  & \mchip.aa.accmulate.dff_gen[9].d2.Q );
	assign _104_ = \mchip.aa.i0.dff_gen[9].d2.Q  ^ \mchip.aa.accmulate.dff_gen[9].d2.Q ;
	assign _105_ = ~(\mchip.aa.i0.dff_gen[8].d2.Q  | \mchip.aa.accmulate.dff_gen[8].d2.Q );
	assign _106_ = _104_ & ~_105_;
	assign _107_ = _103_ & ~_106_;
	assign _108_ = _102_ & ~_107_;
	assign _109_ = _108_ | _101_;
	assign _110_ = \mchip.aa.i0.dff_gen[11].d2.Q  ^ \mchip.aa.accmulate.dff_gen[11].d2.Q ;
	assign _111_ = _110_ & _109_;
	assign _112_ = ~(_111_ | _100_);
	assign _113_ = \mchip.aa.i0.dff_gen[6].d2.Q  & \mchip.aa.accmulate.dff_gen[6].d2.Q ;
	assign _114_ = \mchip.aa.i0.dff_gen[6].d2.Q  ^ \mchip.aa.accmulate.dff_gen[6].d2.Q ;
	assign _115_ = ~(\mchip.aa.i0.dff_gen[5].d2.Q  & \mchip.aa.accmulate.dff_gen[5].d2.Q );
	assign _116_ = \mchip.aa.i0.dff_gen[5].d2.Q  ^ \mchip.aa.accmulate.dff_gen[5].d2.Q ;
	assign _117_ = ~(\mchip.aa.i0.dff_gen[4].d2.Q  | \mchip.aa.accmulate.dff_gen[4].d2.Q );
	assign _118_ = _116_ & ~_117_;
	assign _119_ = _115_ & ~_118_;
	assign _120_ = _114_ & ~_119_;
	assign _121_ = _120_ | _113_;
	assign _122_ = \mchip.aa.i0.dff_gen[7].d2.Q  ^ \mchip.aa.accmulate.dff_gen[7].d2.Q ;
	assign _123_ = ~(_122_ & _121_);
	assign _124_ = \mchip.aa.i0.dff_gen[7].d2.Q  & \mchip.aa.accmulate.dff_gen[7].d2.Q ;
	assign _125_ = _123_ & ~_124_;
	assign _126_ = \mchip.aa.i0.dff_gen[3].d2.Q  ^ \mchip.aa.accmulate.dff_gen[3].d2.Q ;
	assign _127_ = ~(\mchip.aa.i0.dff_gen[2].d2.Q  & \mchip.aa.accmulate.dff_gen[2].d2.Q );
	assign _128_ = \mchip.aa.i0.dff_gen[2].d2.Q  ^ \mchip.aa.accmulate.dff_gen[2].d2.Q ;
	assign _129_ = ~(\mchip.aa.i0.dff_gen[1].d2.Q  & \mchip.aa.accmulate.dff_gen[1].d2.Q );
	assign _130_ = \mchip.aa.i0.dff_gen[1].d2.Q  ^ \mchip.aa.accmulate.dff_gen[1].d2.Q ;
	assign _131_ = ~(\mchip.aa.i0.dff_gen[0].d2.Q  & \mchip.aa.accmulate.dff_gen[0].d2.Q );
	assign _132_ = _130_ & ~_131_;
	assign _133_ = _129_ & ~_132_;
	assign _134_ = _128_ & ~_133_;
	assign _135_ = _127_ & ~_134_;
	assign _136_ = _126_ & ~_135_;
	assign _137_ = \mchip.aa.i0.dff_gen[3].d2.Q  & \mchip.aa.accmulate.dff_gen[3].d2.Q ;
	assign _138_ = _137_ | _136_;
	assign _139_ = _138_ & ~_125_;
	assign _140_ = ~(\mchip.aa.i0.dff_gen[4].d2.Q  & \mchip.aa.accmulate.dff_gen[4].d2.Q );
	assign _141_ = _116_ & ~_140_;
	assign _142_ = _115_ & ~_141_;
	assign _143_ = _114_ & ~_142_;
	assign _144_ = ~(_143_ | _113_);
	assign _145_ = _122_ & ~_144_;
	assign _146_ = _145_ | _124_;
	assign _147_ = _146_ | _139_;
	assign _148_ = _112_ | ~_147_;
	assign _149_ = ~(\mchip.aa.i0.dff_gen[8].d2.Q  & \mchip.aa.accmulate.dff_gen[8].d2.Q );
	assign _150_ = _104_ & ~_149_;
	assign _151_ = _103_ & ~_150_;
	assign _152_ = _102_ & ~_151_;
	assign _153_ = ~(_152_ | _101_);
	assign _154_ = _110_ & ~_153_;
	assign _155_ = _154_ | _100_;
	assign _156_ = _155_ | ~_148_;
	assign _157_ = \mchip.aa.i0.dff_gen[12].d2.Q  | \mchip.aa.accmulate.dff_gen[12].d2.Q ;
	assign _158_ = \mchip.aa.i0.dff_gen[12].d2.Q  & \mchip.aa.accmulate.dff_gen[12].d2.Q ;
	assign _159_ = _157_ & ~_158_;
	assign \mchip.aa.accmulate.dff_gen[12].d2.D  = _159_ ^ _156_;
	assign _160_ = _149_ & ~_105_;
	assign \mchip.aa.accmulate.dff_gen[8].d2.D  = _160_ ^ _147_;
	assign _161_ = _140_ & ~_117_;
	assign \mchip.aa.accmulate.dff_gen[4].d2.D  = _161_ ^ _138_;
	assign _017_ = ~(_063_ | \mchip.mult.i0.temp_count [0]);
	assign _018_ = \mchip.mult.i0.temp_count [0] ^ \mchip.mult.i0.temp_count [1];
	assign _019_ = _062_ ^ \mchip.mult.i0.temp_count [2];
	assign _162_ = ~\mchip.mult.i0.state [1];
	assign _053_ = (\mchip.mult.i3.temp_Add  ? _162_ : \mchip.mult.i0.state [4]);
	assign _054_ = (\mchip.mult.i0.state [3] ? \mchip.opb.dff_gen[0].d1.Q  : \mchip.mult.i3.temp_register [1]);
	assign _055_ = (\mchip.mult.i0.state [3] ? \mchip.opb.dff_gen[1].d1.Q  : \mchip.mult.i3.temp_register [2]);
	assign _056_ = (\mchip.mult.i0.state [3] ? \mchip.opb.dff_gen[2].d1.Q  : \mchip.mult.i3.temp_register [3]);
	assign _057_ = (\mchip.mult.i0.state [3] ? \mchip.opb.dff_gen[3].d1.Q  : \mchip.mult.i3.temp_register [4]);
	assign _058_ = (\mchip.mult.i0.state [3] ? \mchip.opb.dff_gen[4].d1.Q  : \mchip.mult.i3.temp_register [5]);
	assign _059_ = (\mchip.mult.i0.state [3] ? \mchip.opb.dff_gen[5].d1.Q  : \mchip.mult.i3.temp_register [6]);
	assign _060_ = (\mchip.mult.i0.state [3] ? \mchip.opb.dff_gen[6].d1.Q  : \mchip.mult.i3.temp_register [7]);
	assign _163_ = \mchip.mult.i3.temp_register [8] ^ \mchip.mult.i1.r1.dff_gen[0].d1.Q ;
	assign _164_ = (\mchip.mult.i3.temp_Add  ? _163_ : \mchip.mult.i3.temp_register [8]);
	assign _061_ = (\mchip.mult.i0.state [3] ? \mchip.opb.dff_gen[7].d1.Q  : _164_);
	assign _165_ = \mchip.mult.i3.temp_register [8] & \mchip.mult.i1.r1.dff_gen[0].d1.Q ;
	assign _166_ = ~(\mchip.mult.i3.temp_register [9] ^ \mchip.mult.i1.r1.dff_gen[1].d1.Q );
	assign _167_ = ~(_166_ ^ _165_);
	assign _020_ = (\mchip.mult.i3.temp_Add  ? _167_ : \mchip.mult.i3.temp_register [9]);
	assign _168_ = \mchip.mult.i3.temp_register [9] & \mchip.mult.i1.r1.dff_gen[1].d1.Q ;
	assign _169_ = _165_ & ~_166_;
	assign _170_ = _169_ | _168_;
	assign _171_ = \mchip.mult.i3.temp_register [10] ^ \mchip.mult.i1.r1.dff_gen[2].d1.Q ;
	assign _172_ = _171_ ^ _170_;
	assign _021_ = (\mchip.mult.i3.temp_Add  ? _172_ : \mchip.mult.i3.temp_register [10]);
	assign _173_ = \mchip.mult.i3.temp_register [10] & \mchip.mult.i1.r1.dff_gen[2].d1.Q ;
	assign _174_ = _171_ & _170_;
	assign _175_ = _174_ | _173_;
	assign _176_ = \mchip.mult.i3.temp_register [11] ^ \mchip.mult.i1.r1.dff_gen[3].d1.Q ;
	assign _177_ = _176_ ^ _175_;
	assign _022_ = (\mchip.mult.i3.temp_Add  ? _177_ : \mchip.mult.i3.temp_register [11]);
	assign _178_ = \mchip.mult.i3.temp_register [11] & \mchip.mult.i1.r1.dff_gen[3].d1.Q ;
	assign _179_ = _176_ & _175_;
	assign _180_ = _179_ | _178_;
	assign _181_ = \mchip.mult.i3.temp_register [12] | \mchip.mult.i1.r1.dff_gen[4].d1.Q ;
	assign _182_ = \mchip.mult.i3.temp_register [12] & \mchip.mult.i1.r1.dff_gen[4].d1.Q ;
	assign _183_ = _181_ & ~_182_;
	assign _184_ = _183_ ^ _180_;
	assign _023_ = (\mchip.mult.i3.temp_Add  ? _184_ : \mchip.mult.i3.temp_register [12]);
	assign _185_ = (_180_ ? _181_ : _182_);
	assign _186_ = ~(\mchip.mult.i3.temp_register [13] ^ \mchip.mult.i1.r1.dff_gen[5].d1.Q );
	assign _187_ = ~(_186_ ^ _185_);
	assign _024_ = (\mchip.mult.i3.temp_Add  ? _187_ : \mchip.mult.i3.temp_register [13]);
	assign _188_ = \mchip.mult.i3.temp_register [13] & \mchip.mult.i1.r1.dff_gen[5].d1.Q ;
	assign _189_ = _181_ & ~_186_;
	assign _190_ = _189_ | _188_;
	assign _191_ = _182_ & ~_186_;
	assign _192_ = _191_ | _188_;
	assign _193_ = (_180_ ? _190_ : _192_);
	assign _194_ = \mchip.mult.i3.temp_register [14] ^ \mchip.mult.i1.r1.dff_gen[6].d1.Q ;
	assign _195_ = _194_ ^ _193_;
	assign _025_ = (\mchip.mult.i3.temp_Add  ? _195_ : \mchip.mult.i3.temp_register [14]);
	assign _196_ = \mchip.mult.i3.temp_register [14] & \mchip.mult.i1.r1.dff_gen[6].d1.Q ;
	assign _197_ = ~_194_;
	assign _198_ = _190_ & ~_197_;
	assign _199_ = _198_ | _196_;
	assign _200_ = _192_ & ~_197_;
	assign _201_ = _200_ | _196_;
	assign _202_ = (_180_ ? _199_ : _201_);
	assign _203_ = \mchip.mult.i3.temp_register [15] ^ \mchip.mult.i1.r1.dff_gen[7].d1.Q ;
	assign _204_ = _203_ ^ _202_;
	assign _026_ = (\mchip.mult.i3.temp_Add  ? _204_ : \mchip.mult.i3.temp_register [15]);
	assign _205_ = \mchip.mult.i3.temp_register [15] & \mchip.mult.i1.r1.dff_gen[7].d1.Q ;
	assign _206_ = ~_203_;
	assign _207_ = _199_ & ~_206_;
	assign _208_ = _207_ | _205_;
	assign _209_ = ~(_208_ & _180_);
	assign _210_ = _201_ & ~_206_;
	assign _211_ = _210_ | _205_;
	assign _212_ = _209_ & ~_211_;
	assign _027_ = \mchip.mult.i3.temp_Add  & ~_212_;
	assign _049_ = ~(\mchip.control.state [3] & \mchip.control.temp_count [0]);
	assign \mchip.aa.adder.S4.S1.fa0.sum  = ~\mchip.aa.accmulate.dff_gen[16].d2.Q ;
	assign _213_ = _012_ | ~\mchip.mult.i3.temp_register [0];
	assign _004_ = \mchip.mult.i0.state [2] & ~_213_;
	assign _214_ = _012_ | ~\mchip.control.state [6];
	assign _003_ = \mchip.mult.i0.state [0] & ~_214_;
	assign \mchip.aa.accmulate.dff_gen[0].d2.D  = \mchip.aa.i0.dff_gen[0].d2.Q  ^ \mchip.aa.accmulate.dff_gen[0].d2.Q ;
	assign _215_ = \mchip.aa.i0.dff_gen[15].d2.Q  & \mchip.aa.accmulate.dff_gen[15].d2.Q ;
	assign _216_ = \mchip.aa.i0.dff_gen[14].d2.Q  & \mchip.aa.accmulate.dff_gen[14].d2.Q ;
	assign _217_ = \mchip.aa.i0.dff_gen[14].d2.Q  ^ \mchip.aa.accmulate.dff_gen[14].d2.Q ;
	assign _218_ = \mchip.aa.i0.dff_gen[13].d2.Q  & \mchip.aa.accmulate.dff_gen[13].d2.Q ;
	assign _219_ = ~_218_;
	assign _220_ = ~(\mchip.aa.i0.dff_gen[13].d2.Q  ^ \mchip.aa.accmulate.dff_gen[13].d2.Q );
	assign _221_ = _158_ & ~_220_;
	assign _222_ = _219_ & ~_221_;
	assign _223_ = _217_ & ~_222_;
	assign _224_ = _223_ | _216_;
	assign _225_ = \mchip.aa.i0.dff_gen[15].d2.Q  ^ \mchip.aa.accmulate.dff_gen[15].d2.Q ;
	assign _226_ = _225_ & _224_;
	assign _227_ = _226_ | _215_;
	assign _228_ = _157_ & ~_220_;
	assign _229_ = _219_ & ~_228_;
	assign _230_ = _217_ & ~_229_;
	assign _231_ = ~(_230_ | _216_);
	assign _232_ = _231_ | ~_225_;
	assign _233_ = _232_ & ~_215_;
	assign _234_ = _156_ & ~_233_;
	assign \mchip.aa.adder.S4.carry_in  = _234_ | _227_;
	assign _235_ = \mchip.aa.accmulate.dff_gen[17].d2.Q  & \mchip.aa.accmulate.dff_gen[16].d2.Q ;
	assign _236_ = _235_ & \mchip.aa.accmulate.dff_gen[18].d2.Q ;
	assign _237_ = ~(_236_ & \mchip.aa.accmulate.dff_gen[19].d2.Q );
	assign \mchip.aa.adder.S4.carry_out  = \mchip.aa.adder.S4.carry_in  & ~_237_;
	assign _002_ = \mchip.control.state [2] & ~io_in[13];
	assign _238_ = io_in[13] | ~\mchip.mult.i0.state [0];
	assign _001_ = \mchip.control.state [1] & ~_238_;
	assign \mchip.aa.adder.S4.S1.fa3.sum  = _236_ ^ \mchip.aa.accmulate.dff_gen[19].d2.Q ;
	assign \mchip.aa.adder.S4.S1.fa2.sum  = _235_ ^ \mchip.aa.accmulate.dff_gen[18].d2.Q ;
	assign \mchip.aa.adder.S4.S1.fa1.sum  = \mchip.aa.accmulate.dff_gen[17].d2.Q  ^ \mchip.aa.accmulate.dff_gen[16].d2.Q ;
	assign _239_ = _148_ & ~_155_;
	assign _240_ = ~_231_;
	assign _241_ = (_239_ ? _224_ : _240_);
	assign \mchip.aa.accmulate.dff_gen[15].d2.D  = _241_ ^ _225_;
	assign _242_ = (_239_ ? _222_ : _229_);
	assign \mchip.aa.accmulate.dff_gen[14].d2.D  = ~(_242_ ^ _217_);
	assign _243_ = (_156_ ? _157_ : _158_);
	assign \mchip.aa.accmulate.dff_gen[13].d2.D  = ~(_243_ ^ _220_);
	assign _244_ = ~_153_;
	assign _245_ = (_147_ ? _109_ : _244_);
	assign \mchip.aa.accmulate.dff_gen[11].d2.D  = _245_ ^ _110_;
	assign _246_ = (_147_ ? _107_ : _151_);
	assign \mchip.aa.accmulate.dff_gen[10].d2.D  = ~(_246_ ^ _102_);
	assign _247_ = (_147_ ? _105_ : _149_);
	assign \mchip.aa.accmulate.dff_gen[9].d2.D  = ~(_247_ ^ _104_);
	assign _248_ = ~_144_;
	assign _249_ = (_138_ ? _121_ : _248_);
	assign \mchip.aa.accmulate.dff_gen[7].d2.D  = _249_ ^ _122_;
	assign _250_ = (_138_ ? _119_ : _142_);
	assign \mchip.aa.accmulate.dff_gen[6].d2.D  = ~(_250_ ^ _114_);
	assign _251_ = (_138_ ? _117_ : _140_);
	assign \mchip.aa.accmulate.dff_gen[5].d2.D  = ~(_251_ ^ _116_);
	assign \mchip.aa.accmulate.dff_gen[3].d2.D  = ~(_135_ ^ _126_);
	assign \mchip.aa.accmulate.dff_gen[2].d2.D  = ~(_133_ ^ _128_);
	assign \mchip.aa.accmulate.dff_gen[1].d2.D  = ~(_131_ ^ _130_);
	assign _252_ = io_in[13] | ~io_in[11];
	assign _000_ = \mchip.control.state [0] & ~_252_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.control.temp_count [0] <= 1'h1;
		else if (_015_)
			\mchip.control.temp_count [0] <= _049_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.control.temp_count [1] <= 1'h0;
		else if (_015_)
			\mchip.control.temp_count [1] <= _050_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.control.temp_count [2] <= 1'h0;
		else if (_015_)
			\mchip.control.temp_count [2] <= _051_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.control.temp_count [3] <= 1'h1;
		else if (_015_)
			\mchip.control.temp_count [3] <= _052_;
	always @(posedge io_in[12]) \mchip.control._do_next  <= io_in[7];
	always @(posedge io_in[12]) \mchip._Finish  <= \mchip.control.state [0];
	always @(posedge io_in[12]) \mchip.shiftin  <= io_in[8];
	always @(posedge io_in[12])
		if (_047_)
			\mchip.op_b_in [0] <= io_in[9];
	always @(posedge io_in[12])
		if (_047_)
			\mchip.op_b_in [1] <= \mchip.op_b_in [0];
	always @(posedge io_in[12])
		if (_047_)
			\mchip.op_b_in [2] <= \mchip.op_b_in [1];
	always @(posedge io_in[12])
		if (_047_)
			\mchip.op_b_in [3] <= \mchip.op_b_in [2];
	always @(posedge io_in[12])
		if (_047_)
			\mchip.op_b_in [4] <= \mchip.op_b_in [3];
	always @(posedge io_in[12])
		if (_047_)
			\mchip.op_b_in [5] <= \mchip.op_b_in [4];
	always @(posedge io_in[12])
		if (_047_)
			\mchip.op_b_in [6] <= \mchip.op_b_in [5];
	always @(posedge io_in[12])
		if (_047_)
			\mchip.op_b_in [7] <= \mchip.op_b_in [6];
	always @(posedge io_in[12])
		if (_047_)
			\mchip.op_a_in [0] <= io_in[10];
	always @(posedge io_in[12])
		if (_047_)
			\mchip.op_a_in [1] <= \mchip.op_a_in [0];
	always @(posedge io_in[12])
		if (_047_)
			\mchip.op_a_in [2] <= \mchip.op_a_in [1];
	always @(posedge io_in[12])
		if (_047_)
			\mchip.op_a_in [3] <= \mchip.op_a_in [2];
	always @(posedge io_in[12])
		if (_047_)
			\mchip.op_a_in [4] <= \mchip.op_a_in [3];
	always @(posedge io_in[12])
		if (_047_)
			\mchip.op_a_in [5] <= \mchip.op_a_in [4];
	always @(posedge io_in[12])
		if (_047_)
			\mchip.op_a_in [6] <= \mchip.op_a_in [5];
	always @(posedge io_in[12])
		if (_047_)
			\mchip.op_a_in [7] <= \mchip.op_a_in [6];
	always @(posedge io_in[12])
		if (_014_)
			\mchip.shiftout [0] <= _028_;
	always @(posedge io_in[12])
		if (_014_)
			\mchip.shiftout [1] <= _038_;
	always @(posedge io_in[12])
		if (_014_)
			\mchip.shiftout [2] <= _039_;
	always @(posedge io_in[12])
		if (_014_)
			\mchip.shiftout [3] <= _040_;
	always @(posedge io_in[12])
		if (_014_)
			\mchip.shiftout [4] <= _041_;
	always @(posedge io_in[12])
		if (_014_)
			\mchip.shiftout [5] <= _042_;
	always @(posedge io_in[12])
		if (_014_)
			\mchip.shiftout [6] <= _043_;
	always @(posedge io_in[12])
		if (_014_)
			\mchip.shiftout [7] <= _044_;
	always @(posedge io_in[12])
		if (_014_)
			\mchip.shiftout [8] <= _045_;
	always @(posedge io_in[12])
		if (_014_)
			\mchip.shiftout [9] <= _046_;
	always @(posedge io_in[12])
		if (_014_)
			\mchip.shiftout [10] <= _029_;
	always @(posedge io_in[12])
		if (_014_)
			\mchip.shiftout [11] <= _030_;
	always @(posedge io_in[12])
		if (_014_)
			\mchip.shiftout [12] <= _031_;
	always @(posedge io_in[12])
		if (_014_)
			\mchip.shiftout [13] <= _032_;
	always @(posedge io_in[12])
		if (_014_)
			\mchip.shiftout [14] <= _033_;
	always @(posedge io_in[12])
		if (_014_)
			\mchip.shiftout [15] <= _034_;
	always @(posedge io_in[12])
		if (_014_)
			\mchip.shiftout [16] <= _035_;
	always @(posedge io_in[12])
		if (_014_)
			\mchip.shiftout [17] <= _036_;
	always @(posedge io_in[12])
		if (_014_)
			\mchip.shiftout [18] <= _037_;
	always @(posedge io_in[12])
		if (_014_)
			if (!_048_)
				\mchip.shiftout [19] <= 1'h0;
			else
				\mchip.shiftout [19] <= \mchip.aa.accmulate.dff_gen[19].d2.Q ;
	always @(posedge \mchip.control.state [2])
		if (_012_)
			\mchip.opb.dff_gen[7].d1.Q  <= 1'h0;
		else
			\mchip.opb.dff_gen[7].d1.Q  <= \mchip.op_b_in [7];
	always @(posedge \mchip.control.state [5])
		if (_012_)
			\mchip.aa.i0.dff_gen[14].d2.Q  <= 1'h0;
		else
			\mchip.aa.i0.dff_gen[14].d2.Q  <= \mchip.mult.i3.temp_register [14];
	always @(posedge \mchip.control.state [5])
		if (_012_)
			\mchip.aa.i0.dff_gen[13].d2.Q  <= 1'h0;
		else
			\mchip.aa.i0.dff_gen[13].d2.Q  <= \mchip.mult.i3.temp_register [13];
	always @(posedge \mchip.control.state [5])
		if (_012_)
			\mchip.aa.i0.dff_gen[12].d2.Q  <= 1'h0;
		else
			\mchip.aa.i0.dff_gen[12].d2.Q  <= \mchip.mult.i3.temp_register [12];
	always @(posedge \mchip.control.state [5])
		if (_012_)
			\mchip.aa.i0.dff_gen[11].d2.Q  <= 1'h0;
		else
			\mchip.aa.i0.dff_gen[11].d2.Q  <= \mchip.mult.i3.temp_register [11];
	always @(posedge \mchip.control.state [5])
		if (_012_)
			\mchip.aa.i0.dff_gen[10].d2.Q  <= 1'h0;
		else
			\mchip.aa.i0.dff_gen[10].d2.Q  <= \mchip.mult.i3.temp_register [10];
	always @(posedge \mchip.control.state [5])
		if (_012_)
			\mchip.aa.i0.dff_gen[0].d2.Q  <= 1'h0;
		else
			\mchip.aa.i0.dff_gen[0].d2.Q  <= \mchip.mult.i3.temp_register [0];
	always @(posedge \mchip.control.state [5])
		if (_012_)
			\mchip.aa.i0.dff_gen[8].d2.Q  <= 1'h0;
		else
			\mchip.aa.i0.dff_gen[8].d2.Q  <= \mchip.mult.i3.temp_register [8];
	always @(posedge \mchip.control.state [5])
		if (_012_)
			\mchip.aa.i0.dff_gen[7].d2.Q  <= 1'h0;
		else
			\mchip.aa.i0.dff_gen[7].d2.Q  <= \mchip.mult.i3.temp_register [7];
	always @(posedge \mchip.control.state [5])
		if (_012_)
			\mchip.aa.i0.dff_gen[6].d2.Q  <= 1'h0;
		else
			\mchip.aa.i0.dff_gen[6].d2.Q  <= \mchip.mult.i3.temp_register [6];
	always @(posedge \mchip.control.state [5])
		if (_012_)
			\mchip.aa.i0.dff_gen[5].d2.Q  <= 1'h0;
		else
			\mchip.aa.i0.dff_gen[5].d2.Q  <= \mchip.mult.i3.temp_register [5];
	always @(posedge \mchip.control.state [5])
		if (_012_)
			\mchip.aa.i0.dff_gen[4].d2.Q  <= 1'h0;
		else
			\mchip.aa.i0.dff_gen[4].d2.Q  <= \mchip.mult.i3.temp_register [4];
	always @(posedge \mchip.control.state [5])
		if (_012_)
			\mchip.aa.i0.dff_gen[3].d2.Q  <= 1'h0;
		else
			\mchip.aa.i0.dff_gen[3].d2.Q  <= \mchip.mult.i3.temp_register [3];
	always @(posedge \mchip.control.state [5])
		if (_012_)
			\mchip.aa.i0.dff_gen[2].d2.Q  <= 1'h0;
		else
			\mchip.aa.i0.dff_gen[2].d2.Q  <= \mchip.mult.i3.temp_register [2];
	always @(posedge \mchip.control.state [5])
		if (_012_)
			\mchip.aa.i0.dff_gen[1].d2.Q  <= 1'h0;
		else
			\mchip.aa.i0.dff_gen[1].d2.Q  <= \mchip.mult.i3.temp_register [1];
	always @(posedge \mchip.control.state [5])
		if (_012_)
			\mchip.aa.i0.dff_gen[15].d2.Q  <= 1'h0;
		else
			\mchip.aa.i0.dff_gen[15].d2.Q  <= \mchip.mult.i3.temp_register [15];
	always @(negedge \mchip.control.state [5])
		if (_012_)
			\mchip.aa.accmulate.dff_gen[9].d2.Q  <= 1'h0;
		else
			\mchip.aa.accmulate.dff_gen[9].d2.Q  <= \mchip.aa.accmulate.dff_gen[9].d2.D ;
	always @(posedge io_in[12]) \mchip.mult.i0.state [0] <= _009_;
	always @(posedge io_in[12]) \mchip.mult.i0.state [1] <= _010_;
	always @(posedge io_in[12]) \mchip.mult.i0.state [2] <= _011_;
	always @(posedge io_in[12]) \mchip.mult.i0.state [3] <= _003_;
	always @(posedge io_in[12]) \mchip.mult.i0.state [4] <= _004_;
	always @(posedge io_in[12]) \mchip.control.state [0] <= _005_;
	always @(posedge io_in[12]) \mchip.control.state [1] <= _006_;
	always @(posedge io_in[12]) \mchip.control.state [2] <= _007_;
	always @(posedge io_in[12]) \mchip.control.state [3] <= _008_;
	always @(posedge io_in[12]) \mchip.control.state [4] <= _000_;
	always @(posedge io_in[12]) \mchip.control.state [5] <= _001_;
	always @(posedge io_in[12]) \mchip.control.state [6] <= _002_;
	always @(negedge \mchip.control.state [5])
		if (_012_)
			\mchip.aa.accmulate.dff_gen[19].d2.Q  <= 1'h0;
		else if (\mchip.aa.adder.S4.carry_in )
			\mchip.aa.accmulate.dff_gen[19].d2.Q  <= \mchip.aa.adder.S4.S1.fa3.sum ;
	always @(negedge \mchip.control.state [5])
		if (_012_)
			\mchip.aa.accmulate.dff_gen[18].d2.Q  <= 1'h0;
		else if (\mchip.aa.adder.S4.carry_in )
			\mchip.aa.accmulate.dff_gen[18].d2.Q  <= \mchip.aa.adder.S4.S1.fa2.sum ;
	always @(negedge \mchip.control.state [5])
		if (_012_)
			\mchip.aa.accmulate.dff_gen[17].d2.Q  <= 1'h0;
		else if (\mchip.aa.adder.S4.carry_in )
			\mchip.aa.accmulate.dff_gen[17].d2.Q  <= \mchip.aa.adder.S4.S1.fa1.sum ;
	always @(negedge \mchip.control.state [5])
		if (_012_)
			\mchip.aa.accmulate.dff_gen[16].d2.Q  <= 1'h0;
		else if (\mchip.aa.adder.S4.carry_in )
			\mchip.aa.accmulate.dff_gen[16].d2.Q  <= \mchip.aa.adder.S4.S1.fa0.sum ;
	always @(negedge \mchip.control.state [5])
		if (_012_)
			\mchip.aa.accmulate.dff_gen[14].d2.Q  <= 1'h0;
		else
			\mchip.aa.accmulate.dff_gen[14].d2.Q  <= \mchip.aa.accmulate.dff_gen[14].d2.D ;
	always @(negedge \mchip.control.state [5])
		if (_012_)
			\mchip.aa.accmulate.dff_gen[13].d2.Q  <= 1'h0;
		else
			\mchip.aa.accmulate.dff_gen[13].d2.Q  <= \mchip.aa.accmulate.dff_gen[13].d2.D ;
	always @(negedge \mchip.control.state [5])
		if (_012_)
			\mchip.aa.accmulate.dff_gen[12].d2.Q  <= 1'h0;
		else
			\mchip.aa.accmulate.dff_gen[12].d2.Q  <= \mchip.aa.accmulate.dff_gen[12].d2.D ;
	always @(negedge \mchip.control.state [5])
		if (_012_)
			\mchip.aa.accmulate.dff_gen[11].d2.Q  <= 1'h0;
		else
			\mchip.aa.accmulate.dff_gen[11].d2.Q  <= \mchip.aa.accmulate.dff_gen[11].d2.D ;
	always @(negedge \mchip.control.state [5])
		if (_012_)
			\mchip.aa.accmulate.dff_gen[10].d2.Q  <= 1'h0;
		else
			\mchip.aa.accmulate.dff_gen[10].d2.Q  <= \mchip.aa.accmulate.dff_gen[10].d2.D ;
	always @(negedge \mchip.control.state [5])
		if (_012_)
			\mchip.aa.accmulate.dff_gen[0].d2.Q  <= 1'h0;
		else
			\mchip.aa.accmulate.dff_gen[0].d2.Q  <= \mchip.aa.accmulate.dff_gen[0].d2.D ;
	always @(negedge \mchip.control.state [5])
		if (_012_)
			\mchip.aa.accmulate.dff_gen[8].d2.Q  <= 1'h0;
		else
			\mchip.aa.accmulate.dff_gen[8].d2.Q  <= \mchip.aa.accmulate.dff_gen[8].d2.D ;
	always @(negedge \mchip.control.state [5])
		if (_012_)
			\mchip.aa.accmulate.dff_gen[7].d2.Q  <= 1'h0;
		else
			\mchip.aa.accmulate.dff_gen[7].d2.Q  <= \mchip.aa.accmulate.dff_gen[7].d2.D ;
	always @(negedge \mchip.control.state [5])
		if (_012_)
			\mchip.aa.accmulate.dff_gen[6].d2.Q  <= 1'h0;
		else
			\mchip.aa.accmulate.dff_gen[6].d2.Q  <= \mchip.aa.accmulate.dff_gen[6].d2.D ;
	always @(negedge \mchip.control.state [5])
		if (_012_)
			\mchip.aa.accmulate.dff_gen[5].d2.Q  <= 1'h0;
		else
			\mchip.aa.accmulate.dff_gen[5].d2.Q  <= \mchip.aa.accmulate.dff_gen[5].d2.D ;
	always @(negedge \mchip.control.state [5])
		if (_012_)
			\mchip.aa.accmulate.dff_gen[4].d2.Q  <= 1'h0;
		else
			\mchip.aa.accmulate.dff_gen[4].d2.Q  <= \mchip.aa.accmulate.dff_gen[4].d2.D ;
	always @(negedge \mchip.control.state [5])
		if (_012_)
			\mchip.aa.accmulate.dff_gen[3].d2.Q  <= 1'h0;
		else
			\mchip.aa.accmulate.dff_gen[3].d2.Q  <= \mchip.aa.accmulate.dff_gen[3].d2.D ;
	always @(negedge \mchip.control.state [5])
		if (_012_)
			\mchip.aa.accmulate.dff_gen[2].d2.Q  <= 1'h0;
		else
			\mchip.aa.accmulate.dff_gen[2].d2.Q  <= \mchip.aa.accmulate.dff_gen[2].d2.D ;
	always @(negedge \mchip.control.state [5])
		if (_012_)
			\mchip.aa.accmulate.dff_gen[1].d2.Q  <= 1'h0;
		else
			\mchip.aa.accmulate.dff_gen[1].d2.Q  <= \mchip.aa.accmulate.dff_gen[1].d2.D ;
	always @(negedge \mchip.control.state [5])
		if (_012_)
			\mchip.aa.accmulate.dff_gen[15].d2.Q  <= 1'h0;
		else
			\mchip.aa.accmulate.dff_gen[15].d2.Q  <= \mchip.aa.accmulate.dff_gen[15].d2.D ;
	always @(posedge io_in[12])
		if (_012_)
			\mchip.mult.i0.temp_count [0] <= 1'h0;
		else if (\mchip.mult.i0.state [1])
			\mchip.mult.i0.temp_count [0] <= _017_;
	always @(posedge io_in[12])
		if (_012_)
			\mchip.mult.i0.temp_count [1] <= 1'h0;
		else if (\mchip.mult.i0.state [1])
			\mchip.mult.i0.temp_count [1] <= _018_;
	always @(posedge io_in[12])
		if (_012_)
			\mchip.mult.i0.temp_count [2] <= 1'h0;
		else if (\mchip.mult.i0.state [1])
			\mchip.mult.i0.temp_count [2] <= _019_;
	reg \mchip.mult.i3.temp_register_reg[8] ;
	always @(posedge io_in[12])
		if (_016_)
			\mchip.mult.i3.temp_register_reg[8]  <= 1'h0;
		else if (\mchip.mult.i0.state [1])
			\mchip.mult.i3.temp_register_reg[8]  <= _020_;
	assign \mchip.mult.i3.temp_register [8] = \mchip.mult.i3.temp_register_reg[8] ;
	reg \mchip.mult.i3.temp_register_reg[9] ;
	always @(posedge io_in[12])
		if (_016_)
			\mchip.mult.i3.temp_register_reg[9]  <= 1'h0;
		else if (\mchip.mult.i0.state [1])
			\mchip.mult.i3.temp_register_reg[9]  <= _021_;
	assign \mchip.mult.i3.temp_register [9] = \mchip.mult.i3.temp_register_reg[9] ;
	reg \mchip.mult.i3.temp_register_reg[10] ;
	always @(posedge io_in[12])
		if (_016_)
			\mchip.mult.i3.temp_register_reg[10]  <= 1'h0;
		else if (\mchip.mult.i0.state [1])
			\mchip.mult.i3.temp_register_reg[10]  <= _022_;
	assign \mchip.mult.i3.temp_register [10] = \mchip.mult.i3.temp_register_reg[10] ;
	reg \mchip.mult.i3.temp_register_reg[11] ;
	always @(posedge io_in[12])
		if (_016_)
			\mchip.mult.i3.temp_register_reg[11]  <= 1'h0;
		else if (\mchip.mult.i0.state [1])
			\mchip.mult.i3.temp_register_reg[11]  <= _023_;
	assign \mchip.mult.i3.temp_register [11] = \mchip.mult.i3.temp_register_reg[11] ;
	reg \mchip.mult.i3.temp_register_reg[12] ;
	always @(posedge io_in[12])
		if (_016_)
			\mchip.mult.i3.temp_register_reg[12]  <= 1'h0;
		else if (\mchip.mult.i0.state [1])
			\mchip.mult.i3.temp_register_reg[12]  <= _024_;
	assign \mchip.mult.i3.temp_register [12] = \mchip.mult.i3.temp_register_reg[12] ;
	reg \mchip.mult.i3.temp_register_reg[13] ;
	always @(posedge io_in[12])
		if (_016_)
			\mchip.mult.i3.temp_register_reg[13]  <= 1'h0;
		else if (\mchip.mult.i0.state [1])
			\mchip.mult.i3.temp_register_reg[13]  <= _025_;
	assign \mchip.mult.i3.temp_register [13] = \mchip.mult.i3.temp_register_reg[13] ;
	reg \mchip.mult.i3.temp_register_reg[14] ;
	always @(posedge io_in[12])
		if (_016_)
			\mchip.mult.i3.temp_register_reg[14]  <= 1'h0;
		else if (\mchip.mult.i0.state [1])
			\mchip.mult.i3.temp_register_reg[14]  <= _026_;
	assign \mchip.mult.i3.temp_register [14] = \mchip.mult.i3.temp_register_reg[14] ;
	reg \mchip.mult.i3.temp_register_reg[15] ;
	always @(posedge io_in[12])
		if (_016_)
			\mchip.mult.i3.temp_register_reg[15]  <= 1'h0;
		else if (\mchip.mult.i0.state [1])
			\mchip.mult.i3.temp_register_reg[15]  <= _027_;
	assign \mchip.mult.i3.temp_register [15] = \mchip.mult.i3.temp_register_reg[15] ;
	always @(posedge \mchip.control.state [5])
		if (_012_)
			\mchip.aa.i0.dff_gen[9].d2.Q  <= 1'h0;
		else
			\mchip.aa.i0.dff_gen[9].d2.Q  <= \mchip.mult.i3.temp_register [9];
	always @(posedge \mchip.mult.i0.state [3])
		if (_012_)
			\mchip.mult.i1.r1.dff_gen[0].d1.Q  <= 1'h0;
		else
			\mchip.mult.i1.r1.dff_gen[0].d1.Q  <= \mchip.opa.dff_gen[0].d1.Q ;
	always @(posedge \mchip.mult.i0.state [3])
		if (_012_)
			\mchip.mult.i1.r1.dff_gen[1].d1.Q  <= 1'h0;
		else
			\mchip.mult.i1.r1.dff_gen[1].d1.Q  <= \mchip.opa.dff_gen[1].d1.Q ;
	always @(posedge \mchip.mult.i0.state [3])
		if (_012_)
			\mchip.mult.i1.r1.dff_gen[2].d1.Q  <= 1'h0;
		else
			\mchip.mult.i1.r1.dff_gen[2].d1.Q  <= \mchip.opa.dff_gen[2].d1.Q ;
	always @(posedge \mchip.mult.i0.state [3])
		if (_012_)
			\mchip.mult.i1.r1.dff_gen[3].d1.Q  <= 1'h0;
		else
			\mchip.mult.i1.r1.dff_gen[3].d1.Q  <= \mchip.opa.dff_gen[3].d1.Q ;
	always @(posedge \mchip.mult.i0.state [3])
		if (_012_)
			\mchip.mult.i1.r1.dff_gen[4].d1.Q  <= 1'h0;
		else
			\mchip.mult.i1.r1.dff_gen[4].d1.Q  <= \mchip.opa.dff_gen[4].d1.Q ;
	always @(posedge \mchip.mult.i0.state [3])
		if (_012_)
			\mchip.mult.i1.r1.dff_gen[5].d1.Q  <= 1'h0;
		else
			\mchip.mult.i1.r1.dff_gen[5].d1.Q  <= \mchip.opa.dff_gen[5].d1.Q ;
	always @(posedge \mchip.mult.i0.state [3])
		if (_012_)
			\mchip.mult.i1.r1.dff_gen[6].d1.Q  <= 1'h0;
		else
			\mchip.mult.i1.r1.dff_gen[6].d1.Q  <= \mchip.opa.dff_gen[6].d1.Q ;
	always @(posedge io_in[12])
		if (_012_)
			\mchip.mult.i3.temp_Add  <= 1'h0;
		else if (!\mchip.mult.i0.state [3])
			\mchip.mult.i3.temp_Add  <= _053_;
	always @(posedge \mchip.control.state [2])
		if (_012_)
			\mchip.opa.dff_gen[7].d1.Q  <= 1'h0;
		else
			\mchip.opa.dff_gen[7].d1.Q  <= \mchip.op_a_in [7];
	always @(posedge \mchip.control.state [2])
		if (_012_)
			\mchip.opb.dff_gen[0].d1.Q  <= 1'h0;
		else
			\mchip.opb.dff_gen[0].d1.Q  <= \mchip.op_b_in [0];
	always @(posedge \mchip.control.state [2])
		if (_012_)
			\mchip.opb.dff_gen[1].d1.Q  <= 1'h0;
		else
			\mchip.opb.dff_gen[1].d1.Q  <= \mchip.op_b_in [1];
	always @(posedge \mchip.control.state [2])
		if (_012_)
			\mchip.opb.dff_gen[2].d1.Q  <= 1'h0;
		else
			\mchip.opb.dff_gen[2].d1.Q  <= \mchip.op_b_in [2];
	always @(posedge \mchip.control.state [2])
		if (_012_)
			\mchip.opb.dff_gen[3].d1.Q  <= 1'h0;
		else
			\mchip.opb.dff_gen[3].d1.Q  <= \mchip.op_b_in [3];
	always @(posedge \mchip.control.state [2])
		if (_012_)
			\mchip.opb.dff_gen[4].d1.Q  <= 1'h0;
		else
			\mchip.opb.dff_gen[4].d1.Q  <= \mchip.op_b_in [4];
	always @(posedge \mchip.control.state [2])
		if (_012_)
			\mchip.opb.dff_gen[5].d1.Q  <= 1'h0;
		else
			\mchip.opb.dff_gen[5].d1.Q  <= \mchip.op_b_in [5];
	always @(posedge \mchip.control.state [2])
		if (_012_)
			\mchip.opb.dff_gen[6].d1.Q  <= 1'h0;
		else
			\mchip.opb.dff_gen[6].d1.Q  <= \mchip.op_b_in [6];
	always @(posedge \mchip.mult.i0.state [3])
		if (_012_)
			\mchip.mult.i1.r1.dff_gen[7].d1.Q  <= 1'h0;
		else
			\mchip.mult.i1.r1.dff_gen[7].d1.Q  <= \mchip.opa.dff_gen[7].d1.Q ;
	always @(posedge \mchip.control.state [2])
		if (_012_)
			\mchip.opa.dff_gen[0].d1.Q  <= 1'h0;
		else
			\mchip.opa.dff_gen[0].d1.Q  <= \mchip.op_a_in [0];
	always @(posedge \mchip.control.state [2])
		if (_012_)
			\mchip.opa.dff_gen[1].d1.Q  <= 1'h0;
		else
			\mchip.opa.dff_gen[1].d1.Q  <= \mchip.op_a_in [1];
	always @(posedge \mchip.control.state [2])
		if (_012_)
			\mchip.opa.dff_gen[2].d1.Q  <= 1'h0;
		else
			\mchip.opa.dff_gen[2].d1.Q  <= \mchip.op_a_in [2];
	always @(posedge \mchip.control.state [2])
		if (_012_)
			\mchip.opa.dff_gen[3].d1.Q  <= 1'h0;
		else
			\mchip.opa.dff_gen[3].d1.Q  <= \mchip.op_a_in [3];
	always @(posedge \mchip.control.state [2])
		if (_012_)
			\mchip.opa.dff_gen[4].d1.Q  <= 1'h0;
		else
			\mchip.opa.dff_gen[4].d1.Q  <= \mchip.op_a_in [4];
	always @(posedge \mchip.control.state [2])
		if (_012_)
			\mchip.opa.dff_gen[5].d1.Q  <= 1'h0;
		else
			\mchip.opa.dff_gen[5].d1.Q  <= \mchip.op_a_in [5];
	always @(posedge \mchip.control.state [2])
		if (_012_)
			\mchip.opa.dff_gen[6].d1.Q  <= 1'h0;
		else
			\mchip.opa.dff_gen[6].d1.Q  <= \mchip.op_a_in [6];
	reg \mchip.mult.i3.temp_register_reg[0] ;
	always @(posedge io_in[12])
		if (_012_)
			\mchip.mult.i3.temp_register_reg[0]  <= 1'h0;
		else if (_013_)
			\mchip.mult.i3.temp_register_reg[0]  <= _054_;
	assign \mchip.mult.i3.temp_register [0] = \mchip.mult.i3.temp_register_reg[0] ;
	reg \mchip.mult.i3.temp_register_reg[1] ;
	always @(posedge io_in[12])
		if (_012_)
			\mchip.mult.i3.temp_register_reg[1]  <= 1'h0;
		else if (_013_)
			\mchip.mult.i3.temp_register_reg[1]  <= _055_;
	assign \mchip.mult.i3.temp_register [1] = \mchip.mult.i3.temp_register_reg[1] ;
	reg \mchip.mult.i3.temp_register_reg[2] ;
	always @(posedge io_in[12])
		if (_012_)
			\mchip.mult.i3.temp_register_reg[2]  <= 1'h0;
		else if (_013_)
			\mchip.mult.i3.temp_register_reg[2]  <= _056_;
	assign \mchip.mult.i3.temp_register [2] = \mchip.mult.i3.temp_register_reg[2] ;
	reg \mchip.mult.i3.temp_register_reg[3] ;
	always @(posedge io_in[12])
		if (_012_)
			\mchip.mult.i3.temp_register_reg[3]  <= 1'h0;
		else if (_013_)
			\mchip.mult.i3.temp_register_reg[3]  <= _057_;
	assign \mchip.mult.i3.temp_register [3] = \mchip.mult.i3.temp_register_reg[3] ;
	reg \mchip.mult.i3.temp_register_reg[4] ;
	always @(posedge io_in[12])
		if (_012_)
			\mchip.mult.i3.temp_register_reg[4]  <= 1'h0;
		else if (_013_)
			\mchip.mult.i3.temp_register_reg[4]  <= _058_;
	assign \mchip.mult.i3.temp_register [4] = \mchip.mult.i3.temp_register_reg[4] ;
	reg \mchip.mult.i3.temp_register_reg[5] ;
	always @(posedge io_in[12])
		if (_012_)
			\mchip.mult.i3.temp_register_reg[5]  <= 1'h0;
		else if (_013_)
			\mchip.mult.i3.temp_register_reg[5]  <= _059_;
	assign \mchip.mult.i3.temp_register [5] = \mchip.mult.i3.temp_register_reg[5] ;
	reg \mchip.mult.i3.temp_register_reg[6] ;
	always @(posedge io_in[12])
		if (_012_)
			\mchip.mult.i3.temp_register_reg[6]  <= 1'h0;
		else if (_013_)
			\mchip.mult.i3.temp_register_reg[6]  <= _060_;
	assign \mchip.mult.i3.temp_register [6] = \mchip.mult.i3.temp_register_reg[6] ;
	reg \mchip.mult.i3.temp_register_reg[7] ;
	always @(posedge io_in[12])
		if (_012_)
			\mchip.mult.i3.temp_register_reg[7]  <= 1'h0;
		else if (_013_)
			\mchip.mult.i3.temp_register_reg[7]  <= _061_;
	assign \mchip.mult.i3.temp_register [7] = \mchip.mult.i3.temp_register_reg[7] ;
	assign io_out = {2'h0, \mchip.aa.adder.S4.carry_out , \mchip.control.state [0], \mchip.shiftout [0], \mchip.mult.i0.state [0], 8'h00};
	assign \mchip.Begin_mul  = \mchip.control.state [6];
	assign \mchip.End_mul  = \mchip.mult.i0.state [0];
	assign \mchip.Finish  = \mchip.control.state [0];
	assign \mchip.Load_op  = \mchip.control.state [2];
	assign \mchip.START  = io_in[11];
	assign \mchip.aa.accmulate.in  = {4'h0, \mchip.aa.accmulate.dff_gen[15].d2.D , \mchip.aa.accmulate.dff_gen[14].d2.D , \mchip.aa.accmulate.dff_gen[13].d2.D , \mchip.aa.accmulate.dff_gen[12].d2.D , \mchip.aa.accmulate.dff_gen[11].d2.D , \mchip.aa.accmulate.dff_gen[10].d2.D , \mchip.aa.accmulate.dff_gen[9].d2.D , \mchip.aa.accmulate.dff_gen[8].d2.D , \mchip.aa.accmulate.dff_gen[7].d2.D , \mchip.aa.accmulate.dff_gen[6].d2.D , \mchip.aa.accmulate.dff_gen[5].d2.D , \mchip.aa.accmulate.dff_gen[4].d2.D , \mchip.aa.accmulate.dff_gen[3].d2.D , \mchip.aa.accmulate.dff_gen[2].d2.D , \mchip.aa.accmulate.dff_gen[1].d2.D , \mchip.aa.accmulate.dff_gen[0].d2.D };
	assign \mchip.aa.accmulate.out  = {\mchip.aa.accmulate.dff_gen[19].d2.Q , \mchip.aa.accmulate.dff_gen[18].d2.Q , \mchip.aa.accmulate.dff_gen[17].d2.Q , \mchip.aa.accmulate.dff_gen[16].d2.Q , \mchip.aa.accmulate.dff_gen[15].d2.Q , \mchip.aa.accmulate.dff_gen[14].d2.Q , \mchip.aa.accmulate.dff_gen[13].d2.Q , \mchip.aa.accmulate.dff_gen[12].d2.Q , \mchip.aa.accmulate.dff_gen[11].d2.Q , \mchip.aa.accmulate.dff_gen[10].d2.Q , \mchip.aa.accmulate.dff_gen[9].d2.Q , \mchip.aa.accmulate.dff_gen[8].d2.Q , \mchip.aa.accmulate.dff_gen[7].d2.Q , \mchip.aa.accmulate.dff_gen[6].d2.Q , \mchip.aa.accmulate.dff_gen[5].d2.Q , \mchip.aa.accmulate.dff_gen[4].d2.Q , \mchip.aa.accmulate.dff_gen[3].d2.Q , \mchip.aa.accmulate.dff_gen[2].d2.Q , \mchip.aa.accmulate.dff_gen[1].d2.Q , \mchip.aa.accmulate.dff_gen[0].d2.Q };
	assign \mchip.aa.accmulate.temp_out  = {\mchip.aa.accmulate.dff_gen[19].d2.Q , \mchip.aa.accmulate.dff_gen[18].d2.Q , \mchip.aa.accmulate.dff_gen[17].d2.Q , \mchip.aa.accmulate.dff_gen[16].d2.Q , \mchip.aa.accmulate.dff_gen[15].d2.Q , \mchip.aa.accmulate.dff_gen[14].d2.Q , \mchip.aa.accmulate.dff_gen[13].d2.Q , \mchip.aa.accmulate.dff_gen[12].d2.Q , \mchip.aa.accmulate.dff_gen[11].d2.Q , \mchip.aa.accmulate.dff_gen[10].d2.Q , \mchip.aa.accmulate.dff_gen[9].d2.Q , \mchip.aa.accmulate.dff_gen[8].d2.Q , \mchip.aa.accmulate.dff_gen[7].d2.Q , \mchip.aa.accmulate.dff_gen[6].d2.Q , \mchip.aa.accmulate.dff_gen[5].d2.Q , \mchip.aa.accmulate.dff_gen[4].d2.Q , \mchip.aa.accmulate.dff_gen[3].d2.Q , \mchip.aa.accmulate.dff_gen[2].d2.Q , \mchip.aa.accmulate.dff_gen[1].d2.Q , \mchip.aa.accmulate.dff_gen[0].d2.Q };
	assign \mchip.aa.add  = \mchip.control.state [5];
	assign \mchip.aa.add_in  = {\mchip.aa.accmulate.dff_gen[19].d2.Q , \mchip.aa.accmulate.dff_gen[18].d2.Q , \mchip.aa.accmulate.dff_gen[17].d2.Q , \mchip.aa.accmulate.dff_gen[16].d2.Q , \mchip.aa.accmulate.dff_gen[15].d2.Q , \mchip.aa.accmulate.dff_gen[14].d2.Q , \mchip.aa.accmulate.dff_gen[13].d2.Q , \mchip.aa.accmulate.dff_gen[12].d2.Q , \mchip.aa.accmulate.dff_gen[11].d2.Q , \mchip.aa.accmulate.dff_gen[10].d2.Q , \mchip.aa.accmulate.dff_gen[9].d2.Q , \mchip.aa.accmulate.dff_gen[8].d2.Q , \mchip.aa.accmulate.dff_gen[7].d2.Q , \mchip.aa.accmulate.dff_gen[6].d2.Q , \mchip.aa.accmulate.dff_gen[5].d2.Q , \mchip.aa.accmulate.dff_gen[4].d2.Q , \mchip.aa.accmulate.dff_gen[3].d2.Q , \mchip.aa.accmulate.dff_gen[2].d2.Q , \mchip.aa.accmulate.dff_gen[1].d2.Q , \mchip.aa.accmulate.dff_gen[0].d2.Q };
	assign \mchip.aa.add_out  = {4'h0, \mchip.aa.accmulate.dff_gen[15].d2.D , \mchip.aa.accmulate.dff_gen[14].d2.D , \mchip.aa.accmulate.dff_gen[13].d2.D , \mchip.aa.accmulate.dff_gen[12].d2.D , \mchip.aa.accmulate.dff_gen[11].d2.D , \mchip.aa.accmulate.dff_gen[10].d2.D , \mchip.aa.accmulate.dff_gen[9].d2.D , \mchip.aa.accmulate.dff_gen[8].d2.D , \mchip.aa.accmulate.dff_gen[7].d2.D , \mchip.aa.accmulate.dff_gen[6].d2.D , \mchip.aa.accmulate.dff_gen[5].d2.D , \mchip.aa.accmulate.dff_gen[4].d2.D , \mchip.aa.accmulate.dff_gen[3].d2.D , \mchip.aa.accmulate.dff_gen[2].d2.D , \mchip.aa.accmulate.dff_gen[1].d2.D , \mchip.aa.accmulate.dff_gen[0].d2.D };
	assign \mchip.aa.adder.S0.S0.a  = {\mchip.aa.i0.dff_gen[3].d2.Q , \mchip.aa.i0.dff_gen[2].d2.Q , \mchip.aa.i0.dff_gen[1].d2.Q , \mchip.aa.i0.dff_gen[0].d2.Q };
	assign \mchip.aa.adder.S0.S0.b  = {\mchip.aa.accmulate.dff_gen[3].d2.Q , \mchip.aa.accmulate.dff_gen[2].d2.Q , \mchip.aa.accmulate.dff_gen[1].d2.Q , \mchip.aa.accmulate.dff_gen[0].d2.Q };
	assign \mchip.aa.adder.S0.S0.carry_in  = 1'h0;
	assign \mchip.aa.adder.S0.S0.fa0.a  = \mchip.aa.i0.dff_gen[0].d2.Q ;
	assign \mchip.aa.adder.S0.S0.fa0.b  = \mchip.aa.accmulate.dff_gen[0].d2.Q ;
	assign \mchip.aa.adder.S0.S0.fa0.carry_in  = 1'h0;
	assign \mchip.aa.adder.S0.S0.fa0.sum  = \mchip.aa.accmulate.dff_gen[0].d2.D ;
	assign \mchip.aa.adder.S0.S0.fa0.w1  = \mchip.aa.accmulate.dff_gen[0].d2.D ;
	assign \mchip.aa.adder.S0.S0.fa0.w3  = 1'h0;
	assign \mchip.aa.adder.S0.S0.fa1.a  = \mchip.aa.i0.dff_gen[1].d2.Q ;
	assign \mchip.aa.adder.S0.S0.fa1.b  = \mchip.aa.accmulate.dff_gen[1].d2.Q ;
	assign \mchip.aa.adder.S0.S0.fa1.sum  = \mchip.aa.accmulate.dff_gen[1].d2.D ;
	assign \mchip.aa.adder.S0.S0.fa2.a  = \mchip.aa.i0.dff_gen[2].d2.Q ;
	assign \mchip.aa.adder.S0.S0.fa2.b  = \mchip.aa.accmulate.dff_gen[2].d2.Q ;
	assign \mchip.aa.adder.S0.S0.fa2.sum  = \mchip.aa.accmulate.dff_gen[2].d2.D ;
	assign \mchip.aa.adder.S0.S0.fa3.a  = \mchip.aa.i0.dff_gen[3].d2.Q ;
	assign \mchip.aa.adder.S0.S0.fa3.b  = \mchip.aa.accmulate.dff_gen[3].d2.Q ;
	assign \mchip.aa.adder.S0.S0.fa3.sum  = \mchip.aa.accmulate.dff_gen[3].d2.D ;
	assign \mchip.aa.adder.S0.S0.sum  = {\mchip.aa.accmulate.dff_gen[3].d2.D , \mchip.aa.accmulate.dff_gen[2].d2.D , \mchip.aa.accmulate.dff_gen[1].d2.D , \mchip.aa.accmulate.dff_gen[0].d2.D };
	assign \mchip.aa.adder.S0.S1.a  = {\mchip.aa.i0.dff_gen[3].d2.Q , \mchip.aa.i0.dff_gen[2].d2.Q , \mchip.aa.i0.dff_gen[1].d2.Q , \mchip.aa.i0.dff_gen[0].d2.Q };
	assign \mchip.aa.adder.S0.S1.b  = {\mchip.aa.accmulate.dff_gen[3].d2.Q , \mchip.aa.accmulate.dff_gen[2].d2.Q , \mchip.aa.accmulate.dff_gen[1].d2.Q , \mchip.aa.accmulate.dff_gen[0].d2.Q };
	assign \mchip.aa.adder.S0.S1.carry_in  = 1'h1;
	assign \mchip.aa.adder.S0.S1.fa0.a  = \mchip.aa.i0.dff_gen[0].d2.Q ;
	assign \mchip.aa.adder.S0.S1.fa0.b  = \mchip.aa.accmulate.dff_gen[0].d2.Q ;
	assign \mchip.aa.adder.S0.S1.fa0.carry_in  = 1'h1;
	assign \mchip.aa.adder.S0.S1.fa1.a  = \mchip.aa.i0.dff_gen[1].d2.Q ;
	assign \mchip.aa.adder.S0.S1.fa1.b  = \mchip.aa.accmulate.dff_gen[1].d2.Q ;
	assign \mchip.aa.adder.S0.S1.fa2.a  = \mchip.aa.i0.dff_gen[2].d2.Q ;
	assign \mchip.aa.adder.S0.S1.fa2.b  = \mchip.aa.accmulate.dff_gen[2].d2.Q ;
	assign \mchip.aa.adder.S0.S1.fa3.a  = \mchip.aa.i0.dff_gen[3].d2.Q ;
	assign \mchip.aa.adder.S0.S1.fa3.b  = \mchip.aa.accmulate.dff_gen[3].d2.Q ;
	assign \mchip.aa.adder.S0.SUM0  = {\mchip.aa.accmulate.dff_gen[3].d2.D , \mchip.aa.accmulate.dff_gen[2].d2.D , \mchip.aa.accmulate.dff_gen[1].d2.D , \mchip.aa.accmulate.dff_gen[0].d2.D };
	assign \mchip.aa.adder.S0.a  = {\mchip.aa.i0.dff_gen[3].d2.Q , \mchip.aa.i0.dff_gen[2].d2.Q , \mchip.aa.i0.dff_gen[1].d2.Q , \mchip.aa.i0.dff_gen[0].d2.Q };
	assign \mchip.aa.adder.S0.b  = {\mchip.aa.accmulate.dff_gen[3].d2.Q , \mchip.aa.accmulate.dff_gen[2].d2.Q , \mchip.aa.accmulate.dff_gen[1].d2.Q , \mchip.aa.accmulate.dff_gen[0].d2.Q };
	assign \mchip.aa.adder.S0.carry_in  = 1'h0;
	assign \mchip.aa.adder.S0.sum  = {\mchip.aa.accmulate.dff_gen[3].d2.D , \mchip.aa.accmulate.dff_gen[2].d2.D , \mchip.aa.accmulate.dff_gen[1].d2.D , \mchip.aa.accmulate.dff_gen[0].d2.D };
	assign \mchip.aa.adder.S1.S0.a  = {\mchip.aa.i0.dff_gen[7].d2.Q , \mchip.aa.i0.dff_gen[6].d2.Q , \mchip.aa.i0.dff_gen[5].d2.Q , \mchip.aa.i0.dff_gen[4].d2.Q };
	assign \mchip.aa.adder.S1.S0.b  = {\mchip.aa.accmulate.dff_gen[7].d2.Q , \mchip.aa.accmulate.dff_gen[6].d2.Q , \mchip.aa.accmulate.dff_gen[5].d2.Q , \mchip.aa.accmulate.dff_gen[4].d2.Q };
	assign \mchip.aa.adder.S1.S0.carry_in  = 1'h0;
	assign \mchip.aa.adder.S1.S0.fa0.a  = \mchip.aa.i0.dff_gen[4].d2.Q ;
	assign \mchip.aa.adder.S1.S0.fa0.b  = \mchip.aa.accmulate.dff_gen[4].d2.Q ;
	assign \mchip.aa.adder.S1.S0.fa0.carry_in  = 1'h0;
	assign \mchip.aa.adder.S1.S0.fa0.w3  = 1'h0;
	assign \mchip.aa.adder.S1.S0.fa1.a  = \mchip.aa.i0.dff_gen[5].d2.Q ;
	assign \mchip.aa.adder.S1.S0.fa1.b  = \mchip.aa.accmulate.dff_gen[5].d2.Q ;
	assign \mchip.aa.adder.S1.S0.fa2.a  = \mchip.aa.i0.dff_gen[6].d2.Q ;
	assign \mchip.aa.adder.S1.S0.fa2.b  = \mchip.aa.accmulate.dff_gen[6].d2.Q ;
	assign \mchip.aa.adder.S1.S0.fa3.a  = \mchip.aa.i0.dff_gen[7].d2.Q ;
	assign \mchip.aa.adder.S1.S0.fa3.b  = \mchip.aa.accmulate.dff_gen[7].d2.Q ;
	assign \mchip.aa.adder.S1.S0.sum  = 4'h0;
	assign \mchip.aa.adder.S1.S1.a  = {\mchip.aa.i0.dff_gen[7].d2.Q , \mchip.aa.i0.dff_gen[6].d2.Q , \mchip.aa.i0.dff_gen[5].d2.Q , \mchip.aa.i0.dff_gen[4].d2.Q };
	assign \mchip.aa.adder.S1.S1.b  = {\mchip.aa.accmulate.dff_gen[7].d2.Q , \mchip.aa.accmulate.dff_gen[6].d2.Q , \mchip.aa.accmulate.dff_gen[5].d2.Q , \mchip.aa.accmulate.dff_gen[4].d2.Q };
	assign \mchip.aa.adder.S1.S1.carry_in  = 1'h1;
	assign \mchip.aa.adder.S1.S1.fa0.a  = \mchip.aa.i0.dff_gen[4].d2.Q ;
	assign \mchip.aa.adder.S1.S1.fa0.b  = \mchip.aa.accmulate.dff_gen[4].d2.Q ;
	assign \mchip.aa.adder.S1.S1.fa0.carry_in  = 1'h1;
	assign \mchip.aa.adder.S1.S1.fa1.a  = \mchip.aa.i0.dff_gen[5].d2.Q ;
	assign \mchip.aa.adder.S1.S1.fa1.b  = \mchip.aa.accmulate.dff_gen[5].d2.Q ;
	assign \mchip.aa.adder.S1.S1.fa2.a  = \mchip.aa.i0.dff_gen[6].d2.Q ;
	assign \mchip.aa.adder.S1.S1.fa2.b  = \mchip.aa.accmulate.dff_gen[6].d2.Q ;
	assign \mchip.aa.adder.S1.S1.fa3.a  = \mchip.aa.i0.dff_gen[7].d2.Q ;
	assign \mchip.aa.adder.S1.S1.fa3.b  = \mchip.aa.accmulate.dff_gen[7].d2.Q ;
	assign \mchip.aa.adder.S1.S1.sum  = 4'h0;
	assign \mchip.aa.adder.S1.SUM0  = 4'h0;
	assign \mchip.aa.adder.S1.SUM1  = 4'h0;
	assign \mchip.aa.adder.S1.a  = {\mchip.aa.i0.dff_gen[7].d2.Q , \mchip.aa.i0.dff_gen[6].d2.Q , \mchip.aa.i0.dff_gen[5].d2.Q , \mchip.aa.i0.dff_gen[4].d2.Q };
	assign \mchip.aa.adder.S1.b  = {\mchip.aa.accmulate.dff_gen[7].d2.Q , \mchip.aa.accmulate.dff_gen[6].d2.Q , \mchip.aa.accmulate.dff_gen[5].d2.Q , \mchip.aa.accmulate.dff_gen[4].d2.Q };
	assign \mchip.aa.adder.S1.sum  = {\mchip.aa.accmulate.dff_gen[7].d2.D , \mchip.aa.accmulate.dff_gen[6].d2.D , \mchip.aa.accmulate.dff_gen[5].d2.D , \mchip.aa.accmulate.dff_gen[4].d2.D };
	assign \mchip.aa.adder.S2.S0.a  = {\mchip.aa.i0.dff_gen[11].d2.Q , \mchip.aa.i0.dff_gen[10].d2.Q , \mchip.aa.i0.dff_gen[9].d2.Q , \mchip.aa.i0.dff_gen[8].d2.Q };
	assign \mchip.aa.adder.S2.S0.b  = {\mchip.aa.accmulate.dff_gen[11].d2.Q , \mchip.aa.accmulate.dff_gen[10].d2.Q , \mchip.aa.accmulate.dff_gen[9].d2.Q , \mchip.aa.accmulate.dff_gen[8].d2.Q };
	assign \mchip.aa.adder.S2.S0.carry_in  = 1'h0;
	assign \mchip.aa.adder.S2.S0.fa0.a  = \mchip.aa.i0.dff_gen[8].d2.Q ;
	assign \mchip.aa.adder.S2.S0.fa0.b  = \mchip.aa.accmulate.dff_gen[8].d2.Q ;
	assign \mchip.aa.adder.S2.S0.fa0.carry_in  = 1'h0;
	assign \mchip.aa.adder.S2.S0.fa0.w3  = 1'h0;
	assign \mchip.aa.adder.S2.S0.fa1.a  = \mchip.aa.i0.dff_gen[9].d2.Q ;
	assign \mchip.aa.adder.S2.S0.fa1.b  = \mchip.aa.accmulate.dff_gen[9].d2.Q ;
	assign \mchip.aa.adder.S2.S0.fa2.a  = \mchip.aa.i0.dff_gen[10].d2.Q ;
	assign \mchip.aa.adder.S2.S0.fa2.b  = \mchip.aa.accmulate.dff_gen[10].d2.Q ;
	assign \mchip.aa.adder.S2.S0.fa3.a  = \mchip.aa.i0.dff_gen[11].d2.Q ;
	assign \mchip.aa.adder.S2.S0.fa3.b  = \mchip.aa.accmulate.dff_gen[11].d2.Q ;
	assign \mchip.aa.adder.S2.S0.sum  = 4'h0;
	assign \mchip.aa.adder.S2.S1.a  = {\mchip.aa.i0.dff_gen[11].d2.Q , \mchip.aa.i0.dff_gen[10].d2.Q , \mchip.aa.i0.dff_gen[9].d2.Q , \mchip.aa.i0.dff_gen[8].d2.Q };
	assign \mchip.aa.adder.S2.S1.b  = {\mchip.aa.accmulate.dff_gen[11].d2.Q , \mchip.aa.accmulate.dff_gen[10].d2.Q , \mchip.aa.accmulate.dff_gen[9].d2.Q , \mchip.aa.accmulate.dff_gen[8].d2.Q };
	assign \mchip.aa.adder.S2.S1.carry_in  = 1'h1;
	assign \mchip.aa.adder.S2.S1.fa0.a  = \mchip.aa.i0.dff_gen[8].d2.Q ;
	assign \mchip.aa.adder.S2.S1.fa0.b  = \mchip.aa.accmulate.dff_gen[8].d2.Q ;
	assign \mchip.aa.adder.S2.S1.fa0.carry_in  = 1'h1;
	assign \mchip.aa.adder.S2.S1.fa1.a  = \mchip.aa.i0.dff_gen[9].d2.Q ;
	assign \mchip.aa.adder.S2.S1.fa1.b  = \mchip.aa.accmulate.dff_gen[9].d2.Q ;
	assign \mchip.aa.adder.S2.S1.fa2.a  = \mchip.aa.i0.dff_gen[10].d2.Q ;
	assign \mchip.aa.adder.S2.S1.fa2.b  = \mchip.aa.accmulate.dff_gen[10].d2.Q ;
	assign \mchip.aa.adder.S2.S1.fa3.a  = \mchip.aa.i0.dff_gen[11].d2.Q ;
	assign \mchip.aa.adder.S2.S1.fa3.b  = \mchip.aa.accmulate.dff_gen[11].d2.Q ;
	assign \mchip.aa.adder.S2.S1.sum  = 4'h0;
	assign \mchip.aa.adder.S2.SUM0  = 4'h0;
	assign \mchip.aa.adder.S2.SUM1  = 4'h0;
	assign \mchip.aa.adder.S2.a  = {\mchip.aa.i0.dff_gen[11].d2.Q , \mchip.aa.i0.dff_gen[10].d2.Q , \mchip.aa.i0.dff_gen[9].d2.Q , \mchip.aa.i0.dff_gen[8].d2.Q };
	assign \mchip.aa.adder.S2.b  = {\mchip.aa.accmulate.dff_gen[11].d2.Q , \mchip.aa.accmulate.dff_gen[10].d2.Q , \mchip.aa.accmulate.dff_gen[9].d2.Q , \mchip.aa.accmulate.dff_gen[8].d2.Q };
	assign \mchip.aa.adder.S2.sum  = {\mchip.aa.accmulate.dff_gen[11].d2.D , \mchip.aa.accmulate.dff_gen[10].d2.D , \mchip.aa.accmulate.dff_gen[9].d2.D , \mchip.aa.accmulate.dff_gen[8].d2.D };
	assign \mchip.aa.adder.S3.S0.a  = {\mchip.aa.i0.dff_gen[15].d2.Q , \mchip.aa.i0.dff_gen[14].d2.Q , \mchip.aa.i0.dff_gen[13].d2.Q , \mchip.aa.i0.dff_gen[12].d2.Q };
	assign \mchip.aa.adder.S3.S0.b  = {\mchip.aa.accmulate.dff_gen[15].d2.Q , \mchip.aa.accmulate.dff_gen[14].d2.Q , \mchip.aa.accmulate.dff_gen[13].d2.Q , \mchip.aa.accmulate.dff_gen[12].d2.Q };
	assign \mchip.aa.adder.S3.S0.carry_in  = 1'h0;
	assign \mchip.aa.adder.S3.S0.fa0.a  = \mchip.aa.i0.dff_gen[12].d2.Q ;
	assign \mchip.aa.adder.S3.S0.fa0.b  = \mchip.aa.accmulate.dff_gen[12].d2.Q ;
	assign \mchip.aa.adder.S3.S0.fa0.carry_in  = 1'h0;
	assign \mchip.aa.adder.S3.S0.fa0.w3  = 1'h0;
	assign \mchip.aa.adder.S3.S0.fa1.a  = \mchip.aa.i0.dff_gen[13].d2.Q ;
	assign \mchip.aa.adder.S3.S0.fa1.b  = \mchip.aa.accmulate.dff_gen[13].d2.Q ;
	assign \mchip.aa.adder.S3.S0.fa2.a  = \mchip.aa.i0.dff_gen[14].d2.Q ;
	assign \mchip.aa.adder.S3.S0.fa2.b  = \mchip.aa.accmulate.dff_gen[14].d2.Q ;
	assign \mchip.aa.adder.S3.S0.fa3.a  = \mchip.aa.i0.dff_gen[15].d2.Q ;
	assign \mchip.aa.adder.S3.S0.fa3.b  = \mchip.aa.accmulate.dff_gen[15].d2.Q ;
	assign \mchip.aa.adder.S3.S0.sum  = 4'h0;
	assign \mchip.aa.adder.S3.S1.a  = {\mchip.aa.i0.dff_gen[15].d2.Q , \mchip.aa.i0.dff_gen[14].d2.Q , \mchip.aa.i0.dff_gen[13].d2.Q , \mchip.aa.i0.dff_gen[12].d2.Q };
	assign \mchip.aa.adder.S3.S1.b  = {\mchip.aa.accmulate.dff_gen[15].d2.Q , \mchip.aa.accmulate.dff_gen[14].d2.Q , \mchip.aa.accmulate.dff_gen[13].d2.Q , \mchip.aa.accmulate.dff_gen[12].d2.Q };
	assign \mchip.aa.adder.S3.S1.carry_in  = 1'h1;
	assign \mchip.aa.adder.S3.S1.fa0.a  = \mchip.aa.i0.dff_gen[12].d2.Q ;
	assign \mchip.aa.adder.S3.S1.fa0.b  = \mchip.aa.accmulate.dff_gen[12].d2.Q ;
	assign \mchip.aa.adder.S3.S1.fa0.carry_in  = 1'h1;
	assign \mchip.aa.adder.S3.S1.fa1.a  = \mchip.aa.i0.dff_gen[13].d2.Q ;
	assign \mchip.aa.adder.S3.S1.fa1.b  = \mchip.aa.accmulate.dff_gen[13].d2.Q ;
	assign \mchip.aa.adder.S3.S1.fa2.a  = \mchip.aa.i0.dff_gen[14].d2.Q ;
	assign \mchip.aa.adder.S3.S1.fa2.b  = \mchip.aa.accmulate.dff_gen[14].d2.Q ;
	assign \mchip.aa.adder.S3.S1.fa3.a  = \mchip.aa.i0.dff_gen[15].d2.Q ;
	assign \mchip.aa.adder.S3.S1.fa3.b  = \mchip.aa.accmulate.dff_gen[15].d2.Q ;
	assign \mchip.aa.adder.S3.S1.sum  = 4'h0;
	assign \mchip.aa.adder.S3.SUM0  = 4'h0;
	assign \mchip.aa.adder.S3.SUM1  = 4'h0;
	assign \mchip.aa.adder.S3.a  = {\mchip.aa.i0.dff_gen[15].d2.Q , \mchip.aa.i0.dff_gen[14].d2.Q , \mchip.aa.i0.dff_gen[13].d2.Q , \mchip.aa.i0.dff_gen[12].d2.Q };
	assign \mchip.aa.adder.S3.b  = {\mchip.aa.accmulate.dff_gen[15].d2.Q , \mchip.aa.accmulate.dff_gen[14].d2.Q , \mchip.aa.accmulate.dff_gen[13].d2.Q , \mchip.aa.accmulate.dff_gen[12].d2.Q };
	assign \mchip.aa.adder.S3.carry_out  = \mchip.aa.adder.S4.carry_in ;
	assign \mchip.aa.adder.S3.sum  = {\mchip.aa.accmulate.dff_gen[15].d2.D , \mchip.aa.accmulate.dff_gen[14].d2.D , \mchip.aa.accmulate.dff_gen[13].d2.D , \mchip.aa.accmulate.dff_gen[12].d2.D };
	assign \mchip.aa.adder.S4.S0.a  = 4'h0;
	assign \mchip.aa.adder.S4.S0.b  = {\mchip.aa.accmulate.dff_gen[19].d2.Q , \mchip.aa.accmulate.dff_gen[18].d2.Q , \mchip.aa.accmulate.dff_gen[17].d2.Q , \mchip.aa.accmulate.dff_gen[16].d2.Q };
	assign \mchip.aa.adder.S4.S0.carry_in  = 1'h0;
	assign \mchip.aa.adder.S4.S0.carry_out  = 1'h0;
	assign \mchip.aa.adder.S4.S0.fa0.a  = 1'h0;
	assign \mchip.aa.adder.S4.S0.fa0.b  = \mchip.aa.accmulate.dff_gen[16].d2.Q ;
	assign \mchip.aa.adder.S4.S0.fa0.carry_in  = 1'h0;
	assign \mchip.aa.adder.S4.S0.fa0.carry_out  = 1'h0;
	assign \mchip.aa.adder.S4.S0.fa0.sum  = \mchip.aa.accmulate.dff_gen[16].d2.Q ;
	assign \mchip.aa.adder.S4.S0.fa0.w1  = \mchip.aa.accmulate.dff_gen[16].d2.Q ;
	assign \mchip.aa.adder.S4.S0.fa0.w2  = 1'h0;
	assign \mchip.aa.adder.S4.S0.fa0.w3  = 1'h0;
	assign \mchip.aa.adder.S4.S0.fa1.a  = 1'h0;
	assign \mchip.aa.adder.S4.S0.fa1.b  = \mchip.aa.accmulate.dff_gen[17].d2.Q ;
	assign \mchip.aa.adder.S4.S0.fa1.carry_in  = 1'h0;
	assign \mchip.aa.adder.S4.S0.fa1.carry_out  = 1'h0;
	assign \mchip.aa.adder.S4.S0.fa1.sum  = \mchip.aa.accmulate.dff_gen[17].d2.Q ;
	assign \mchip.aa.adder.S4.S0.fa1.w1  = \mchip.aa.accmulate.dff_gen[17].d2.Q ;
	assign \mchip.aa.adder.S4.S0.fa1.w2  = 1'h0;
	assign \mchip.aa.adder.S4.S0.fa1.w3  = 1'h0;
	assign \mchip.aa.adder.S4.S0.fa2.a  = 1'h0;
	assign \mchip.aa.adder.S4.S0.fa2.b  = \mchip.aa.accmulate.dff_gen[18].d2.Q ;
	assign \mchip.aa.adder.S4.S0.fa2.carry_in  = 1'h0;
	assign \mchip.aa.adder.S4.S0.fa2.carry_out  = 1'h0;
	assign \mchip.aa.adder.S4.S0.fa2.sum  = \mchip.aa.accmulate.dff_gen[18].d2.Q ;
	assign \mchip.aa.adder.S4.S0.fa2.w1  = \mchip.aa.accmulate.dff_gen[18].d2.Q ;
	assign \mchip.aa.adder.S4.S0.fa2.w2  = 1'h0;
	assign \mchip.aa.adder.S4.S0.fa2.w3  = 1'h0;
	assign \mchip.aa.adder.S4.S0.fa3.a  = 1'h0;
	assign \mchip.aa.adder.S4.S0.fa3.b  = \mchip.aa.accmulate.dff_gen[19].d2.Q ;
	assign \mchip.aa.adder.S4.S0.fa3.carry_in  = 1'h0;
	assign \mchip.aa.adder.S4.S0.fa3.carry_out  = 1'h0;
	assign \mchip.aa.adder.S4.S0.fa3.sum  = \mchip.aa.accmulate.dff_gen[19].d2.Q ;
	assign \mchip.aa.adder.S4.S0.fa3.w1  = \mchip.aa.accmulate.dff_gen[19].d2.Q ;
	assign \mchip.aa.adder.S4.S0.fa3.w2  = 1'h0;
	assign \mchip.aa.adder.S4.S0.fa3.w3  = 1'h0;
	assign \mchip.aa.adder.S4.S0.sum  = {\mchip.aa.accmulate.dff_gen[19].d2.Q , \mchip.aa.accmulate.dff_gen[18].d2.Q , \mchip.aa.accmulate.dff_gen[17].d2.Q , \mchip.aa.accmulate.dff_gen[16].d2.Q };
	assign \mchip.aa.adder.S4.S0.w1  = 1'h0;
	assign \mchip.aa.adder.S4.S0.w2  = 1'h0;
	assign \mchip.aa.adder.S4.S0.w3  = 1'h0;
	assign \mchip.aa.adder.S4.S1.a  = 4'h0;
	assign \mchip.aa.adder.S4.S1.b  = {\mchip.aa.accmulate.dff_gen[19].d2.Q , \mchip.aa.accmulate.dff_gen[18].d2.Q , \mchip.aa.accmulate.dff_gen[17].d2.Q , \mchip.aa.accmulate.dff_gen[16].d2.Q };
	assign \mchip.aa.adder.S4.S1.carry_in  = 1'h1;
	assign \mchip.aa.adder.S4.S1.fa0.a  = 1'h0;
	assign \mchip.aa.adder.S4.S1.fa0.b  = \mchip.aa.accmulate.dff_gen[16].d2.Q ;
	assign \mchip.aa.adder.S4.S1.fa0.carry_in  = 1'h1;
	assign \mchip.aa.adder.S4.S1.fa0.carry_out  = \mchip.aa.accmulate.dff_gen[16].d2.Q ;
	assign \mchip.aa.adder.S4.S1.fa0.w1  = \mchip.aa.accmulate.dff_gen[16].d2.Q ;
	assign \mchip.aa.adder.S4.S1.fa0.w2  = 1'h0;
	assign \mchip.aa.adder.S4.S1.fa0.w3  = \mchip.aa.accmulate.dff_gen[16].d2.Q ;
	assign \mchip.aa.adder.S4.S1.fa1.a  = 1'h0;
	assign \mchip.aa.adder.S4.S1.fa1.b  = \mchip.aa.accmulate.dff_gen[17].d2.Q ;
	assign \mchip.aa.adder.S4.S1.fa1.carry_in  = \mchip.aa.accmulate.dff_gen[16].d2.Q ;
	assign \mchip.aa.adder.S4.S1.fa1.w1  = \mchip.aa.accmulate.dff_gen[17].d2.Q ;
	assign \mchip.aa.adder.S4.S1.fa1.w2  = 1'h0;
	assign \mchip.aa.adder.S4.S1.fa2.a  = 1'h0;
	assign \mchip.aa.adder.S4.S1.fa2.b  = \mchip.aa.accmulate.dff_gen[18].d2.Q ;
	assign \mchip.aa.adder.S4.S1.fa2.w1  = \mchip.aa.accmulate.dff_gen[18].d2.Q ;
	assign \mchip.aa.adder.S4.S1.fa2.w2  = 1'h0;
	assign \mchip.aa.adder.S4.S1.fa3.a  = 1'h0;
	assign \mchip.aa.adder.S4.S1.fa3.b  = \mchip.aa.accmulate.dff_gen[19].d2.Q ;
	assign \mchip.aa.adder.S4.S1.fa3.w1  = \mchip.aa.accmulate.dff_gen[19].d2.Q ;
	assign \mchip.aa.adder.S4.S1.fa3.w2  = 1'h0;
	assign \mchip.aa.adder.S4.S1.sum  = {\mchip.aa.adder.S4.S1.fa3.sum , \mchip.aa.adder.S4.S1.fa2.sum , \mchip.aa.adder.S4.S1.fa1.sum , \mchip.aa.adder.S4.S1.fa0.sum };
	assign \mchip.aa.adder.S4.S1.w1  = \mchip.aa.accmulate.dff_gen[16].d2.Q ;
	assign \mchip.aa.adder.S4.SUM0  = {\mchip.aa.accmulate.dff_gen[19].d2.Q , \mchip.aa.accmulate.dff_gen[18].d2.Q , \mchip.aa.accmulate.dff_gen[17].d2.Q , \mchip.aa.accmulate.dff_gen[16].d2.Q };
	assign \mchip.aa.adder.S4.SUM1  = {\mchip.aa.adder.S4.S1.fa3.sum , \mchip.aa.adder.S4.S1.fa2.sum , \mchip.aa.adder.S4.S1.fa1.sum , \mchip.aa.adder.S4.S1.fa0.sum };
	assign \mchip.aa.adder.S4.a  = 4'h0;
	assign \mchip.aa.adder.S4.b  = {\mchip.aa.accmulate.dff_gen[19].d2.Q , \mchip.aa.accmulate.dff_gen[18].d2.Q , \mchip.aa.accmulate.dff_gen[17].d2.Q , \mchip.aa.accmulate.dff_gen[16].d2.Q };
	assign \mchip.aa.adder.S4.carry0  = 1'h0;
	assign \mchip.aa.adder.a  = {4'h0, \mchip.aa.i0.dff_gen[15].d2.Q , \mchip.aa.i0.dff_gen[14].d2.Q , \mchip.aa.i0.dff_gen[13].d2.Q , \mchip.aa.i0.dff_gen[12].d2.Q , \mchip.aa.i0.dff_gen[11].d2.Q , \mchip.aa.i0.dff_gen[10].d2.Q , \mchip.aa.i0.dff_gen[9].d2.Q , \mchip.aa.i0.dff_gen[8].d2.Q , \mchip.aa.i0.dff_gen[7].d2.Q , \mchip.aa.i0.dff_gen[6].d2.Q , \mchip.aa.i0.dff_gen[5].d2.Q , \mchip.aa.i0.dff_gen[4].d2.Q , \mchip.aa.i0.dff_gen[3].d2.Q , \mchip.aa.i0.dff_gen[2].d2.Q , \mchip.aa.i0.dff_gen[1].d2.Q , \mchip.aa.i0.dff_gen[0].d2.Q };
	assign \mchip.aa.adder.b  = {\mchip.aa.accmulate.dff_gen[19].d2.Q , \mchip.aa.accmulate.dff_gen[18].d2.Q , \mchip.aa.accmulate.dff_gen[17].d2.Q , \mchip.aa.accmulate.dff_gen[16].d2.Q , \mchip.aa.accmulate.dff_gen[15].d2.Q , \mchip.aa.accmulate.dff_gen[14].d2.Q , \mchip.aa.accmulate.dff_gen[13].d2.Q , \mchip.aa.accmulate.dff_gen[12].d2.Q , \mchip.aa.accmulate.dff_gen[11].d2.Q , \mchip.aa.accmulate.dff_gen[10].d2.Q , \mchip.aa.accmulate.dff_gen[9].d2.Q , \mchip.aa.accmulate.dff_gen[8].d2.Q , \mchip.aa.accmulate.dff_gen[7].d2.Q , \mchip.aa.accmulate.dff_gen[6].d2.Q , \mchip.aa.accmulate.dff_gen[5].d2.Q , \mchip.aa.accmulate.dff_gen[4].d2.Q , \mchip.aa.accmulate.dff_gen[3].d2.Q , \mchip.aa.accmulate.dff_gen[2].d2.Q , \mchip.aa.accmulate.dff_gen[1].d2.Q , \mchip.aa.accmulate.dff_gen[0].d2.Q };
	assign \mchip.aa.adder.carry_in  = 1'h0;
	assign \mchip.aa.adder.carry_out  = \mchip.aa.adder.S4.carry_out ;
	assign \mchip.aa.adder.sum  = {4'h0, \mchip.aa.accmulate.dff_gen[15].d2.D , \mchip.aa.accmulate.dff_gen[14].d2.D , \mchip.aa.accmulate.dff_gen[13].d2.D , \mchip.aa.accmulate.dff_gen[12].d2.D , \mchip.aa.accmulate.dff_gen[11].d2.D , \mchip.aa.accmulate.dff_gen[10].d2.D , \mchip.aa.accmulate.dff_gen[9].d2.D , \mchip.aa.accmulate.dff_gen[8].d2.D , \mchip.aa.accmulate.dff_gen[7].d2.D , \mchip.aa.accmulate.dff_gen[6].d2.D , \mchip.aa.accmulate.dff_gen[5].d2.D , \mchip.aa.accmulate.dff_gen[4].d2.D , \mchip.aa.accmulate.dff_gen[3].d2.D , \mchip.aa.accmulate.dff_gen[2].d2.D , \mchip.aa.accmulate.dff_gen[1].d2.D , \mchip.aa.accmulate.dff_gen[0].d2.D };
	assign \mchip.aa.adder.temp_carry4  = \mchip.aa.adder.S4.carry_in ;
	assign \mchip.aa.i0.add  = \mchip.control.state [5];
	assign \mchip.aa.i0.dff_gen[0].d2.D  = \mchip.mult.i3.temp_register [0];
	assign \mchip.aa.i0.dff_gen[0].d2.clk  = \mchip.control.state [5];
	assign \mchip.aa.i0.dff_gen[10].d2.D  = \mchip.mult.i3.temp_register [10];
	assign \mchip.aa.i0.dff_gen[10].d2.clk  = \mchip.control.state [5];
	assign \mchip.aa.i0.dff_gen[11].d2.D  = \mchip.mult.i3.temp_register [11];
	assign \mchip.aa.i0.dff_gen[11].d2.clk  = \mchip.control.state [5];
	assign \mchip.aa.i0.dff_gen[12].d2.D  = \mchip.mult.i3.temp_register [12];
	assign \mchip.aa.i0.dff_gen[12].d2.clk  = \mchip.control.state [5];
	assign \mchip.aa.i0.dff_gen[13].d2.D  = \mchip.mult.i3.temp_register [13];
	assign \mchip.aa.i0.dff_gen[13].d2.clk  = \mchip.control.state [5];
	assign \mchip.aa.i0.dff_gen[14].d2.D  = \mchip.mult.i3.temp_register [14];
	assign \mchip.aa.i0.dff_gen[14].d2.clk  = \mchip.control.state [5];
	assign \mchip.aa.i0.dff_gen[15].d2.D  = \mchip.mult.i3.temp_register [15];
	assign \mchip.aa.i0.dff_gen[15].d2.clk  = \mchip.control.state [5];
	assign \mchip.aa.i0.dff_gen[16].d2.D  = 1'h0;
	assign \mchip.aa.i0.dff_gen[16].d2.Q  = 1'h0;
	assign \mchip.aa.i0.dff_gen[16].d2.clk  = \mchip.control.state [5];
	assign \mchip.aa.i0.dff_gen[17].d2.D  = 1'h0;
	assign \mchip.aa.i0.dff_gen[17].d2.Q  = 1'h0;
	assign \mchip.aa.i0.dff_gen[17].d2.clk  = \mchip.control.state [5];
	assign \mchip.aa.i0.dff_gen[18].d2.D  = 1'h0;
	assign \mchip.aa.i0.dff_gen[18].d2.Q  = 1'h0;
	assign \mchip.aa.i0.dff_gen[18].d2.clk  = \mchip.control.state [5];
	assign \mchip.aa.i0.dff_gen[19].d2.D  = 1'h0;
	assign \mchip.aa.i0.dff_gen[19].d2.Q  = 1'h0;
	assign \mchip.aa.i0.dff_gen[19].d2.clk  = \mchip.control.state [5];
	assign \mchip.aa.i0.dff_gen[1].d2.D  = \mchip.mult.i3.temp_register [1];
	assign \mchip.aa.i0.dff_gen[1].d2.clk  = \mchip.control.state [5];
	assign \mchip.aa.i0.dff_gen[2].d2.D  = \mchip.mult.i3.temp_register [2];
	assign \mchip.aa.i0.dff_gen[2].d2.clk  = \mchip.control.state [5];
	assign \mchip.aa.i0.dff_gen[3].d2.D  = \mchip.mult.i3.temp_register [3];
	assign \mchip.aa.i0.dff_gen[3].d2.clk  = \mchip.control.state [5];
	assign \mchip.aa.i0.dff_gen[4].d2.D  = \mchip.mult.i3.temp_register [4];
	assign \mchip.aa.i0.dff_gen[4].d2.clk  = \mchip.control.state [5];
	assign \mchip.aa.i0.dff_gen[5].d2.D  = \mchip.mult.i3.temp_register [5];
	assign \mchip.aa.i0.dff_gen[5].d2.clk  = \mchip.control.state [5];
	assign \mchip.aa.i0.dff_gen[6].d2.D  = \mchip.mult.i3.temp_register [6];
	assign \mchip.aa.i0.dff_gen[6].d2.clk  = \mchip.control.state [5];
	assign \mchip.aa.i0.dff_gen[7].d2.D  = \mchip.mult.i3.temp_register [7];
	assign \mchip.aa.i0.dff_gen[7].d2.clk  = \mchip.control.state [5];
	assign \mchip.aa.i0.dff_gen[8].d2.D  = \mchip.mult.i3.temp_register [8];
	assign \mchip.aa.i0.dff_gen[8].d2.clk  = \mchip.control.state [5];
	assign \mchip.aa.i0.dff_gen[9].d2.D  = \mchip.mult.i3.temp_register [9];
	assign \mchip.aa.i0.dff_gen[9].d2.clk  = \mchip.control.state [5];
	assign \mchip.aa.i0.in  = {4'h0, \mchip.mult.i3.temp_register [15:0]};
	assign \mchip.aa.i0.out  = {4'h0, \mchip.aa.i0.dff_gen[15].d2.Q , \mchip.aa.i0.dff_gen[14].d2.Q , \mchip.aa.i0.dff_gen[13].d2.Q , \mchip.aa.i0.dff_gen[12].d2.Q , \mchip.aa.i0.dff_gen[11].d2.Q , \mchip.aa.i0.dff_gen[10].d2.Q , \mchip.aa.i0.dff_gen[9].d2.Q , \mchip.aa.i0.dff_gen[8].d2.Q , \mchip.aa.i0.dff_gen[7].d2.Q , \mchip.aa.i0.dff_gen[6].d2.Q , \mchip.aa.i0.dff_gen[5].d2.Q , \mchip.aa.i0.dff_gen[4].d2.Q , \mchip.aa.i0.dff_gen[3].d2.Q , \mchip.aa.i0.dff_gen[2].d2.Q , \mchip.aa.i0.dff_gen[1].d2.Q , \mchip.aa.i0.dff_gen[0].d2.Q };
	assign \mchip.aa.i0.temp_out  = {4'h0, \mchip.aa.i0.dff_gen[15].d2.Q , \mchip.aa.i0.dff_gen[14].d2.Q , \mchip.aa.i0.dff_gen[13].d2.Q , \mchip.aa.i0.dff_gen[12].d2.Q , \mchip.aa.i0.dff_gen[11].d2.Q , \mchip.aa.i0.dff_gen[10].d2.Q , \mchip.aa.i0.dff_gen[9].d2.Q , \mchip.aa.i0.dff_gen[8].d2.Q , \mchip.aa.i0.dff_gen[7].d2.Q , \mchip.aa.i0.dff_gen[6].d2.Q , \mchip.aa.i0.dff_gen[5].d2.Q , \mchip.aa.i0.dff_gen[4].d2.Q , \mchip.aa.i0.dff_gen[3].d2.Q , \mchip.aa.i0.dff_gen[2].d2.Q , \mchip.aa.i0.dff_gen[1].d2.Q , \mchip.aa.i0.dff_gen[0].d2.Q };
	assign \mchip.aa.mult_res_in  = \mchip.mult.i3.temp_register [15:0];
	assign \mchip.aa.mult_res_out  = {4'h0, \mchip.aa.i0.dff_gen[15].d2.Q , \mchip.aa.i0.dff_gen[14].d2.Q , \mchip.aa.i0.dff_gen[13].d2.Q , \mchip.aa.i0.dff_gen[12].d2.Q , \mchip.aa.i0.dff_gen[11].d2.Q , \mchip.aa.i0.dff_gen[10].d2.Q , \mchip.aa.i0.dff_gen[9].d2.Q , \mchip.aa.i0.dff_gen[8].d2.Q , \mchip.aa.i0.dff_gen[7].d2.Q , \mchip.aa.i0.dff_gen[6].d2.Q , \mchip.aa.i0.dff_gen[5].d2.Q , \mchip.aa.i0.dff_gen[4].d2.Q , \mchip.aa.i0.dff_gen[3].d2.Q , \mchip.aa.i0.dff_gen[2].d2.Q , \mchip.aa.i0.dff_gen[1].d2.Q , \mchip.aa.i0.dff_gen[0].d2.Q };
	assign \mchip.aa.result  = {\mchip.aa.accmulate.dff_gen[19].d2.Q , \mchip.aa.accmulate.dff_gen[18].d2.Q , \mchip.aa.accmulate.dff_gen[17].d2.Q , \mchip.aa.accmulate.dff_gen[16].d2.Q , \mchip.aa.accmulate.dff_gen[15].d2.Q , \mchip.aa.accmulate.dff_gen[14].d2.Q , \mchip.aa.accmulate.dff_gen[13].d2.Q , \mchip.aa.accmulate.dff_gen[12].d2.Q , \mchip.aa.accmulate.dff_gen[11].d2.Q , \mchip.aa.accmulate.dff_gen[10].d2.Q , \mchip.aa.accmulate.dff_gen[9].d2.Q , \mchip.aa.accmulate.dff_gen[8].d2.Q , \mchip.aa.accmulate.dff_gen[7].d2.Q , \mchip.aa.accmulate.dff_gen[6].d2.Q , \mchip.aa.accmulate.dff_gen[5].d2.Q , \mchip.aa.accmulate.dff_gen[4].d2.Q , \mchip.aa.accmulate.dff_gen[3].d2.Q , \mchip.aa.accmulate.dff_gen[2].d2.Q , \mchip.aa.accmulate.dff_gen[1].d2.Q , \mchip.aa.accmulate.dff_gen[0].d2.Q };
	assign \mchip.aa.result_carry_out  = \mchip.aa.adder.S4.carry_out ;
	assign \mchip.aa.temp_mult_res_in  = {4'h0, \mchip.mult.i3.temp_register [15:0]};
	assign \mchip.aa.temp_result  = {\mchip.aa.accmulate.dff_gen[19].d2.Q , \mchip.aa.accmulate.dff_gen[18].d2.Q , \mchip.aa.accmulate.dff_gen[17].d2.Q , \mchip.aa.accmulate.dff_gen[16].d2.Q , \mchip.aa.accmulate.dff_gen[15].d2.Q , \mchip.aa.accmulate.dff_gen[14].d2.Q , \mchip.aa.accmulate.dff_gen[13].d2.Q , \mchip.aa.accmulate.dff_gen[12].d2.Q , \mchip.aa.accmulate.dff_gen[11].d2.Q , \mchip.aa.accmulate.dff_gen[10].d2.Q , \mchip.aa.accmulate.dff_gen[9].d2.Q , \mchip.aa.accmulate.dff_gen[8].d2.Q , \mchip.aa.accmulate.dff_gen[7].d2.Q , \mchip.aa.accmulate.dff_gen[6].d2.Q , \mchip.aa.accmulate.dff_gen[5].d2.Q , \mchip.aa.accmulate.dff_gen[4].d2.Q , \mchip.aa.accmulate.dff_gen[3].d2.Q , \mchip.aa.accmulate.dff_gen[2].d2.Q , \mchip.aa.accmulate.dff_gen[1].d2.Q , \mchip.aa.accmulate.dff_gen[0].d2.Q };
	assign \mchip.add  = \mchip.control.state [5];
	assign \mchip.clock  = io_in[12];
	assign \mchip.control.Begin_mul  = \mchip.control.state [6];
	assign \mchip.control.End_mul  = \mchip.mult.i0.state [0];
	assign \mchip.control.Finish  = \mchip.control.state [0];
	assign \mchip.control.Load_op  = \mchip.control.state [2];
	assign \mchip.control.START  = io_in[11];
	assign \mchip.control.add  = \mchip.control.state [5];
	assign \mchip.control.clk  = io_in[12];
	assign \mchip.control.do_next  = io_in[7];
	assign \mchip.do_next  = io_in[7];
	assign \mchip.io_in  = io_in[11:0];
	assign \mchip.io_out  = {\mchip.aa.adder.S4.carry_out , \mchip.control.state [0], \mchip.shiftout [0], \mchip.mult.i0.state [0], 8'h00};
	assign \mchip.mac_carry_out  = \mchip.aa.adder.S4.carry_out ;
	assign \mchip.mac_res  = {\mchip.aa.accmulate.dff_gen[19].d2.Q , \mchip.aa.accmulate.dff_gen[18].d2.Q , \mchip.aa.accmulate.dff_gen[17].d2.Q , \mchip.aa.accmulate.dff_gen[16].d2.Q , \mchip.aa.accmulate.dff_gen[15].d2.Q , \mchip.aa.accmulate.dff_gen[14].d2.Q , \mchip.aa.accmulate.dff_gen[13].d2.Q , \mchip.aa.accmulate.dff_gen[12].d2.Q , \mchip.aa.accmulate.dff_gen[11].d2.Q , \mchip.aa.accmulate.dff_gen[10].d2.Q , \mchip.aa.accmulate.dff_gen[9].d2.Q , \mchip.aa.accmulate.dff_gen[8].d2.Q , \mchip.aa.accmulate.dff_gen[7].d2.Q , \mchip.aa.accmulate.dff_gen[6].d2.Q , \mchip.aa.accmulate.dff_gen[5].d2.Q , \mchip.aa.accmulate.dff_gen[4].d2.Q , \mchip.aa.accmulate.dff_gen[3].d2.Q , \mchip.aa.accmulate.dff_gen[2].d2.Q , \mchip.aa.accmulate.dff_gen[1].d2.Q , \mchip.aa.accmulate.dff_gen[0].d2.Q };
	assign \mchip.mult.Begin_mul  = \mchip.control.state [6];
	assign \mchip.mult.End_mul  = \mchip.mult.i0.state [0];
	assign \mchip.mult.LSB  = \mchip.mult.i3.temp_register [0];
	assign \mchip.mult.Load_mul  = \mchip.mult.i0.state [3];
	assign \mchip.mult.a_in  = {\mchip.opa.dff_gen[7].d1.Q , \mchip.opa.dff_gen[6].d1.Q , \mchip.opa.dff_gen[5].d1.Q , \mchip.opa.dff_gen[4].d1.Q , \mchip.opa.dff_gen[3].d1.Q , \mchip.opa.dff_gen[2].d1.Q , \mchip.opa.dff_gen[1].d1.Q , \mchip.opa.dff_gen[0].d1.Q };
	assign \mchip.mult.a_out  = {\mchip.mult.i1.r1.dff_gen[7].d1.Q , \mchip.mult.i1.r1.dff_gen[6].d1.Q , \mchip.mult.i1.r1.dff_gen[5].d1.Q , \mchip.mult.i1.r1.dff_gen[4].d1.Q , \mchip.mult.i1.r1.dff_gen[3].d1.Q , \mchip.mult.i1.r1.dff_gen[2].d1.Q , \mchip.mult.i1.r1.dff_gen[1].d1.Q , \mchip.mult.i1.r1.dff_gen[0].d1.Q };
	assign \mchip.mult.b_in  = {\mchip.opb.dff_gen[7].d1.Q , \mchip.opb.dff_gen[6].d1.Q , \mchip.opb.dff_gen[5].d1.Q , \mchip.opb.dff_gen[4].d1.Q , \mchip.opb.dff_gen[3].d1.Q , \mchip.opb.dff_gen[2].d1.Q , \mchip.opb.dff_gen[1].d1.Q , \mchip.opb.dff_gen[0].d1.Q };
	assign \mchip.mult.b_out  = \mchip.mult.i3.temp_register [15:8];
	assign \mchip.mult.clk  = io_in[12];
	assign \mchip.mult.do_add  = \mchip.mult.i0.state [4];
	assign \mchip.mult.do_shift  = \mchip.mult.i0.state [1];
	assign \mchip.mult.i0.Begin_mul  = \mchip.control.state [6];
	assign \mchip.mult.i0.End_mul  = \mchip.mult.i0.state [0];
	assign \mchip.mult.i0.LSB  = \mchip.mult.i3.temp_register [0];
	assign \mchip.mult.i0.Load_mul  = \mchip.mult.i0.state [3];
	assign \mchip.mult.i0.clk  = io_in[12];
	assign \mchip.mult.i0.do_add  = \mchip.mult.i0.state [4];
	assign \mchip.mult.i0.do_shift  = \mchip.mult.i0.state [1];
	assign \mchip.mult.i1.Load_mul  = \mchip.mult.i0.state [3];
	assign \mchip.mult.i1.a_in  = {\mchip.opa.dff_gen[7].d1.Q , \mchip.opa.dff_gen[6].d1.Q , \mchip.opa.dff_gen[5].d1.Q , \mchip.opa.dff_gen[4].d1.Q , \mchip.opa.dff_gen[3].d1.Q , \mchip.opa.dff_gen[2].d1.Q , \mchip.opa.dff_gen[1].d1.Q , \mchip.opa.dff_gen[0].d1.Q };
	assign \mchip.mult.i1.a_out  = {\mchip.mult.i1.r1.dff_gen[7].d1.Q , \mchip.mult.i1.r1.dff_gen[6].d1.Q , \mchip.mult.i1.r1.dff_gen[5].d1.Q , \mchip.mult.i1.r1.dff_gen[4].d1.Q , \mchip.mult.i1.r1.dff_gen[3].d1.Q , \mchip.mult.i1.r1.dff_gen[2].d1.Q , \mchip.mult.i1.r1.dff_gen[1].d1.Q , \mchip.mult.i1.r1.dff_gen[0].d1.Q };
	assign \mchip.mult.i1.r1.Load_op  = \mchip.mult.i0.state [3];
	assign \mchip.mult.i1.r1.dff_gen[0].d1.D  = \mchip.opa.dff_gen[0].d1.Q ;
	assign \mchip.mult.i1.r1.dff_gen[0].d1.clk  = \mchip.mult.i0.state [3];
	assign \mchip.mult.i1.r1.dff_gen[1].d1.D  = \mchip.opa.dff_gen[1].d1.Q ;
	assign \mchip.mult.i1.r1.dff_gen[1].d1.clk  = \mchip.mult.i0.state [3];
	assign \mchip.mult.i1.r1.dff_gen[2].d1.D  = \mchip.opa.dff_gen[2].d1.Q ;
	assign \mchip.mult.i1.r1.dff_gen[2].d1.clk  = \mchip.mult.i0.state [3];
	assign \mchip.mult.i1.r1.dff_gen[3].d1.D  = \mchip.opa.dff_gen[3].d1.Q ;
	assign \mchip.mult.i1.r1.dff_gen[3].d1.clk  = \mchip.mult.i0.state [3];
	assign \mchip.mult.i1.r1.dff_gen[4].d1.D  = \mchip.opa.dff_gen[4].d1.Q ;
	assign \mchip.mult.i1.r1.dff_gen[4].d1.clk  = \mchip.mult.i0.state [3];
	assign \mchip.mult.i1.r1.dff_gen[5].d1.D  = \mchip.opa.dff_gen[5].d1.Q ;
	assign \mchip.mult.i1.r1.dff_gen[5].d1.clk  = \mchip.mult.i0.state [3];
	assign \mchip.mult.i1.r1.dff_gen[6].d1.D  = \mchip.opa.dff_gen[6].d1.Q ;
	assign \mchip.mult.i1.r1.dff_gen[6].d1.clk  = \mchip.mult.i0.state [3];
	assign \mchip.mult.i1.r1.dff_gen[7].d1.D  = \mchip.opa.dff_gen[7].d1.Q ;
	assign \mchip.mult.i1.r1.dff_gen[7].d1.clk  = \mchip.mult.i0.state [3];
	assign \mchip.mult.i1.r1.in  = {\mchip.opa.dff_gen[7].d1.Q , \mchip.opa.dff_gen[6].d1.Q , \mchip.opa.dff_gen[5].d1.Q , \mchip.opa.dff_gen[4].d1.Q , \mchip.opa.dff_gen[3].d1.Q , \mchip.opa.dff_gen[2].d1.Q , \mchip.opa.dff_gen[1].d1.Q , \mchip.opa.dff_gen[0].d1.Q };
	assign \mchip.mult.i1.r1.out  = {\mchip.mult.i1.r1.dff_gen[7].d1.Q , \mchip.mult.i1.r1.dff_gen[6].d1.Q , \mchip.mult.i1.r1.dff_gen[5].d1.Q , \mchip.mult.i1.r1.dff_gen[4].d1.Q , \mchip.mult.i1.r1.dff_gen[3].d1.Q , \mchip.mult.i1.r1.dff_gen[2].d1.Q , \mchip.mult.i1.r1.dff_gen[1].d1.Q , \mchip.mult.i1.r1.dff_gen[0].d1.Q };
	assign \mchip.mult.i1.r1.temp_out  = {\mchip.mult.i1.r1.dff_gen[7].d1.Q , \mchip.mult.i1.r1.dff_gen[6].d1.Q , \mchip.mult.i1.r1.dff_gen[5].d1.Q , \mchip.mult.i1.r1.dff_gen[4].d1.Q , \mchip.mult.i1.r1.dff_gen[3].d1.Q , \mchip.mult.i1.r1.dff_gen[2].d1.Q , \mchip.mult.i1.r1.dff_gen[1].d1.Q , \mchip.mult.i1.r1.dff_gen[0].d1.Q };
	assign \mchip.mult.i2.S0.S0.a  = {\mchip.mult.i1.r1.dff_gen[3].d1.Q , \mchip.mult.i1.r1.dff_gen[2].d1.Q , \mchip.mult.i1.r1.dff_gen[1].d1.Q , \mchip.mult.i1.r1.dff_gen[0].d1.Q };
	assign \mchip.mult.i2.S0.S0.b  = \mchip.mult.i3.temp_register [11:8];
	assign \mchip.mult.i2.S0.S0.carry_in  = 1'h0;
	assign \mchip.mult.i2.S0.S0.fa0.a  = \mchip.mult.i1.r1.dff_gen[0].d1.Q ;
	assign \mchip.mult.i2.S0.S0.fa0.b  = \mchip.mult.i3.temp_register [8];
	assign \mchip.mult.i2.S0.S0.fa0.carry_in  = 1'h0;
	assign \mchip.mult.i2.S0.S0.fa0.w3  = 1'h0;
	assign \mchip.mult.i2.S0.S0.fa1.a  = \mchip.mult.i1.r1.dff_gen[1].d1.Q ;
	assign \mchip.mult.i2.S0.S0.fa1.b  = \mchip.mult.i3.temp_register [9];
	assign \mchip.mult.i2.S0.S0.fa2.a  = \mchip.mult.i1.r1.dff_gen[2].d1.Q ;
	assign \mchip.mult.i2.S0.S0.fa2.b  = \mchip.mult.i3.temp_register [10];
	assign \mchip.mult.i2.S0.S0.fa3.a  = \mchip.mult.i1.r1.dff_gen[3].d1.Q ;
	assign \mchip.mult.i2.S0.S0.fa3.b  = \mchip.mult.i3.temp_register [11];
	assign \mchip.mult.i2.S0.S1.a  = {\mchip.mult.i1.r1.dff_gen[3].d1.Q , \mchip.mult.i1.r1.dff_gen[2].d1.Q , \mchip.mult.i1.r1.dff_gen[1].d1.Q , \mchip.mult.i1.r1.dff_gen[0].d1.Q };
	assign \mchip.mult.i2.S0.S1.b  = \mchip.mult.i3.temp_register [11:8];
	assign \mchip.mult.i2.S0.S1.carry_in  = 1'h1;
	assign \mchip.mult.i2.S0.S1.fa0.a  = \mchip.mult.i1.r1.dff_gen[0].d1.Q ;
	assign \mchip.mult.i2.S0.S1.fa0.b  = \mchip.mult.i3.temp_register [8];
	assign \mchip.mult.i2.S0.S1.fa0.carry_in  = 1'h1;
	assign \mchip.mult.i2.S0.S1.fa1.a  = \mchip.mult.i1.r1.dff_gen[1].d1.Q ;
	assign \mchip.mult.i2.S0.S1.fa1.b  = \mchip.mult.i3.temp_register [9];
	assign \mchip.mult.i2.S0.S1.fa2.a  = \mchip.mult.i1.r1.dff_gen[2].d1.Q ;
	assign \mchip.mult.i2.S0.S1.fa2.b  = \mchip.mult.i3.temp_register [10];
	assign \mchip.mult.i2.S0.S1.fa3.a  = \mchip.mult.i1.r1.dff_gen[3].d1.Q ;
	assign \mchip.mult.i2.S0.S1.fa3.b  = \mchip.mult.i3.temp_register [11];
	assign \mchip.mult.i2.S0.a  = {\mchip.mult.i1.r1.dff_gen[3].d1.Q , \mchip.mult.i1.r1.dff_gen[2].d1.Q , \mchip.mult.i1.r1.dff_gen[1].d1.Q , \mchip.mult.i1.r1.dff_gen[0].d1.Q };
	assign \mchip.mult.i2.S0.b  = \mchip.mult.i3.temp_register [11:8];
	assign \mchip.mult.i2.S0.carry_in  = 1'h0;
	assign \mchip.mult.i2.S1.S0.a  = {\mchip.mult.i1.r1.dff_gen[7].d1.Q , \mchip.mult.i1.r1.dff_gen[6].d1.Q , \mchip.mult.i1.r1.dff_gen[5].d1.Q , \mchip.mult.i1.r1.dff_gen[4].d1.Q };
	assign \mchip.mult.i2.S1.S0.b  = \mchip.mult.i3.temp_register [15:12];
	assign \mchip.mult.i2.S1.S0.carry_in  = 1'h0;
	assign \mchip.mult.i2.S1.S0.fa0.a  = \mchip.mult.i1.r1.dff_gen[4].d1.Q ;
	assign \mchip.mult.i2.S1.S0.fa0.b  = \mchip.mult.i3.temp_register [12];
	assign \mchip.mult.i2.S1.S0.fa0.carry_in  = 1'h0;
	assign \mchip.mult.i2.S1.S0.fa0.w3  = 1'h0;
	assign \mchip.mult.i2.S1.S0.fa1.a  = \mchip.mult.i1.r1.dff_gen[5].d1.Q ;
	assign \mchip.mult.i2.S1.S0.fa1.b  = \mchip.mult.i3.temp_register [13];
	assign \mchip.mult.i2.S1.S0.fa2.a  = \mchip.mult.i1.r1.dff_gen[6].d1.Q ;
	assign \mchip.mult.i2.S1.S0.fa2.b  = \mchip.mult.i3.temp_register [14];
	assign \mchip.mult.i2.S1.S0.fa3.a  = \mchip.mult.i1.r1.dff_gen[7].d1.Q ;
	assign \mchip.mult.i2.S1.S0.fa3.b  = \mchip.mult.i3.temp_register [15];
	assign \mchip.mult.i2.S1.S0.sum  = 4'h0;
	assign \mchip.mult.i2.S1.S1.a  = {\mchip.mult.i1.r1.dff_gen[7].d1.Q , \mchip.mult.i1.r1.dff_gen[6].d1.Q , \mchip.mult.i1.r1.dff_gen[5].d1.Q , \mchip.mult.i1.r1.dff_gen[4].d1.Q };
	assign \mchip.mult.i2.S1.S1.b  = \mchip.mult.i3.temp_register [15:12];
	assign \mchip.mult.i2.S1.S1.carry_in  = 1'h1;
	assign \mchip.mult.i2.S1.S1.fa0.a  = \mchip.mult.i1.r1.dff_gen[4].d1.Q ;
	assign \mchip.mult.i2.S1.S1.fa0.b  = \mchip.mult.i3.temp_register [12];
	assign \mchip.mult.i2.S1.S1.fa0.carry_in  = 1'h1;
	assign \mchip.mult.i2.S1.S1.fa1.a  = \mchip.mult.i1.r1.dff_gen[5].d1.Q ;
	assign \mchip.mult.i2.S1.S1.fa1.b  = \mchip.mult.i3.temp_register [13];
	assign \mchip.mult.i2.S1.S1.fa2.a  = \mchip.mult.i1.r1.dff_gen[6].d1.Q ;
	assign \mchip.mult.i2.S1.S1.fa2.b  = \mchip.mult.i3.temp_register [14];
	assign \mchip.mult.i2.S1.S1.fa3.a  = \mchip.mult.i1.r1.dff_gen[7].d1.Q ;
	assign \mchip.mult.i2.S1.S1.fa3.b  = \mchip.mult.i3.temp_register [15];
	assign \mchip.mult.i2.S1.S1.sum  = 4'h0;
	assign \mchip.mult.i2.S1.SUM0  = 4'h0;
	assign \mchip.mult.i2.S1.SUM1  = 4'h0;
	assign \mchip.mult.i2.S1.a  = {\mchip.mult.i1.r1.dff_gen[7].d1.Q , \mchip.mult.i1.r1.dff_gen[6].d1.Q , \mchip.mult.i1.r1.dff_gen[5].d1.Q , \mchip.mult.i1.r1.dff_gen[4].d1.Q };
	assign \mchip.mult.i2.S1.b  = \mchip.mult.i3.temp_register [15:12];
	assign \mchip.mult.i2.a  = {\mchip.mult.i1.r1.dff_gen[7].d1.Q , \mchip.mult.i1.r1.dff_gen[6].d1.Q , \mchip.mult.i1.r1.dff_gen[5].d1.Q , \mchip.mult.i1.r1.dff_gen[4].d1.Q , \mchip.mult.i1.r1.dff_gen[3].d1.Q , \mchip.mult.i1.r1.dff_gen[2].d1.Q , \mchip.mult.i1.r1.dff_gen[1].d1.Q , \mchip.mult.i1.r1.dff_gen[0].d1.Q };
	assign \mchip.mult.i2.b  = \mchip.mult.i3.temp_register [15:8];
	assign \mchip.mult.i2.carry_in  = 1'h0;
	assign \mchip.mult.i3.LSB  = \mchip.mult.i3.temp_register [0];
	assign \mchip.mult.i3.Load_mul  = \mchip.mult.i0.state [3];
	assign \mchip.mult.i3.b_in  = {\mchip.opb.dff_gen[7].d1.Q , \mchip.opb.dff_gen[6].d1.Q , \mchip.opb.dff_gen[5].d1.Q , \mchip.opb.dff_gen[4].d1.Q , \mchip.opb.dff_gen[3].d1.Q , \mchip.opb.dff_gen[2].d1.Q , \mchip.opb.dff_gen[1].d1.Q , \mchip.opb.dff_gen[0].d1.Q };
	assign \mchip.mult.i3.b_out  = \mchip.mult.i3.temp_register [15:8];
	assign \mchip.mult.i3.clk  = io_in[12];
	assign \mchip.mult.i3.do_add  = \mchip.mult.i0.state [4];
	assign \mchip.mult.i3.do_shift  = \mchip.mult.i0.state [1];
	assign \mchip.mult.i3.mult_out  = \mchip.mult.i3.temp_register [15:0];
	assign \mchip.mult.i3.temp_register [16] = 1'h0;
	assign \mchip.mult.mult_out  = \mchip.mult.i3.temp_register [15:0];
	assign \mchip.mult_res  = \mchip.mult.i3.temp_register [15:0];
	assign \mchip.op_a_out  = {\mchip.opa.dff_gen[7].d1.Q , \mchip.opa.dff_gen[6].d1.Q , \mchip.opa.dff_gen[5].d1.Q , \mchip.opa.dff_gen[4].d1.Q , \mchip.opa.dff_gen[3].d1.Q , \mchip.opa.dff_gen[2].d1.Q , \mchip.opa.dff_gen[1].d1.Q , \mchip.opa.dff_gen[0].d1.Q };
	assign \mchip.op_b_out  = {\mchip.opb.dff_gen[7].d1.Q , \mchip.opb.dff_gen[6].d1.Q , \mchip.opb.dff_gen[5].d1.Q , \mchip.opb.dff_gen[4].d1.Q , \mchip.opb.dff_gen[3].d1.Q , \mchip.opb.dff_gen[2].d1.Q , \mchip.opb.dff_gen[1].d1.Q , \mchip.opb.dff_gen[0].d1.Q };
	assign \mchip.opa.Load_op  = \mchip.control.state [2];
	assign \mchip.opa.dff_gen[0].d1.D  = \mchip.op_a_in [0];
	assign \mchip.opa.dff_gen[0].d1.clk  = \mchip.control.state [2];
	assign \mchip.opa.dff_gen[1].d1.D  = \mchip.op_a_in [1];
	assign \mchip.opa.dff_gen[1].d1.clk  = \mchip.control.state [2];
	assign \mchip.opa.dff_gen[2].d1.D  = \mchip.op_a_in [2];
	assign \mchip.opa.dff_gen[2].d1.clk  = \mchip.control.state [2];
	assign \mchip.opa.dff_gen[3].d1.D  = \mchip.op_a_in [3];
	assign \mchip.opa.dff_gen[3].d1.clk  = \mchip.control.state [2];
	assign \mchip.opa.dff_gen[4].d1.D  = \mchip.op_a_in [4];
	assign \mchip.opa.dff_gen[4].d1.clk  = \mchip.control.state [2];
	assign \mchip.opa.dff_gen[5].d1.D  = \mchip.op_a_in [5];
	assign \mchip.opa.dff_gen[5].d1.clk  = \mchip.control.state [2];
	assign \mchip.opa.dff_gen[6].d1.D  = \mchip.op_a_in [6];
	assign \mchip.opa.dff_gen[6].d1.clk  = \mchip.control.state [2];
	assign \mchip.opa.dff_gen[7].d1.D  = \mchip.op_a_in [7];
	assign \mchip.opa.dff_gen[7].d1.clk  = \mchip.control.state [2];
	assign \mchip.opa.in  = \mchip.op_a_in ;
	assign \mchip.opa.out  = {\mchip.opa.dff_gen[7].d1.Q , \mchip.opa.dff_gen[6].d1.Q , \mchip.opa.dff_gen[5].d1.Q , \mchip.opa.dff_gen[4].d1.Q , \mchip.opa.dff_gen[3].d1.Q , \mchip.opa.dff_gen[2].d1.Q , \mchip.opa.dff_gen[1].d1.Q , \mchip.opa.dff_gen[0].d1.Q };
	assign \mchip.opa.temp_out  = {\mchip.opa.dff_gen[7].d1.Q , \mchip.opa.dff_gen[6].d1.Q , \mchip.opa.dff_gen[5].d1.Q , \mchip.opa.dff_gen[4].d1.Q , \mchip.opa.dff_gen[3].d1.Q , \mchip.opa.dff_gen[2].d1.Q , \mchip.opa.dff_gen[1].d1.Q , \mchip.opa.dff_gen[0].d1.Q };
	assign \mchip.opb.Load_op  = \mchip.control.state [2];
	assign \mchip.opb.dff_gen[0].d1.D  = \mchip.op_b_in [0];
	assign \mchip.opb.dff_gen[0].d1.clk  = \mchip.control.state [2];
	assign \mchip.opb.dff_gen[1].d1.D  = \mchip.op_b_in [1];
	assign \mchip.opb.dff_gen[1].d1.clk  = \mchip.control.state [2];
	assign \mchip.opb.dff_gen[2].d1.D  = \mchip.op_b_in [2];
	assign \mchip.opb.dff_gen[2].d1.clk  = \mchip.control.state [2];
	assign \mchip.opb.dff_gen[3].d1.D  = \mchip.op_b_in [3];
	assign \mchip.opb.dff_gen[3].d1.clk  = \mchip.control.state [2];
	assign \mchip.opb.dff_gen[4].d1.D  = \mchip.op_b_in [4];
	assign \mchip.opb.dff_gen[4].d1.clk  = \mchip.control.state [2];
	assign \mchip.opb.dff_gen[5].d1.D  = \mchip.op_b_in [5];
	assign \mchip.opb.dff_gen[5].d1.clk  = \mchip.control.state [2];
	assign \mchip.opb.dff_gen[6].d1.D  = \mchip.op_b_in [6];
	assign \mchip.opb.dff_gen[6].d1.clk  = \mchip.control.state [2];
	assign \mchip.opb.dff_gen[7].d1.D  = \mchip.op_b_in [7];
	assign \mchip.opb.dff_gen[7].d1.clk  = \mchip.control.state [2];
	assign \mchip.opb.in  = \mchip.op_b_in ;
	assign \mchip.opb.out  = {\mchip.opb.dff_gen[7].d1.Q , \mchip.opb.dff_gen[6].d1.Q , \mchip.opb.dff_gen[5].d1.Q , \mchip.opb.dff_gen[4].d1.Q , \mchip.opb.dff_gen[3].d1.Q , \mchip.opb.dff_gen[2].d1.Q , \mchip.opb.dff_gen[1].d1.Q , \mchip.opb.dff_gen[0].d1.Q };
	assign \mchip.opb.temp_out  = {\mchip.opb.dff_gen[7].d1.Q , \mchip.opb.dff_gen[6].d1.Q , \mchip.opb.dff_gen[5].d1.Q , \mchip.opb.dff_gen[4].d1.Q , \mchip.opb.dff_gen[3].d1.Q , \mchip.opb.dff_gen[2].d1.Q , \mchip.opb.dff_gen[1].d1.Q , \mchip.opb.dff_gen[0].d1.Q };
	assign \mchip.reset  = io_in[13];
endmodule
module d19_rdkapur_encryptor (
	io_in,
	io_out
);
	wire _00000_;
	wire _00001_;
	wire _00002_;
	wire _00003_;
	wire _00004_;
	wire _00005_;
	wire _00006_;
	wire _00007_;
	wire _00008_;
	wire _00009_;
	wire _00010_;
	wire _00011_;
	wire _00012_;
	wire _00013_;
	wire _00014_;
	wire _00015_;
	wire _00016_;
	wire _00017_;
	wire _00018_;
	wire _00019_;
	wire _00020_;
	wire _00021_;
	wire _00022_;
	wire _00023_;
	wire _00024_;
	wire _00025_;
	wire _00026_;
	wire _00027_;
	wire _00028_;
	wire _00029_;
	wire _00030_;
	wire _00031_;
	wire _00032_;
	wire _00033_;
	wire _00034_;
	wire _00035_;
	wire _00036_;
	wire _00037_;
	wire _00038_;
	wire _00039_;
	wire _00040_;
	wire _00041_;
	wire _00042_;
	wire _00043_;
	wire _00044_;
	wire _00045_;
	wire _00046_;
	wire _00047_;
	wire _00048_;
	wire _00049_;
	wire _00050_;
	wire _00051_;
	wire _00052_;
	wire _00053_;
	wire _00054_;
	wire _00055_;
	wire _00056_;
	wire _00057_;
	wire _00058_;
	wire _00059_;
	wire _00060_;
	wire _00061_;
	wire _00062_;
	wire _00063_;
	wire _00064_;
	wire _00065_;
	wire _00066_;
	wire _00067_;
	wire _00068_;
	wire _00069_;
	wire _00070_;
	wire _00071_;
	wire _00072_;
	wire _00073_;
	wire _00074_;
	wire _00075_;
	wire _00076_;
	wire _00077_;
	wire _00078_;
	wire _00079_;
	wire _00080_;
	wire _00081_;
	wire _00082_;
	wire _00083_;
	wire _00084_;
	wire _00085_;
	wire _00086_;
	wire _00087_;
	wire _00088_;
	wire _00089_;
	wire _00090_;
	wire _00091_;
	wire _00092_;
	wire _00093_;
	wire _00094_;
	wire _00095_;
	wire _00096_;
	wire _00097_;
	wire _00098_;
	wire _00099_;
	wire _00100_;
	wire _00101_;
	wire _00102_;
	wire _00103_;
	wire _00104_;
	wire _00105_;
	wire _00106_;
	wire _00107_;
	wire _00108_;
	wire _00109_;
	wire _00110_;
	wire _00111_;
	wire _00112_;
	wire _00113_;
	wire _00114_;
	wire _00115_;
	wire _00116_;
	wire _00117_;
	wire _00118_;
	wire _00119_;
	wire _00120_;
	wire _00121_;
	wire _00122_;
	wire _00123_;
	wire _00124_;
	wire _00125_;
	wire _00126_;
	wire _00127_;
	wire _00128_;
	wire _00129_;
	wire _00130_;
	wire _00131_;
	wire _00132_;
	wire _00133_;
	wire _00134_;
	wire _00135_;
	wire _00136_;
	wire _00137_;
	wire _00138_;
	wire _00139_;
	wire _00140_;
	wire _00141_;
	wire _00142_;
	wire _00143_;
	wire _00144_;
	wire _00145_;
	wire _00146_;
	wire _00147_;
	wire _00148_;
	wire _00149_;
	wire _00150_;
	wire _00151_;
	wire _00152_;
	wire _00153_;
	wire _00154_;
	wire _00155_;
	wire _00156_;
	wire _00157_;
	wire _00158_;
	wire _00159_;
	wire _00160_;
	wire _00161_;
	wire _00162_;
	wire _00163_;
	wire _00164_;
	wire _00165_;
	wire _00166_;
	wire _00167_;
	wire _00168_;
	wire _00169_;
	wire _00170_;
	wire _00171_;
	wire _00172_;
	wire _00173_;
	wire _00174_;
	wire _00175_;
	wire _00176_;
	wire _00177_;
	wire _00178_;
	wire _00179_;
	wire _00180_;
	wire _00181_;
	wire _00182_;
	wire _00183_;
	wire _00184_;
	wire _00185_;
	wire _00186_;
	wire _00187_;
	wire _00188_;
	wire _00189_;
	wire _00190_;
	wire _00191_;
	wire _00192_;
	wire _00193_;
	wire _00194_;
	wire _00195_;
	wire _00196_;
	wire _00197_;
	wire _00198_;
	wire _00199_;
	wire _00200_;
	wire _00201_;
	wire _00202_;
	wire _00203_;
	wire _00204_;
	wire _00205_;
	wire _00206_;
	wire _00207_;
	wire _00208_;
	wire _00209_;
	wire _00210_;
	wire _00211_;
	wire _00212_;
	wire _00213_;
	wire _00214_;
	wire _00215_;
	wire _00216_;
	wire _00217_;
	wire _00218_;
	wire _00219_;
	wire _00220_;
	wire _00221_;
	wire _00222_;
	wire _00223_;
	wire _00224_;
	wire _00225_;
	wire _00226_;
	wire _00227_;
	wire _00228_;
	wire _00229_;
	wire _00230_;
	wire _00231_;
	wire _00232_;
	wire _00233_;
	wire _00234_;
	wire _00235_;
	wire _00236_;
	wire _00237_;
	wire _00238_;
	wire _00239_;
	wire _00240_;
	wire _00241_;
	wire _00242_;
	wire _00243_;
	wire _00244_;
	wire _00245_;
	wire _00246_;
	wire _00247_;
	wire _00248_;
	wire _00249_;
	wire _00250_;
	wire _00251_;
	wire _00252_;
	wire _00253_;
	wire _00254_;
	wire _00255_;
	wire _00256_;
	wire _00257_;
	wire _00258_;
	wire _00259_;
	wire _00260_;
	wire _00261_;
	wire _00262_;
	wire _00263_;
	wire _00264_;
	wire _00265_;
	wire _00266_;
	wire _00267_;
	wire _00268_;
	wire _00269_;
	wire _00270_;
	wire _00271_;
	wire _00272_;
	wire _00273_;
	wire _00274_;
	wire _00275_;
	wire _00276_;
	wire _00277_;
	wire _00278_;
	wire _00279_;
	wire _00280_;
	wire _00281_;
	wire _00282_;
	wire _00283_;
	wire _00284_;
	wire _00285_;
	wire _00286_;
	wire _00287_;
	wire _00288_;
	wire _00289_;
	wire _00290_;
	wire _00291_;
	wire _00292_;
	wire _00293_;
	wire _00294_;
	wire _00295_;
	wire _00296_;
	wire _00297_;
	wire _00298_;
	wire _00299_;
	wire _00300_;
	wire _00301_;
	wire _00302_;
	wire _00303_;
	wire _00304_;
	wire _00305_;
	wire _00306_;
	wire _00307_;
	wire _00308_;
	wire _00309_;
	wire _00310_;
	wire _00311_;
	wire _00312_;
	wire _00313_;
	wire _00314_;
	wire _00315_;
	wire _00316_;
	wire _00317_;
	wire _00318_;
	wire _00319_;
	wire _00320_;
	wire _00321_;
	wire _00322_;
	wire _00323_;
	wire _00324_;
	wire _00325_;
	wire _00326_;
	wire _00327_;
	wire _00328_;
	wire _00329_;
	wire _00330_;
	wire _00331_;
	wire _00332_;
	wire _00333_;
	wire _00334_;
	wire _00335_;
	wire _00336_;
	wire _00337_;
	wire _00338_;
	wire _00339_;
	wire _00340_;
	wire _00341_;
	wire _00342_;
	wire _00343_;
	wire _00344_;
	wire _00345_;
	wire _00346_;
	wire _00347_;
	wire _00348_;
	wire _00349_;
	wire _00350_;
	wire _00351_;
	wire _00352_;
	wire _00353_;
	wire _00354_;
	wire _00355_;
	wire _00356_;
	wire _00357_;
	wire _00358_;
	wire _00359_;
	wire _00360_;
	wire _00361_;
	wire _00362_;
	wire _00363_;
	wire _00364_;
	wire _00365_;
	wire _00366_;
	wire _00367_;
	wire _00368_;
	wire _00369_;
	wire _00370_;
	wire _00371_;
	wire _00372_;
	wire _00373_;
	wire _00374_;
	wire _00375_;
	wire _00376_;
	wire _00377_;
	wire _00378_;
	wire _00379_;
	wire _00380_;
	wire _00381_;
	wire _00382_;
	wire _00383_;
	wire _00384_;
	wire _00385_;
	wire _00386_;
	wire _00387_;
	wire _00388_;
	wire _00389_;
	wire _00390_;
	wire _00391_;
	wire _00392_;
	wire _00393_;
	wire _00394_;
	wire _00395_;
	wire _00396_;
	wire _00397_;
	wire _00398_;
	wire _00399_;
	wire _00400_;
	wire _00401_;
	wire _00402_;
	wire _00403_;
	wire _00404_;
	wire _00405_;
	wire _00406_;
	wire _00407_;
	wire _00408_;
	wire _00409_;
	wire _00410_;
	wire _00411_;
	wire _00412_;
	wire _00413_;
	wire _00414_;
	wire _00415_;
	wire _00416_;
	wire _00417_;
	wire _00418_;
	wire _00419_;
	wire _00420_;
	wire _00421_;
	wire _00422_;
	wire _00423_;
	wire _00424_;
	wire _00425_;
	wire _00426_;
	wire _00427_;
	wire _00428_;
	wire _00429_;
	wire _00430_;
	wire _00431_;
	wire _00432_;
	wire _00433_;
	wire _00434_;
	wire _00435_;
	wire _00436_;
	wire _00437_;
	wire _00438_;
	wire _00439_;
	wire _00440_;
	wire _00441_;
	wire _00442_;
	wire _00443_;
	wire _00444_;
	wire _00445_;
	wire _00446_;
	wire _00447_;
	wire _00448_;
	wire _00449_;
	wire _00450_;
	wire _00451_;
	wire _00452_;
	wire _00453_;
	wire _00454_;
	wire _00455_;
	wire _00456_;
	wire _00457_;
	wire _00458_;
	wire _00459_;
	wire _00460_;
	wire _00461_;
	wire _00462_;
	wire _00463_;
	wire _00464_;
	wire _00465_;
	wire _00466_;
	wire _00467_;
	wire _00468_;
	wire _00469_;
	wire _00470_;
	wire _00471_;
	wire _00472_;
	wire _00473_;
	wire _00474_;
	wire _00475_;
	wire _00476_;
	wire _00477_;
	wire _00478_;
	wire _00479_;
	wire _00480_;
	wire _00481_;
	wire _00482_;
	wire _00483_;
	wire _00484_;
	wire _00485_;
	wire _00486_;
	wire _00487_;
	wire _00488_;
	wire _00489_;
	wire _00490_;
	wire _00491_;
	wire _00492_;
	wire _00493_;
	wire _00494_;
	wire _00495_;
	wire _00496_;
	wire _00497_;
	wire _00498_;
	wire _00499_;
	wire _00500_;
	wire _00501_;
	wire _00502_;
	wire _00503_;
	wire _00504_;
	wire _00505_;
	wire _00506_;
	wire _00507_;
	wire _00508_;
	wire _00509_;
	wire _00510_;
	wire _00511_;
	wire _00512_;
	wire _00513_;
	wire _00514_;
	wire _00515_;
	wire _00516_;
	wire _00517_;
	wire _00518_;
	wire _00519_;
	wire _00520_;
	wire _00521_;
	wire _00522_;
	wire _00523_;
	wire _00524_;
	wire _00525_;
	wire _00526_;
	wire _00527_;
	wire _00528_;
	wire _00529_;
	wire _00530_;
	wire _00531_;
	wire _00532_;
	wire _00533_;
	wire _00534_;
	wire _00535_;
	wire _00536_;
	wire _00537_;
	wire _00538_;
	wire _00539_;
	wire _00540_;
	wire _00541_;
	wire _00542_;
	wire _00543_;
	wire _00544_;
	wire _00545_;
	wire _00546_;
	wire _00547_;
	wire _00548_;
	wire _00549_;
	wire _00550_;
	wire _00551_;
	wire _00552_;
	wire _00553_;
	wire _00554_;
	wire _00555_;
	wire _00556_;
	wire _00557_;
	wire _00558_;
	wire _00559_;
	wire _00560_;
	wire _00561_;
	wire _00562_;
	wire _00563_;
	wire _00564_;
	wire _00565_;
	wire _00566_;
	wire _00567_;
	wire _00568_;
	wire _00569_;
	wire _00570_;
	wire _00571_;
	wire _00572_;
	wire _00573_;
	wire _00574_;
	wire _00575_;
	wire _00576_;
	wire _00577_;
	wire _00578_;
	wire _00579_;
	wire _00580_;
	wire _00581_;
	wire _00582_;
	wire _00583_;
	wire _00584_;
	wire _00585_;
	wire _00586_;
	wire _00587_;
	wire _00588_;
	wire _00589_;
	wire _00590_;
	wire _00591_;
	wire _00592_;
	wire _00593_;
	wire _00594_;
	wire _00595_;
	wire _00596_;
	wire _00597_;
	wire _00598_;
	wire _00599_;
	wire _00600_;
	wire _00601_;
	wire _00602_;
	wire _00603_;
	wire _00604_;
	wire _00605_;
	wire _00606_;
	wire _00607_;
	wire _00608_;
	wire _00609_;
	wire _00610_;
	wire _00611_;
	wire _00612_;
	wire _00613_;
	wire _00614_;
	wire _00615_;
	wire _00616_;
	wire _00617_;
	wire _00618_;
	wire _00619_;
	wire _00620_;
	wire _00621_;
	wire _00622_;
	wire _00623_;
	wire _00624_;
	wire _00625_;
	wire _00626_;
	wire _00627_;
	wire _00628_;
	wire _00629_;
	wire _00630_;
	wire _00631_;
	wire _00632_;
	wire _00633_;
	wire _00634_;
	wire _00635_;
	wire _00636_;
	wire _00637_;
	wire _00638_;
	wire _00639_;
	wire _00640_;
	wire _00641_;
	wire _00642_;
	wire _00643_;
	wire _00644_;
	wire _00645_;
	wire _00646_;
	wire _00647_;
	wire _00648_;
	wire _00649_;
	wire _00650_;
	wire _00651_;
	wire _00652_;
	wire _00653_;
	wire _00654_;
	wire _00655_;
	wire _00656_;
	wire _00657_;
	wire _00658_;
	wire _00659_;
	wire _00660_;
	wire _00661_;
	wire _00662_;
	wire _00663_;
	wire _00664_;
	wire _00665_;
	wire _00666_;
	wire _00667_;
	wire _00668_;
	wire _00669_;
	wire _00670_;
	wire _00671_;
	wire _00672_;
	wire _00673_;
	wire _00674_;
	wire _00675_;
	wire _00676_;
	wire _00677_;
	wire _00678_;
	wire _00679_;
	wire _00680_;
	wire _00681_;
	wire _00682_;
	wire _00683_;
	wire _00684_;
	wire _00685_;
	wire _00686_;
	wire _00687_;
	wire _00688_;
	wire _00689_;
	wire _00690_;
	wire _00691_;
	wire _00692_;
	wire _00693_;
	wire _00694_;
	wire _00695_;
	wire _00696_;
	wire _00697_;
	wire _00698_;
	wire _00699_;
	wire _00700_;
	wire _00701_;
	wire _00702_;
	wire _00703_;
	wire _00704_;
	wire _00705_;
	wire _00706_;
	wire _00707_;
	wire _00708_;
	wire _00709_;
	wire _00710_;
	wire _00711_;
	wire _00712_;
	wire _00713_;
	wire _00714_;
	wire _00715_;
	wire _00716_;
	wire _00717_;
	wire _00718_;
	wire _00719_;
	wire _00720_;
	wire _00721_;
	wire _00722_;
	wire _00723_;
	wire _00724_;
	wire _00725_;
	wire _00726_;
	wire _00727_;
	wire _00728_;
	wire _00729_;
	wire _00730_;
	wire _00731_;
	wire _00732_;
	wire _00733_;
	wire _00734_;
	wire _00735_;
	wire _00736_;
	wire _00737_;
	wire _00738_;
	wire _00739_;
	wire _00740_;
	wire _00741_;
	wire _00742_;
	wire _00743_;
	wire _00744_;
	wire _00745_;
	wire _00746_;
	wire _00747_;
	wire _00748_;
	wire _00749_;
	wire _00750_;
	wire _00751_;
	wire _00752_;
	wire _00753_;
	wire _00754_;
	wire _00755_;
	wire _00756_;
	wire _00757_;
	wire _00758_;
	wire _00759_;
	wire _00760_;
	wire _00761_;
	wire _00762_;
	wire _00763_;
	wire _00764_;
	wire _00765_;
	wire _00766_;
	wire _00767_;
	wire _00768_;
	wire _00769_;
	wire _00770_;
	wire _00771_;
	wire _00772_;
	wire _00773_;
	wire _00774_;
	wire _00775_;
	wire _00776_;
	wire _00777_;
	wire _00778_;
	wire _00779_;
	wire _00780_;
	wire _00781_;
	wire _00782_;
	wire _00783_;
	wire _00784_;
	wire _00785_;
	wire _00786_;
	wire _00787_;
	wire _00788_;
	wire _00789_;
	wire _00790_;
	wire _00791_;
	wire _00792_;
	wire _00793_;
	wire _00794_;
	wire _00795_;
	wire _00796_;
	wire _00797_;
	wire _00798_;
	wire _00799_;
	wire _00800_;
	wire _00801_;
	wire _00802_;
	wire _00803_;
	wire _00804_;
	wire _00805_;
	wire _00806_;
	wire _00807_;
	wire _00808_;
	wire _00809_;
	wire _00810_;
	wire _00811_;
	wire _00812_;
	wire _00813_;
	wire _00814_;
	wire _00815_;
	wire _00816_;
	wire _00817_;
	wire _00818_;
	wire _00819_;
	wire _00820_;
	wire _00821_;
	wire _00822_;
	wire _00823_;
	wire _00824_;
	wire _00825_;
	wire _00826_;
	wire _00827_;
	wire _00828_;
	wire _00829_;
	wire _00830_;
	wire _00831_;
	wire _00832_;
	wire _00833_;
	wire _00834_;
	wire _00835_;
	wire _00836_;
	wire _00837_;
	wire _00838_;
	wire _00839_;
	wire _00840_;
	wire _00841_;
	wire _00842_;
	wire _00843_;
	wire _00844_;
	wire _00845_;
	wire _00846_;
	wire _00847_;
	wire _00848_;
	wire _00849_;
	wire _00850_;
	wire _00851_;
	wire _00852_;
	wire _00853_;
	wire _00854_;
	wire _00855_;
	wire _00856_;
	wire _00857_;
	wire _00858_;
	wire _00859_;
	wire _00860_;
	wire _00861_;
	wire _00862_;
	wire _00863_;
	wire _00864_;
	wire _00865_;
	wire _00866_;
	wire _00867_;
	wire _00868_;
	wire _00869_;
	wire _00870_;
	wire _00871_;
	wire _00872_;
	wire _00873_;
	wire _00874_;
	wire _00875_;
	wire _00876_;
	wire _00877_;
	wire _00878_;
	wire _00879_;
	wire _00880_;
	wire _00881_;
	wire _00882_;
	wire _00883_;
	wire _00884_;
	wire _00885_;
	wire _00886_;
	wire _00887_;
	wire _00888_;
	wire _00889_;
	wire _00890_;
	wire _00891_;
	wire _00892_;
	wire _00893_;
	wire _00894_;
	wire _00895_;
	wire _00896_;
	wire _00897_;
	wire _00898_;
	wire _00899_;
	wire _00900_;
	wire _00901_;
	wire _00902_;
	wire _00903_;
	wire _00904_;
	wire _00905_;
	wire _00906_;
	wire _00907_;
	wire _00908_;
	wire _00909_;
	wire _00910_;
	wire _00911_;
	wire _00912_;
	wire _00913_;
	wire _00914_;
	wire _00915_;
	wire _00916_;
	wire _00917_;
	wire _00918_;
	wire _00919_;
	wire _00920_;
	wire _00921_;
	wire _00922_;
	wire _00923_;
	wire _00924_;
	wire _00925_;
	wire _00926_;
	wire _00927_;
	wire _00928_;
	wire _00929_;
	wire _00930_;
	wire _00931_;
	wire _00932_;
	wire _00933_;
	wire _00934_;
	wire _00935_;
	wire _00936_;
	wire _00937_;
	wire _00938_;
	wire _00939_;
	wire _00940_;
	wire _00941_;
	wire _00942_;
	wire _00943_;
	wire _00944_;
	wire _00945_;
	wire _00946_;
	wire _00947_;
	wire _00948_;
	wire _00949_;
	wire _00950_;
	wire _00951_;
	wire _00952_;
	wire _00953_;
	wire _00954_;
	wire _00955_;
	wire _00956_;
	wire _00957_;
	wire _00958_;
	wire _00959_;
	wire _00960_;
	wire _00961_;
	wire _00962_;
	wire _00963_;
	wire _00964_;
	wire _00965_;
	wire _00966_;
	wire _00967_;
	wire _00968_;
	wire _00969_;
	wire _00970_;
	wire _00971_;
	wire _00972_;
	wire _00973_;
	wire _00974_;
	wire _00975_;
	wire _00976_;
	wire _00977_;
	wire _00978_;
	wire _00979_;
	wire _00980_;
	wire _00981_;
	wire _00982_;
	wire _00983_;
	wire _00984_;
	wire _00985_;
	wire _00986_;
	wire _00987_;
	wire _00988_;
	wire _00989_;
	wire _00990_;
	wire _00991_;
	wire _00992_;
	wire _00993_;
	wire _00994_;
	wire _00995_;
	wire _00996_;
	wire _00997_;
	wire _00998_;
	wire _00999_;
	wire _01000_;
	wire _01001_;
	wire _01002_;
	wire _01003_;
	wire _01004_;
	wire _01005_;
	wire _01006_;
	wire _01007_;
	wire _01008_;
	wire _01009_;
	wire _01010_;
	wire _01011_;
	wire _01012_;
	wire _01013_;
	wire _01014_;
	wire _01015_;
	wire _01016_;
	wire _01017_;
	wire _01018_;
	wire _01019_;
	wire _01020_;
	wire _01021_;
	wire _01022_;
	wire _01023_;
	wire _01024_;
	wire _01025_;
	wire _01026_;
	wire _01027_;
	wire _01028_;
	wire _01029_;
	wire _01030_;
	wire _01031_;
	wire _01032_;
	wire _01033_;
	wire _01034_;
	wire _01035_;
	wire _01036_;
	wire _01037_;
	wire _01038_;
	wire _01039_;
	wire _01040_;
	wire _01041_;
	wire _01042_;
	wire _01043_;
	wire _01044_;
	wire _01045_;
	wire _01046_;
	wire _01047_;
	wire _01048_;
	wire _01049_;
	wire _01050_;
	wire _01051_;
	wire _01052_;
	wire _01053_;
	wire _01054_;
	wire _01055_;
	wire _01056_;
	wire _01057_;
	wire _01058_;
	wire _01059_;
	wire _01060_;
	wire _01061_;
	wire _01062_;
	wire _01063_;
	wire _01064_;
	wire _01065_;
	wire _01066_;
	wire _01067_;
	wire _01068_;
	wire _01069_;
	wire _01070_;
	wire _01071_;
	wire _01072_;
	wire _01073_;
	wire _01074_;
	wire _01075_;
	wire _01076_;
	wire _01077_;
	wire _01078_;
	wire _01079_;
	wire _01080_;
	wire _01081_;
	wire _01082_;
	wire _01083_;
	wire _01084_;
	wire _01085_;
	wire _01086_;
	wire _01087_;
	wire _01088_;
	wire _01089_;
	wire _01090_;
	wire _01091_;
	wire _01092_;
	wire _01093_;
	wire _01094_;
	wire _01095_;
	wire _01096_;
	wire _01097_;
	wire _01098_;
	wire _01099_;
	wire _01100_;
	wire _01101_;
	wire _01102_;
	wire _01103_;
	wire _01104_;
	wire _01105_;
	wire _01106_;
	wire _01107_;
	wire _01108_;
	wire _01109_;
	wire _01110_;
	wire _01111_;
	wire _01112_;
	wire _01113_;
	wire _01114_;
	wire _01115_;
	wire _01116_;
	wire _01117_;
	wire _01118_;
	wire _01119_;
	wire _01120_;
	wire _01121_;
	wire _01122_;
	wire _01123_;
	wire _01124_;
	wire _01125_;
	wire _01126_;
	wire _01127_;
	wire _01128_;
	wire _01129_;
	wire _01130_;
	wire _01131_;
	wire _01132_;
	wire _01133_;
	wire _01134_;
	wire _01135_;
	wire _01136_;
	wire _01137_;
	wire _01138_;
	wire _01139_;
	wire _01140_;
	wire _01141_;
	wire _01142_;
	wire _01143_;
	wire _01144_;
	wire _01145_;
	wire _01146_;
	wire _01147_;
	wire _01148_;
	wire _01149_;
	wire _01150_;
	wire _01151_;
	wire _01152_;
	wire _01153_;
	wire _01154_;
	wire _01155_;
	wire _01156_;
	wire _01157_;
	wire _01158_;
	wire _01159_;
	wire _01160_;
	wire _01161_;
	wire _01162_;
	wire _01163_;
	wire _01164_;
	wire _01165_;
	wire _01166_;
	wire _01167_;
	wire _01168_;
	wire _01169_;
	wire _01170_;
	wire _01171_;
	wire _01172_;
	wire _01173_;
	wire _01174_;
	wire _01175_;
	wire _01176_;
	wire _01177_;
	wire _01178_;
	wire _01179_;
	wire _01180_;
	wire _01181_;
	wire _01182_;
	wire _01183_;
	wire _01184_;
	wire _01185_;
	wire _01186_;
	wire _01187_;
	wire _01188_;
	wire _01189_;
	wire _01190_;
	wire _01191_;
	wire _01192_;
	wire _01193_;
	wire _01194_;
	wire _01195_;
	wire _01196_;
	wire _01197_;
	wire _01198_;
	wire _01199_;
	wire _01200_;
	wire _01201_;
	wire _01202_;
	wire _01203_;
	wire _01204_;
	wire _01205_;
	wire _01206_;
	wire _01207_;
	wire _01208_;
	wire _01209_;
	wire _01210_;
	wire _01211_;
	wire _01212_;
	wire _01213_;
	wire _01214_;
	wire _01215_;
	wire _01216_;
	wire _01217_;
	wire _01218_;
	wire _01219_;
	wire _01220_;
	wire _01221_;
	wire _01222_;
	wire _01223_;
	wire _01224_;
	wire _01225_;
	wire _01226_;
	wire _01227_;
	wire _01228_;
	wire _01229_;
	wire _01230_;
	wire _01231_;
	wire _01232_;
	wire _01233_;
	wire _01234_;
	wire _01235_;
	wire _01236_;
	wire _01237_;
	wire _01238_;
	wire _01239_;
	wire _01240_;
	wire _01241_;
	wire _01242_;
	wire _01243_;
	wire _01244_;
	wire _01245_;
	wire _01246_;
	wire _01247_;
	wire _01248_;
	wire _01249_;
	wire _01250_;
	wire _01251_;
	wire _01252_;
	wire _01253_;
	wire _01254_;
	wire _01255_;
	wire _01256_;
	wire _01257_;
	wire _01258_;
	wire _01259_;
	wire _01260_;
	wire _01261_;
	wire _01262_;
	wire _01263_;
	wire _01264_;
	wire _01265_;
	wire _01266_;
	wire _01267_;
	wire _01268_;
	wire _01269_;
	wire _01270_;
	wire _01271_;
	wire _01272_;
	wire _01273_;
	wire _01274_;
	wire _01275_;
	wire _01276_;
	wire _01277_;
	wire _01278_;
	wire _01279_;
	wire _01280_;
	wire _01281_;
	wire _01282_;
	wire _01283_;
	wire _01284_;
	wire _01285_;
	wire _01286_;
	wire _01287_;
	wire _01288_;
	wire _01289_;
	wire _01290_;
	wire _01291_;
	wire _01292_;
	wire _01293_;
	wire _01294_;
	wire _01295_;
	wire _01296_;
	wire _01297_;
	wire _01298_;
	wire _01299_;
	wire _01300_;
	wire _01301_;
	wire _01302_;
	wire _01303_;
	wire _01304_;
	wire _01305_;
	wire _01306_;
	wire _01307_;
	wire _01308_;
	wire _01309_;
	wire _01310_;
	wire _01311_;
	wire _01312_;
	wire _01313_;
	wire _01314_;
	wire _01315_;
	wire _01316_;
	wire _01317_;
	wire _01318_;
	wire _01319_;
	wire _01320_;
	wire _01321_;
	wire _01322_;
	wire _01323_;
	wire _01324_;
	wire _01325_;
	wire _01326_;
	wire _01327_;
	wire _01328_;
	wire _01329_;
	wire _01330_;
	wire _01331_;
	wire _01332_;
	wire _01333_;
	wire _01334_;
	wire _01335_;
	wire _01336_;
	wire _01337_;
	wire _01338_;
	wire _01339_;
	wire _01340_;
	wire _01341_;
	wire _01342_;
	wire _01343_;
	wire _01344_;
	wire _01345_;
	wire _01346_;
	wire _01347_;
	wire _01348_;
	wire _01349_;
	wire _01350_;
	wire _01351_;
	wire _01352_;
	wire _01353_;
	wire _01354_;
	wire _01355_;
	wire _01356_;
	wire _01357_;
	wire _01358_;
	wire _01359_;
	wire _01360_;
	wire _01361_;
	wire _01362_;
	wire _01363_;
	wire _01364_;
	wire _01365_;
	wire _01366_;
	wire _01367_;
	wire _01368_;
	wire _01369_;
	wire _01370_;
	wire _01371_;
	wire _01372_;
	wire _01373_;
	wire _01374_;
	wire _01375_;
	wire _01376_;
	wire _01377_;
	wire _01378_;
	wire _01379_;
	wire _01380_;
	wire _01381_;
	wire _01382_;
	wire _01383_;
	wire _01384_;
	wire _01385_;
	wire _01386_;
	wire _01387_;
	wire _01388_;
	wire _01389_;
	wire _01390_;
	wire _01391_;
	wire _01392_;
	wire _01393_;
	wire _01394_;
	wire _01395_;
	wire _01396_;
	wire _01397_;
	wire _01398_;
	wire _01399_;
	wire _01400_;
	wire _01401_;
	wire _01402_;
	wire _01403_;
	wire _01404_;
	wire _01405_;
	wire _01406_;
	wire _01407_;
	wire _01408_;
	wire _01409_;
	wire _01410_;
	wire _01411_;
	wire _01412_;
	wire _01413_;
	wire _01414_;
	wire _01415_;
	wire _01416_;
	wire _01417_;
	wire _01418_;
	wire _01419_;
	wire _01420_;
	wire _01421_;
	wire _01422_;
	wire _01423_;
	wire _01424_;
	wire _01425_;
	wire _01426_;
	wire _01427_;
	wire _01428_;
	wire _01429_;
	wire _01430_;
	wire _01431_;
	wire _01432_;
	wire _01433_;
	wire _01434_;
	wire _01435_;
	wire _01436_;
	wire _01437_;
	wire _01438_;
	wire _01439_;
	wire _01440_;
	wire _01441_;
	wire _01442_;
	wire _01443_;
	wire _01444_;
	wire _01445_;
	wire _01446_;
	wire _01447_;
	wire _01448_;
	wire _01449_;
	wire _01450_;
	wire _01451_;
	wire _01452_;
	wire _01453_;
	wire _01454_;
	wire _01455_;
	wire _01456_;
	wire _01457_;
	wire _01458_;
	wire _01459_;
	wire _01460_;
	wire _01461_;
	wire _01462_;
	wire _01463_;
	wire _01464_;
	wire _01465_;
	wire _01466_;
	wire _01467_;
	wire _01468_;
	wire _01469_;
	wire _01470_;
	wire _01471_;
	wire _01472_;
	wire _01473_;
	wire _01474_;
	wire _01475_;
	wire _01476_;
	wire _01477_;
	wire _01478_;
	wire _01479_;
	wire _01480_;
	wire _01481_;
	wire _01482_;
	wire _01483_;
	wire _01484_;
	wire _01485_;
	wire _01486_;
	wire _01487_;
	wire _01488_;
	wire _01489_;
	wire _01490_;
	wire _01491_;
	wire _01492_;
	wire _01493_;
	wire _01494_;
	wire _01495_;
	wire _01496_;
	wire _01497_;
	wire _01498_;
	wire _01499_;
	wire _01500_;
	wire _01501_;
	wire _01502_;
	wire _01503_;
	wire _01504_;
	wire _01505_;
	wire _01506_;
	wire _01507_;
	wire _01508_;
	wire _01509_;
	wire _01510_;
	wire _01511_;
	wire _01512_;
	wire _01513_;
	wire _01514_;
	wire _01515_;
	wire _01516_;
	wire _01517_;
	wire _01518_;
	wire _01519_;
	wire _01520_;
	wire _01521_;
	wire _01522_;
	wire _01523_;
	wire _01524_;
	wire _01525_;
	wire _01526_;
	wire _01527_;
	wire _01528_;
	wire _01529_;
	wire _01530_;
	wire _01531_;
	wire _01532_;
	wire _01533_;
	wire _01534_;
	wire _01535_;
	wire _01536_;
	wire _01537_;
	wire _01538_;
	wire _01539_;
	wire _01540_;
	wire _01541_;
	wire _01542_;
	wire _01543_;
	wire _01544_;
	wire _01545_;
	wire _01546_;
	wire _01547_;
	wire _01548_;
	wire _01549_;
	wire _01550_;
	wire _01551_;
	wire _01552_;
	wire _01553_;
	wire _01554_;
	wire _01555_;
	wire _01556_;
	wire _01557_;
	wire _01558_;
	wire _01559_;
	wire _01560_;
	wire _01561_;
	wire _01562_;
	wire _01563_;
	wire _01564_;
	wire _01565_;
	wire _01566_;
	wire _01567_;
	wire _01568_;
	wire _01569_;
	wire _01570_;
	wire _01571_;
	wire _01572_;
	wire _01573_;
	wire _01574_;
	wire _01575_;
	wire _01576_;
	wire _01577_;
	wire _01578_;
	wire _01579_;
	wire _01580_;
	wire _01581_;
	wire _01582_;
	wire _01583_;
	wire _01584_;
	wire _01585_;
	wire _01586_;
	wire _01587_;
	wire _01588_;
	wire _01589_;
	wire _01590_;
	wire _01591_;
	wire _01592_;
	wire _01593_;
	wire _01594_;
	wire _01595_;
	wire _01596_;
	wire _01597_;
	wire _01598_;
	wire _01599_;
	wire _01600_;
	wire _01601_;
	wire _01602_;
	wire _01603_;
	wire _01604_;
	wire _01605_;
	wire _01606_;
	wire _01607_;
	wire _01608_;
	wire _01609_;
	wire _01610_;
	wire _01611_;
	wire _01612_;
	wire _01613_;
	wire _01614_;
	wire _01615_;
	wire _01616_;
	wire _01617_;
	wire _01618_;
	wire _01619_;
	wire _01620_;
	wire _01621_;
	wire _01622_;
	wire _01623_;
	wire _01624_;
	wire _01625_;
	wire _01626_;
	wire _01627_;
	wire _01628_;
	wire _01629_;
	wire _01630_;
	wire _01631_;
	wire _01632_;
	wire _01633_;
	wire _01634_;
	wire _01635_;
	wire _01636_;
	wire _01637_;
	wire _01638_;
	wire _01639_;
	wire _01640_;
	wire _01641_;
	wire _01642_;
	wire _01643_;
	wire _01644_;
	wire _01645_;
	wire _01646_;
	wire _01647_;
	wire _01648_;
	wire _01649_;
	wire _01650_;
	wire _01651_;
	wire _01652_;
	wire _01653_;
	wire _01654_;
	wire _01655_;
	wire _01656_;
	wire _01657_;
	wire _01658_;
	wire _01659_;
	wire _01660_;
	wire _01661_;
	wire _01662_;
	wire _01663_;
	wire _01664_;
	wire _01665_;
	wire _01666_;
	wire _01667_;
	wire _01668_;
	wire _01669_;
	wire _01670_;
	wire _01671_;
	wire _01672_;
	wire _01673_;
	wire _01674_;
	wire _01675_;
	wire _01676_;
	wire _01677_;
	wire _01678_;
	wire _01679_;
	wire _01680_;
	wire _01681_;
	wire _01682_;
	wire _01683_;
	wire _01684_;
	wire _01685_;
	wire _01686_;
	wire _01687_;
	wire _01688_;
	wire _01689_;
	wire _01690_;
	wire _01691_;
	wire _01692_;
	wire _01693_;
	wire _01694_;
	wire _01695_;
	wire _01696_;
	wire _01697_;
	wire _01698_;
	wire _01699_;
	wire _01700_;
	wire _01701_;
	wire _01702_;
	wire _01703_;
	wire _01704_;
	wire _01705_;
	wire _01706_;
	wire _01707_;
	wire _01708_;
	wire _01709_;
	wire _01710_;
	wire _01711_;
	wire _01712_;
	wire _01713_;
	wire _01714_;
	wire _01715_;
	wire _01716_;
	wire _01717_;
	wire _01718_;
	wire _01719_;
	wire _01720_;
	wire _01721_;
	wire _01722_;
	wire _01723_;
	wire _01724_;
	wire _01725_;
	wire _01726_;
	wire _01727_;
	wire _01728_;
	wire _01729_;
	wire _01730_;
	wire _01731_;
	wire _01732_;
	wire _01733_;
	wire _01734_;
	wire _01735_;
	wire _01736_;
	wire _01737_;
	wire _01738_;
	wire _01739_;
	wire _01740_;
	wire _01741_;
	wire _01742_;
	wire _01743_;
	wire _01744_;
	wire _01745_;
	wire _01746_;
	wire _01747_;
	wire _01748_;
	wire _01749_;
	wire _01750_;
	wire _01751_;
	wire _01752_;
	wire _01753_;
	wire _01754_;
	wire _01755_;
	wire _01756_;
	wire _01757_;
	wire _01758_;
	wire _01759_;
	wire _01760_;
	wire _01761_;
	wire _01762_;
	wire _01763_;
	wire _01764_;
	wire _01765_;
	wire _01766_;
	wire _01767_;
	wire _01768_;
	wire _01769_;
	wire _01770_;
	wire _01771_;
	wire _01772_;
	wire _01773_;
	wire _01774_;
	wire _01775_;
	wire _01776_;
	wire _01777_;
	wire _01778_;
	wire _01779_;
	wire _01780_;
	wire _01781_;
	wire _01782_;
	wire _01783_;
	wire _01784_;
	wire _01785_;
	wire _01786_;
	wire _01787_;
	wire _01788_;
	wire _01789_;
	wire _01790_;
	wire _01791_;
	wire _01792_;
	wire _01793_;
	wire _01794_;
	wire _01795_;
	wire _01796_;
	wire _01797_;
	wire _01798_;
	wire _01799_;
	wire _01800_;
	wire _01801_;
	wire _01802_;
	wire _01803_;
	wire _01804_;
	wire _01805_;
	wire _01806_;
	wire _01807_;
	wire _01808_;
	wire _01809_;
	wire _01810_;
	wire _01811_;
	wire _01812_;
	wire _01813_;
	wire _01814_;
	wire _01815_;
	wire _01816_;
	wire _01817_;
	wire _01818_;
	wire _01819_;
	wire _01820_;
	wire _01821_;
	wire _01822_;
	wire _01823_;
	wire _01824_;
	wire _01825_;
	wire _01826_;
	wire _01827_;
	wire _01828_;
	wire _01829_;
	wire _01830_;
	wire _01831_;
	wire _01832_;
	wire _01833_;
	wire _01834_;
	wire _01835_;
	wire _01836_;
	wire _01837_;
	wire _01838_;
	wire _01839_;
	wire _01840_;
	wire _01841_;
	wire _01842_;
	wire _01843_;
	wire _01844_;
	wire _01845_;
	wire _01846_;
	wire _01847_;
	wire _01848_;
	wire _01849_;
	wire _01850_;
	wire _01851_;
	wire _01852_;
	wire _01853_;
	wire _01854_;
	wire _01855_;
	wire _01856_;
	wire _01857_;
	wire _01858_;
	wire _01859_;
	wire _01860_;
	wire _01861_;
	wire _01862_;
	wire _01863_;
	wire _01864_;
	wire _01865_;
	wire _01866_;
	wire _01867_;
	wire _01868_;
	wire _01869_;
	wire _01870_;
	wire _01871_;
	wire _01872_;
	wire _01873_;
	wire _01874_;
	wire _01875_;
	wire _01876_;
	wire _01877_;
	wire _01878_;
	wire _01879_;
	wire _01880_;
	wire _01881_;
	wire _01882_;
	wire _01883_;
	wire _01884_;
	wire _01885_;
	wire _01886_;
	wire _01887_;
	wire _01888_;
	wire _01889_;
	wire _01890_;
	wire _01891_;
	wire _01892_;
	wire _01893_;
	wire _01894_;
	wire _01895_;
	wire _01896_;
	wire _01897_;
	wire _01898_;
	wire _01899_;
	wire _01900_;
	wire _01901_;
	wire _01902_;
	wire _01903_;
	wire _01904_;
	wire _01905_;
	wire _01906_;
	wire _01907_;
	wire _01908_;
	wire _01909_;
	wire _01910_;
	wire _01911_;
	wire _01912_;
	wire _01913_;
	wire _01914_;
	wire _01915_;
	wire _01916_;
	wire _01917_;
	wire _01918_;
	wire _01919_;
	wire _01920_;
	wire _01921_;
	wire _01922_;
	wire _01923_;
	wire _01924_;
	wire _01925_;
	wire _01926_;
	wire _01927_;
	wire _01928_;
	wire _01929_;
	wire _01930_;
	wire _01931_;
	wire _01932_;
	wire _01933_;
	wire _01934_;
	wire _01935_;
	wire _01936_;
	wire _01937_;
	wire _01938_;
	wire _01939_;
	wire _01940_;
	wire _01941_;
	wire _01942_;
	wire _01943_;
	wire _01944_;
	wire _01945_;
	wire _01946_;
	wire _01947_;
	wire _01948_;
	wire _01949_;
	wire _01950_;
	wire _01951_;
	wire _01952_;
	wire _01953_;
	wire _01954_;
	wire _01955_;
	wire _01956_;
	wire _01957_;
	wire _01958_;
	wire _01959_;
	wire _01960_;
	wire _01961_;
	wire _01962_;
	wire _01963_;
	wire _01964_;
	wire _01965_;
	wire _01966_;
	wire _01967_;
	wire _01968_;
	wire _01969_;
	wire _01970_;
	wire _01971_;
	wire _01972_;
	wire _01973_;
	wire _01974_;
	wire _01975_;
	wire _01976_;
	wire _01977_;
	wire _01978_;
	wire _01979_;
	wire _01980_;
	wire _01981_;
	wire _01982_;
	wire _01983_;
	wire _01984_;
	wire _01985_;
	wire _01986_;
	wire _01987_;
	wire _01988_;
	wire _01989_;
	wire _01990_;
	wire _01991_;
	wire _01992_;
	wire _01993_;
	wire _01994_;
	wire _01995_;
	wire _01996_;
	wire _01997_;
	wire _01998_;
	wire _01999_;
	wire _02000_;
	wire _02001_;
	wire _02002_;
	wire _02003_;
	wire _02004_;
	wire _02005_;
	wire _02006_;
	wire _02007_;
	wire _02008_;
	wire _02009_;
	wire _02010_;
	wire _02011_;
	wire _02012_;
	wire _02013_;
	wire _02014_;
	wire _02015_;
	wire _02016_;
	wire _02017_;
	wire _02018_;
	wire _02019_;
	wire _02020_;
	wire _02021_;
	wire _02022_;
	wire _02023_;
	wire _02024_;
	wire _02025_;
	wire _02026_;
	wire _02027_;
	wire _02028_;
	wire _02029_;
	wire _02030_;
	wire _02031_;
	wire _02032_;
	wire _02033_;
	wire _02034_;
	wire _02035_;
	wire _02036_;
	wire _02037_;
	wire _02038_;
	wire _02039_;
	wire _02040_;
	wire _02041_;
	wire _02042_;
	wire _02043_;
	wire _02044_;
	wire _02045_;
	wire _02046_;
	wire _02047_;
	wire _02048_;
	wire _02049_;
	wire _02050_;
	wire _02051_;
	wire _02052_;
	wire _02053_;
	wire _02054_;
	wire _02055_;
	wire _02056_;
	wire _02057_;
	wire _02058_;
	wire _02059_;
	wire _02060_;
	wire _02061_;
	wire _02062_;
	wire _02063_;
	wire _02064_;
	wire _02065_;
	wire _02066_;
	wire _02067_;
	wire _02068_;
	wire _02069_;
	wire _02070_;
	wire _02071_;
	wire _02072_;
	wire _02073_;
	wire _02074_;
	wire _02075_;
	wire _02076_;
	wire _02077_;
	wire _02078_;
	wire _02079_;
	wire _02080_;
	wire _02081_;
	wire _02082_;
	wire _02083_;
	wire _02084_;
	wire _02085_;
	wire _02086_;
	wire _02087_;
	wire _02088_;
	wire _02089_;
	wire _02090_;
	wire _02091_;
	wire _02092_;
	wire _02093_;
	wire _02094_;
	wire _02095_;
	wire _02096_;
	wire _02097_;
	wire _02098_;
	wire _02099_;
	wire _02100_;
	wire _02101_;
	wire _02102_;
	wire _02103_;
	wire _02104_;
	wire _02105_;
	wire _02106_;
	wire _02107_;
	wire _02108_;
	wire _02109_;
	wire _02110_;
	wire _02111_;
	wire _02112_;
	wire _02113_;
	wire _02114_;
	wire _02115_;
	wire _02116_;
	wire _02117_;
	wire _02118_;
	wire _02119_;
	wire _02120_;
	wire _02121_;
	wire _02122_;
	wire _02123_;
	wire _02124_;
	wire _02125_;
	wire _02126_;
	wire _02127_;
	wire _02128_;
	wire _02129_;
	wire _02130_;
	wire _02131_;
	wire _02132_;
	wire _02133_;
	wire _02134_;
	wire _02135_;
	wire _02136_;
	wire _02137_;
	wire _02138_;
	wire _02139_;
	wire _02140_;
	wire _02141_;
	wire _02142_;
	wire _02143_;
	wire _02144_;
	wire _02145_;
	wire _02146_;
	wire _02147_;
	wire _02148_;
	wire _02149_;
	wire _02150_;
	wire _02151_;
	wire _02152_;
	wire _02153_;
	wire _02154_;
	wire _02155_;
	wire _02156_;
	wire _02157_;
	wire _02158_;
	wire _02159_;
	wire _02160_;
	wire _02161_;
	wire _02162_;
	wire _02163_;
	wire _02164_;
	wire _02165_;
	wire _02166_;
	wire _02167_;
	wire _02168_;
	wire _02169_;
	wire _02170_;
	wire _02171_;
	wire _02172_;
	wire _02173_;
	wire _02174_;
	wire _02175_;
	wire _02176_;
	wire _02177_;
	wire _02178_;
	wire _02179_;
	wire _02180_;
	wire _02181_;
	wire _02182_;
	wire _02183_;
	wire _02184_;
	wire _02185_;
	wire _02186_;
	wire _02187_;
	wire _02188_;
	wire _02189_;
	wire _02190_;
	wire _02191_;
	wire _02192_;
	wire _02193_;
	wire _02194_;
	wire _02195_;
	wire _02196_;
	wire _02197_;
	wire _02198_;
	wire _02199_;
	wire _02200_;
	wire _02201_;
	wire _02202_;
	wire _02203_;
	wire _02204_;
	wire _02205_;
	wire _02206_;
	wire _02207_;
	wire _02208_;
	wire _02209_;
	wire _02210_;
	wire _02211_;
	wire _02212_;
	wire _02213_;
	wire _02214_;
	wire _02215_;
	wire _02216_;
	wire _02217_;
	wire _02218_;
	wire _02219_;
	wire _02220_;
	wire _02221_;
	wire _02222_;
	wire _02223_;
	wire _02224_;
	wire _02225_;
	wire _02226_;
	wire _02227_;
	wire _02228_;
	wire _02229_;
	wire _02230_;
	wire _02231_;
	wire _02232_;
	wire _02233_;
	wire _02234_;
	wire _02235_;
	wire _02236_;
	wire _02237_;
	wire _02238_;
	wire _02239_;
	wire _02240_;
	wire _02241_;
	wire _02242_;
	wire _02243_;
	wire _02244_;
	wire _02245_;
	wire _02246_;
	wire _02247_;
	wire _02248_;
	wire _02249_;
	wire _02250_;
	wire _02251_;
	wire _02252_;
	wire _02253_;
	wire _02254_;
	wire _02255_;
	wire _02256_;
	wire _02257_;
	wire _02258_;
	wire _02259_;
	wire _02260_;
	wire _02261_;
	wire _02262_;
	wire _02263_;
	wire _02264_;
	wire _02265_;
	wire _02266_;
	wire _02267_;
	wire _02268_;
	wire _02269_;
	wire _02270_;
	wire _02271_;
	wire _02272_;
	wire _02273_;
	wire _02274_;
	wire _02275_;
	wire _02276_;
	wire _02277_;
	wire _02278_;
	wire _02279_;
	wire _02280_;
	wire _02281_;
	wire _02282_;
	wire _02283_;
	wire _02284_;
	wire _02285_;
	wire _02286_;
	wire _02287_;
	wire _02288_;
	wire _02289_;
	wire _02290_;
	wire _02291_;
	wire _02292_;
	wire _02293_;
	wire _02294_;
	wire _02295_;
	wire _02296_;
	wire _02297_;
	wire _02298_;
	wire _02299_;
	wire _02300_;
	wire _02301_;
	wire _02302_;
	wire _02303_;
	wire _02304_;
	wire _02305_;
	wire _02306_;
	wire _02307_;
	wire _02308_;
	wire _02309_;
	wire _02310_;
	wire _02311_;
	wire _02312_;
	wire _02313_;
	wire _02314_;
	wire _02315_;
	wire _02316_;
	wire _02317_;
	wire _02318_;
	wire _02319_;
	wire _02320_;
	wire _02321_;
	wire _02322_;
	wire _02323_;
	wire _02324_;
	wire _02325_;
	wire _02326_;
	wire _02327_;
	wire _02328_;
	wire _02329_;
	wire _02330_;
	wire _02331_;
	wire _02332_;
	wire _02333_;
	wire _02334_;
	wire _02335_;
	wire _02336_;
	wire _02337_;
	wire _02338_;
	wire _02339_;
	wire _02340_;
	wire _02341_;
	wire _02342_;
	wire _02343_;
	wire _02344_;
	wire _02345_;
	wire _02346_;
	wire _02347_;
	wire _02348_;
	wire _02349_;
	wire _02350_;
	wire _02351_;
	wire _02352_;
	wire _02353_;
	wire _02354_;
	wire _02355_;
	wire _02356_;
	wire _02357_;
	wire _02358_;
	wire _02359_;
	wire _02360_;
	wire _02361_;
	wire _02362_;
	wire _02363_;
	wire _02364_;
	wire _02365_;
	wire _02366_;
	wire _02367_;
	wire _02368_;
	wire _02369_;
	wire _02370_;
	wire _02371_;
	wire _02372_;
	wire _02373_;
	wire _02374_;
	wire _02375_;
	wire _02376_;
	wire _02377_;
	wire _02378_;
	wire _02379_;
	wire _02380_;
	wire _02381_;
	wire _02382_;
	wire _02383_;
	wire _02384_;
	wire _02385_;
	wire _02386_;
	wire _02387_;
	wire _02388_;
	wire _02389_;
	wire _02390_;
	wire _02391_;
	wire _02392_;
	wire _02393_;
	wire _02394_;
	wire _02395_;
	wire _02396_;
	wire _02397_;
	wire _02398_;
	wire _02399_;
	wire _02400_;
	wire _02401_;
	wire _02402_;
	wire _02403_;
	wire _02404_;
	wire _02405_;
	wire _02406_;
	wire _02407_;
	wire _02408_;
	wire _02409_;
	wire _02410_;
	wire _02411_;
	wire _02412_;
	wire _02413_;
	wire _02414_;
	wire _02415_;
	wire _02416_;
	wire _02417_;
	wire _02418_;
	wire _02419_;
	wire _02420_;
	wire _02421_;
	wire _02422_;
	wire _02423_;
	wire _02424_;
	wire _02425_;
	wire _02426_;
	wire _02427_;
	wire _02428_;
	wire _02429_;
	wire _02430_;
	wire _02431_;
	wire _02432_;
	wire _02433_;
	wire _02434_;
	wire _02435_;
	wire _02436_;
	wire _02437_;
	wire _02438_;
	wire _02439_;
	wire _02440_;
	wire _02441_;
	wire _02442_;
	wire _02443_;
	wire _02444_;
	wire _02445_;
	wire _02446_;
	wire _02447_;
	wire _02448_;
	wire _02449_;
	wire _02450_;
	wire _02451_;
	wire _02452_;
	wire _02453_;
	wire _02454_;
	wire _02455_;
	wire _02456_;
	wire _02457_;
	wire _02458_;
	wire _02459_;
	wire _02460_;
	wire _02461_;
	wire _02462_;
	wire _02463_;
	wire _02464_;
	wire _02465_;
	wire _02466_;
	wire _02467_;
	wire _02468_;
	wire _02469_;
	wire _02470_;
	wire _02471_;
	wire _02472_;
	wire _02473_;
	wire _02474_;
	wire _02475_;
	wire _02476_;
	wire _02477_;
	wire _02478_;
	wire _02479_;
	wire _02480_;
	wire _02481_;
	wire _02482_;
	wire _02483_;
	wire _02484_;
	wire _02485_;
	wire _02486_;
	wire _02487_;
	wire _02488_;
	wire _02489_;
	wire _02490_;
	wire _02491_;
	wire _02492_;
	wire _02493_;
	wire _02494_;
	wire _02495_;
	wire _02496_;
	wire _02497_;
	wire _02498_;
	wire _02499_;
	wire _02500_;
	wire _02501_;
	wire _02502_;
	wire _02503_;
	wire _02504_;
	wire _02505_;
	wire _02506_;
	wire _02507_;
	wire _02508_;
	wire _02509_;
	wire _02510_;
	wire _02511_;
	wire _02512_;
	wire _02513_;
	wire _02514_;
	wire _02515_;
	wire _02516_;
	wire _02517_;
	wire _02518_;
	wire _02519_;
	wire _02520_;
	wire _02521_;
	wire _02522_;
	wire _02523_;
	wire _02524_;
	wire _02525_;
	wire _02526_;
	wire _02527_;
	wire _02528_;
	wire _02529_;
	wire _02530_;
	wire _02531_;
	wire _02532_;
	wire _02533_;
	wire _02534_;
	wire _02535_;
	wire _02536_;
	wire _02537_;
	wire _02538_;
	wire _02539_;
	wire _02540_;
	wire _02541_;
	wire _02542_;
	wire _02543_;
	wire _02544_;
	wire _02545_;
	wire _02546_;
	wire _02547_;
	wire _02548_;
	wire _02549_;
	wire _02550_;
	wire _02551_;
	wire _02552_;
	wire _02553_;
	wire _02554_;
	wire _02555_;
	wire _02556_;
	wire _02557_;
	wire _02558_;
	wire _02559_;
	wire _02560_;
	wire _02561_;
	wire _02562_;
	wire _02563_;
	wire _02564_;
	wire _02565_;
	wire _02566_;
	wire _02567_;
	wire _02568_;
	wire _02569_;
	wire _02570_;
	wire _02571_;
	wire _02572_;
	wire _02573_;
	wire _02574_;
	wire _02575_;
	wire _02576_;
	wire _02577_;
	wire _02578_;
	wire _02579_;
	wire _02580_;
	wire _02581_;
	wire _02582_;
	wire _02583_;
	wire _02584_;
	wire _02585_;
	wire _02586_;
	wire _02587_;
	wire _02588_;
	wire _02589_;
	wire _02590_;
	wire _02591_;
	wire _02592_;
	wire _02593_;
	wire _02594_;
	wire _02595_;
	wire _02596_;
	wire _02597_;
	wire _02598_;
	wire _02599_;
	wire _02600_;
	wire _02601_;
	wire _02602_;
	wire _02603_;
	wire _02604_;
	wire _02605_;
	wire _02606_;
	wire _02607_;
	wire _02608_;
	wire _02609_;
	wire _02610_;
	wire _02611_;
	wire _02612_;
	wire _02613_;
	wire _02614_;
	wire _02615_;
	wire _02616_;
	wire _02617_;
	wire _02618_;
	wire _02619_;
	wire _02620_;
	wire _02621_;
	wire _02622_;
	wire _02623_;
	wire _02624_;
	wire _02625_;
	wire _02626_;
	wire _02627_;
	wire _02628_;
	wire _02629_;
	wire _02630_;
	wire _02631_;
	wire _02632_;
	wire _02633_;
	wire _02634_;
	wire _02635_;
	wire _02636_;
	wire _02637_;
	wire _02638_;
	wire _02639_;
	wire _02640_;
	wire _02641_;
	wire _02642_;
	wire _02643_;
	wire _02644_;
	wire _02645_;
	wire _02646_;
	wire _02647_;
	wire _02648_;
	wire _02649_;
	wire _02650_;
	wire _02651_;
	wire _02652_;
	wire _02653_;
	wire _02654_;
	wire _02655_;
	wire _02656_;
	wire _02657_;
	wire _02658_;
	wire _02659_;
	wire _02660_;
	wire _02661_;
	wire _02662_;
	wire _02663_;
	wire _02664_;
	wire _02665_;
	wire _02666_;
	wire _02667_;
	wire _02668_;
	wire _02669_;
	wire _02670_;
	wire _02671_;
	wire _02672_;
	wire _02673_;
	wire _02674_;
	wire _02675_;
	wire _02676_;
	wire _02677_;
	wire _02678_;
	wire _02679_;
	wire _02680_;
	wire _02681_;
	wire _02682_;
	wire _02683_;
	wire _02684_;
	wire _02685_;
	wire _02686_;
	wire _02687_;
	wire _02688_;
	wire _02689_;
	wire _02690_;
	wire _02691_;
	wire _02692_;
	wire _02693_;
	wire _02694_;
	wire _02695_;
	wire _02696_;
	wire _02697_;
	wire _02698_;
	wire _02699_;
	wire _02700_;
	wire _02701_;
	wire _02702_;
	wire _02703_;
	wire _02704_;
	wire _02705_;
	wire _02706_;
	wire _02707_;
	wire _02708_;
	wire _02709_;
	wire _02710_;
	wire _02711_;
	wire _02712_;
	wire _02713_;
	wire _02714_;
	wire _02715_;
	wire _02716_;
	wire _02717_;
	wire _02718_;
	wire _02719_;
	wire _02720_;
	wire _02721_;
	wire _02722_;
	wire _02723_;
	wire _02724_;
	wire _02725_;
	wire _02726_;
	wire _02727_;
	wire _02728_;
	wire _02729_;
	wire _02730_;
	wire _02731_;
	wire _02732_;
	wire _02733_;
	wire _02734_;
	wire _02735_;
	wire _02736_;
	wire _02737_;
	wire _02738_;
	wire _02739_;
	wire _02740_;
	wire _02741_;
	wire _02742_;
	wire _02743_;
	wire _02744_;
	wire _02745_;
	wire _02746_;
	wire _02747_;
	wire _02748_;
	wire _02749_;
	wire _02750_;
	wire _02751_;
	wire _02752_;
	wire _02753_;
	wire _02754_;
	wire _02755_;
	wire _02756_;
	wire _02757_;
	wire _02758_;
	wire _02759_;
	wire _02760_;
	wire _02761_;
	wire _02762_;
	wire _02763_;
	wire _02764_;
	wire _02765_;
	wire _02766_;
	wire _02767_;
	wire _02768_;
	wire _02769_;
	wire _02770_;
	wire _02771_;
	wire _02772_;
	wire _02773_;
	wire _02774_;
	wire _02775_;
	wire _02776_;
	wire _02777_;
	wire _02778_;
	wire _02779_;
	wire _02780_;
	wire _02781_;
	wire _02782_;
	wire _02783_;
	wire _02784_;
	wire _02785_;
	wire _02786_;
	wire _02787_;
	wire _02788_;
	wire _02789_;
	wire _02790_;
	wire _02791_;
	wire _02792_;
	wire _02793_;
	wire _02794_;
	wire _02795_;
	wire _02796_;
	wire _02797_;
	wire _02798_;
	wire _02799_;
	wire _02800_;
	wire _02801_;
	wire _02802_;
	wire _02803_;
	wire _02804_;
	wire _02805_;
	wire _02806_;
	wire _02807_;
	wire _02808_;
	wire _02809_;
	wire _02810_;
	wire _02811_;
	wire _02812_;
	wire _02813_;
	wire _02814_;
	wire _02815_;
	wire _02816_;
	wire _02817_;
	wire _02818_;
	wire _02819_;
	wire _02820_;
	wire _02821_;
	wire _02822_;
	wire _02823_;
	wire _02824_;
	wire _02825_;
	wire _02826_;
	wire _02827_;
	wire _02828_;
	wire _02829_;
	wire _02830_;
	wire _02831_;
	wire _02832_;
	wire _02833_;
	wire _02834_;
	wire _02835_;
	wire _02836_;
	wire _02837_;
	wire _02838_;
	wire _02839_;
	wire _02840_;
	wire _02841_;
	wire _02842_;
	wire _02843_;
	wire _02844_;
	wire _02845_;
	wire _02846_;
	wire _02847_;
	wire _02848_;
	wire _02849_;
	wire _02850_;
	wire _02851_;
	wire _02852_;
	wire _02853_;
	wire _02854_;
	wire _02855_;
	wire _02856_;
	wire _02857_;
	wire _02858_;
	wire _02859_;
	wire _02860_;
	wire _02861_;
	wire _02862_;
	wire _02863_;
	wire _02864_;
	wire _02865_;
	wire _02866_;
	wire _02867_;
	wire _02868_;
	wire _02869_;
	wire _02870_;
	wire _02871_;
	wire _02872_;
	wire _02873_;
	wire _02874_;
	wire _02875_;
	wire _02876_;
	wire _02877_;
	wire _02878_;
	wire _02879_;
	wire _02880_;
	wire _02881_;
	wire _02882_;
	wire _02883_;
	wire _02884_;
	wire _02885_;
	wire _02886_;
	wire _02887_;
	wire _02888_;
	wire _02889_;
	wire _02890_;
	wire _02891_;
	wire _02892_;
	wire _02893_;
	wire _02894_;
	wire _02895_;
	wire _02896_;
	wire _02897_;
	wire _02898_;
	wire _02899_;
	wire _02900_;
	wire _02901_;
	wire _02902_;
	wire _02903_;
	wire _02904_;
	wire _02905_;
	wire _02906_;
	wire _02907_;
	wire _02908_;
	wire _02909_;
	wire _02910_;
	wire _02911_;
	wire _02912_;
	wire _02913_;
	wire _02914_;
	wire _02915_;
	wire _02916_;
	wire _02917_;
	wire _02918_;
	wire _02919_;
	wire _02920_;
	wire _02921_;
	wire _02922_;
	wire _02923_;
	wire _02924_;
	wire _02925_;
	wire _02926_;
	wire _02927_;
	wire _02928_;
	wire _02929_;
	wire _02930_;
	wire _02931_;
	wire _02932_;
	wire _02933_;
	wire _02934_;
	wire _02935_;
	wire _02936_;
	wire _02937_;
	wire _02938_;
	wire _02939_;
	wire _02940_;
	wire _02941_;
	wire _02942_;
	wire _02943_;
	wire _02944_;
	wire _02945_;
	wire _02946_;
	wire _02947_;
	wire _02948_;
	wire _02949_;
	wire _02950_;
	wire _02951_;
	wire _02952_;
	wire _02953_;
	wire _02954_;
	wire _02955_;
	wire _02956_;
	wire _02957_;
	wire _02958_;
	wire _02959_;
	wire _02960_;
	wire _02961_;
	wire _02962_;
	wire _02963_;
	wire _02964_;
	wire _02965_;
	wire _02966_;
	wire _02967_;
	wire _02968_;
	wire _02969_;
	wire _02970_;
	wire _02971_;
	wire _02972_;
	wire _02973_;
	wire _02974_;
	wire _02975_;
	wire _02976_;
	wire _02977_;
	wire _02978_;
	wire _02979_;
	wire _02980_;
	wire _02981_;
	wire _02982_;
	wire _02983_;
	wire _02984_;
	wire _02985_;
	wire _02986_;
	wire _02987_;
	wire _02988_;
	wire _02989_;
	wire _02990_;
	wire _02991_;
	wire _02992_;
	wire _02993_;
	wire _02994_;
	wire _02995_;
	wire _02996_;
	wire _02997_;
	wire _02998_;
	wire _02999_;
	wire _03000_;
	wire _03001_;
	wire _03002_;
	wire _03003_;
	wire _03004_;
	wire _03005_;
	wire _03006_;
	wire _03007_;
	wire _03008_;
	wire _03009_;
	wire _03010_;
	wire _03011_;
	wire _03012_;
	wire _03013_;
	wire _03014_;
	wire _03015_;
	wire _03016_;
	wire _03017_;
	wire _03018_;
	wire _03019_;
	wire _03020_;
	wire _03021_;
	wire _03022_;
	wire _03023_;
	wire _03024_;
	wire _03025_;
	wire _03026_;
	wire _03027_;
	wire _03028_;
	wire _03029_;
	wire _03030_;
	wire _03031_;
	wire _03032_;
	wire _03033_;
	wire _03034_;
	wire _03035_;
	wire _03036_;
	wire _03037_;
	wire _03038_;
	wire _03039_;
	wire _03040_;
	wire _03041_;
	wire _03042_;
	wire _03043_;
	wire _03044_;
	wire _03045_;
	wire _03046_;
	wire _03047_;
	wire _03048_;
	wire _03049_;
	wire _03050_;
	wire _03051_;
	wire _03052_;
	wire _03053_;
	wire _03054_;
	wire _03055_;
	wire _03056_;
	wire _03057_;
	wire _03058_;
	wire _03059_;
	wire _03060_;
	wire _03061_;
	wire _03062_;
	wire _03063_;
	wire _03064_;
	wire _03065_;
	wire _03066_;
	wire _03067_;
	wire _03068_;
	wire _03069_;
	wire _03070_;
	wire _03071_;
	wire _03072_;
	wire _03073_;
	wire _03074_;
	wire _03075_;
	wire _03076_;
	wire _03077_;
	wire _03078_;
	wire _03079_;
	wire _03080_;
	wire _03081_;
	wire _03082_;
	wire _03083_;
	wire _03084_;
	wire _03085_;
	wire _03086_;
	wire _03087_;
	wire _03088_;
	wire _03089_;
	wire _03090_;
	wire _03091_;
	wire _03092_;
	wire _03093_;
	wire _03094_;
	wire _03095_;
	wire _03096_;
	wire _03097_;
	wire _03098_;
	wire _03099_;
	wire _03100_;
	wire _03101_;
	wire _03102_;
	wire _03103_;
	wire _03104_;
	wire _03105_;
	wire _03106_;
	wire _03107_;
	wire _03108_;
	wire _03109_;
	wire _03110_;
	wire _03111_;
	wire _03112_;
	wire _03113_;
	wire _03114_;
	wire _03115_;
	wire _03116_;
	wire _03117_;
	wire _03118_;
	wire _03119_;
	wire _03120_;
	wire _03121_;
	wire _03122_;
	wire _03123_;
	wire _03124_;
	wire _03125_;
	wire _03126_;
	wire _03127_;
	wire _03128_;
	wire _03129_;
	wire _03130_;
	wire _03131_;
	wire _03132_;
	wire _03133_;
	wire _03134_;
	wire _03135_;
	wire _03136_;
	wire _03137_;
	wire _03138_;
	wire _03139_;
	wire _03140_;
	wire _03141_;
	wire _03142_;
	wire _03143_;
	wire _03144_;
	wire _03145_;
	wire _03146_;
	wire _03147_;
	wire _03148_;
	wire _03149_;
	wire _03150_;
	wire _03151_;
	wire _03152_;
	wire _03153_;
	wire _03154_;
	wire _03155_;
	wire _03156_;
	wire _03157_;
	wire _03158_;
	wire _03159_;
	wire _03160_;
	wire _03161_;
	wire _03162_;
	wire _03163_;
	wire _03164_;
	wire _03165_;
	wire _03166_;
	wire _03167_;
	wire _03168_;
	wire _03169_;
	wire _03170_;
	wire _03171_;
	wire _03172_;
	wire _03173_;
	wire _03174_;
	wire _03175_;
	wire _03176_;
	wire _03177_;
	wire _03178_;
	wire _03179_;
	wire _03180_;
	wire _03181_;
	wire _03182_;
	wire _03183_;
	wire _03184_;
	wire _03185_;
	wire _03186_;
	wire _03187_;
	wire _03188_;
	wire _03189_;
	wire _03190_;
	wire _03191_;
	wire _03192_;
	wire _03193_;
	wire _03194_;
	wire _03195_;
	wire _03196_;
	wire _03197_;
	wire _03198_;
	wire _03199_;
	wire _03200_;
	wire _03201_;
	wire _03202_;
	wire _03203_;
	wire _03204_;
	wire _03205_;
	wire _03206_;
	wire _03207_;
	wire _03208_;
	wire _03209_;
	wire _03210_;
	wire _03211_;
	wire _03212_;
	wire _03213_;
	wire _03214_;
	wire _03215_;
	wire _03216_;
	wire _03217_;
	wire _03218_;
	wire _03219_;
	wire _03220_;
	wire _03221_;
	wire _03222_;
	wire _03223_;
	wire _03224_;
	wire _03225_;
	wire _03226_;
	wire _03227_;
	wire _03228_;
	wire _03229_;
	wire _03230_;
	wire _03231_;
	wire _03232_;
	wire _03233_;
	wire _03234_;
	wire _03235_;
	wire _03236_;
	wire _03237_;
	wire _03238_;
	wire _03239_;
	wire _03240_;
	wire _03241_;
	wire _03242_;
	wire _03243_;
	wire _03244_;
	wire _03245_;
	wire _03246_;
	wire _03247_;
	wire _03248_;
	wire _03249_;
	wire _03250_;
	wire _03251_;
	wire _03252_;
	wire _03253_;
	wire _03254_;
	wire _03255_;
	wire _03256_;
	wire _03257_;
	wire _03258_;
	wire _03259_;
	wire _03260_;
	wire _03261_;
	wire _03262_;
	wire _03263_;
	wire _03264_;
	wire _03265_;
	wire _03266_;
	wire _03267_;
	wire _03268_;
	wire _03269_;
	wire _03270_;
	wire _03271_;
	wire _03272_;
	wire _03273_;
	wire _03274_;
	wire _03275_;
	wire _03276_;
	wire _03277_;
	wire _03278_;
	wire _03279_;
	wire _03280_;
	wire _03281_;
	wire _03282_;
	wire _03283_;
	wire _03284_;
	wire _03285_;
	wire _03286_;
	wire _03287_;
	wire _03288_;
	wire _03289_;
	wire _03290_;
	wire _03291_;
	wire _03292_;
	wire _03293_;
	wire _03294_;
	wire _03295_;
	wire _03296_;
	wire _03297_;
	wire _03298_;
	wire _03299_;
	wire _03300_;
	wire _03301_;
	wire _03302_;
	wire _03303_;
	wire _03304_;
	wire _03305_;
	wire _03306_;
	wire _03307_;
	wire _03308_;
	wire _03309_;
	wire _03310_;
	wire _03311_;
	wire _03312_;
	wire _03313_;
	wire _03314_;
	wire _03315_;
	wire _03316_;
	wire _03317_;
	wire _03318_;
	wire _03319_;
	wire _03320_;
	wire _03321_;
	wire _03322_;
	wire _03323_;
	wire _03324_;
	wire _03325_;
	wire _03326_;
	wire _03327_;
	wire _03328_;
	wire _03329_;
	wire _03330_;
	wire _03331_;
	wire _03332_;
	wire _03333_;
	wire _03334_;
	wire _03335_;
	wire _03336_;
	wire _03337_;
	wire _03338_;
	wire _03339_;
	wire _03340_;
	wire _03341_;
	wire _03342_;
	wire _03343_;
	wire _03344_;
	wire _03345_;
	wire _03346_;
	wire _03347_;
	wire _03348_;
	wire _03349_;
	wire _03350_;
	wire _03351_;
	wire _03352_;
	wire _03353_;
	wire _03354_;
	wire _03355_;
	wire _03356_;
	wire _03357_;
	wire _03358_;
	wire _03359_;
	wire _03360_;
	wire _03361_;
	wire _03362_;
	wire _03363_;
	wire _03364_;
	wire _03365_;
	wire _03366_;
	wire _03367_;
	wire _03368_;
	wire _03369_;
	wire _03370_;
	wire _03371_;
	wire _03372_;
	wire _03373_;
	wire _03374_;
	wire _03375_;
	wire _03376_;
	wire _03377_;
	wire _03378_;
	wire _03379_;
	wire _03380_;
	wire _03381_;
	wire _03382_;
	wire _03383_;
	wire _03384_;
	wire _03385_;
	wire _03386_;
	wire _03387_;
	wire _03388_;
	wire _03389_;
	wire _03390_;
	wire _03391_;
	wire _03392_;
	wire _03393_;
	wire _03394_;
	wire _03395_;
	wire _03396_;
	wire _03397_;
	wire _03398_;
	wire _03399_;
	wire _03400_;
	wire _03401_;
	wire _03402_;
	wire _03403_;
	wire _03404_;
	wire _03405_;
	wire _03406_;
	wire _03407_;
	wire _03408_;
	wire _03409_;
	wire _03410_;
	wire _03411_;
	wire _03412_;
	wire _03413_;
	wire _03414_;
	wire _03415_;
	wire _03416_;
	wire _03417_;
	wire _03418_;
	wire _03419_;
	wire _03420_;
	wire _03421_;
	wire _03422_;
	wire _03423_;
	wire _03424_;
	wire _03425_;
	wire _03426_;
	wire _03427_;
	wire _03428_;
	wire _03429_;
	wire _03430_;
	wire _03431_;
	wire _03432_;
	wire _03433_;
	wire _03434_;
	wire _03435_;
	wire _03436_;
	wire _03437_;
	wire _03438_;
	wire _03439_;
	wire _03440_;
	wire _03441_;
	wire _03442_;
	wire _03443_;
	wire _03444_;
	wire _03445_;
	wire _03446_;
	wire _03447_;
	wire _03448_;
	wire _03449_;
	wire _03450_;
	wire _03451_;
	wire _03452_;
	wire _03453_;
	wire _03454_;
	wire _03455_;
	wire _03456_;
	wire _03457_;
	wire _03458_;
	wire _03459_;
	wire _03460_;
	wire _03461_;
	wire _03462_;
	wire _03463_;
	wire _03464_;
	wire _03465_;
	wire _03466_;
	wire _03467_;
	wire _03468_;
	wire _03469_;
	wire _03470_;
	wire _03471_;
	wire _03472_;
	wire _03473_;
	wire _03474_;
	wire _03475_;
	wire _03476_;
	wire _03477_;
	wire _03478_;
	wire _03479_;
	wire _03480_;
	wire _03481_;
	wire _03482_;
	wire _03483_;
	wire _03484_;
	wire _03485_;
	wire _03486_;
	wire _03487_;
	wire _03488_;
	wire _03489_;
	wire _03490_;
	wire _03491_;
	wire _03492_;
	wire _03493_;
	wire _03494_;
	wire _03495_;
	wire _03496_;
	wire _03497_;
	wire _03498_;
	wire _03499_;
	wire _03500_;
	wire _03501_;
	wire _03502_;
	wire _03503_;
	wire _03504_;
	wire _03505_;
	wire _03506_;
	wire _03507_;
	wire _03508_;
	wire _03509_;
	wire _03510_;
	wire _03511_;
	wire _03512_;
	wire _03513_;
	wire _03514_;
	wire _03515_;
	wire _03516_;
	wire _03517_;
	wire _03518_;
	wire _03519_;
	wire _03520_;
	wire _03521_;
	wire _03522_;
	wire _03523_;
	wire _03524_;
	wire _03525_;
	wire _03526_;
	wire _03527_;
	wire _03528_;
	wire _03529_;
	wire _03530_;
	wire _03531_;
	wire _03532_;
	wire _03533_;
	wire _03534_;
	wire _03535_;
	wire _03536_;
	wire _03537_;
	wire _03538_;
	wire _03539_;
	wire _03540_;
	wire _03541_;
	wire _03542_;
	wire _03543_;
	wire _03544_;
	wire _03545_;
	wire _03546_;
	wire _03547_;
	wire _03548_;
	wire _03549_;
	wire _03550_;
	wire _03551_;
	wire _03552_;
	wire _03553_;
	wire _03554_;
	wire _03555_;
	wire _03556_;
	wire _03557_;
	wire _03558_;
	wire _03559_;
	wire _03560_;
	wire _03561_;
	wire _03562_;
	wire _03563_;
	wire _03564_;
	wire _03565_;
	wire _03566_;
	wire _03567_;
	wire _03568_;
	wire _03569_;
	wire _03570_;
	wire _03571_;
	wire _03572_;
	wire _03573_;
	wire _03574_;
	wire _03575_;
	wire _03576_;
	wire _03577_;
	wire _03578_;
	wire _03579_;
	wire _03580_;
	wire _03581_;
	wire _03582_;
	wire _03583_;
	wire _03584_;
	wire _03585_;
	wire _03586_;
	wire _03587_;
	wire _03588_;
	wire _03589_;
	wire _03590_;
	wire _03591_;
	wire _03592_;
	wire _03593_;
	wire _03594_;
	wire _03595_;
	wire _03596_;
	wire _03597_;
	wire _03598_;
	wire _03599_;
	wire _03600_;
	wire _03601_;
	wire _03602_;
	wire _03603_;
	wire _03604_;
	wire _03605_;
	wire _03606_;
	wire _03607_;
	wire _03608_;
	wire _03609_;
	wire _03610_;
	wire _03611_;
	wire _03612_;
	wire _03613_;
	wire _03614_;
	wire _03615_;
	wire _03616_;
	wire _03617_;
	wire _03618_;
	wire _03619_;
	wire _03620_;
	wire _03621_;
	wire _03622_;
	wire _03623_;
	wire _03624_;
	wire _03625_;
	wire _03626_;
	wire _03627_;
	wire _03628_;
	wire _03629_;
	wire _03630_;
	wire _03631_;
	wire _03632_;
	wire _03633_;
	wire _03634_;
	wire _03635_;
	wire _03636_;
	wire _03637_;
	wire _03638_;
	wire _03639_;
	wire _03640_;
	wire _03641_;
	wire _03642_;
	wire _03643_;
	wire _03644_;
	wire _03645_;
	wire _03646_;
	wire _03647_;
	wire _03648_;
	wire _03649_;
	wire _03650_;
	wire _03651_;
	wire _03652_;
	wire _03653_;
	wire _03654_;
	wire _03655_;
	wire _03656_;
	wire _03657_;
	wire _03658_;
	wire _03659_;
	wire _03660_;
	wire _03661_;
	wire _03662_;
	wire _03663_;
	wire _03664_;
	wire _03665_;
	wire _03666_;
	wire _03667_;
	wire _03668_;
	wire _03669_;
	wire _03670_;
	wire _03671_;
	wire _03672_;
	wire _03673_;
	wire _03674_;
	wire _03675_;
	wire _03676_;
	wire _03677_;
	wire _03678_;
	wire _03679_;
	wire _03680_;
	wire _03681_;
	wire _03682_;
	wire _03683_;
	wire _03684_;
	wire _03685_;
	wire _03686_;
	wire _03687_;
	wire _03688_;
	wire _03689_;
	wire _03690_;
	wire _03691_;
	wire _03692_;
	wire _03693_;
	wire _03694_;
	wire _03695_;
	wire _03696_;
	wire _03697_;
	wire _03698_;
	wire _03699_;
	wire _03700_;
	wire _03701_;
	wire _03702_;
	wire _03703_;
	wire _03704_;
	wire _03705_;
	wire _03706_;
	wire _03707_;
	wire _03708_;
	wire _03709_;
	wire _03710_;
	wire _03711_;
	wire _03712_;
	wire _03713_;
	wire _03714_;
	wire _03715_;
	wire _03716_;
	wire _03717_;
	wire _03718_;
	wire _03719_;
	wire _03720_;
	wire _03721_;
	wire _03722_;
	wire _03723_;
	wire _03724_;
	wire _03725_;
	wire _03726_;
	wire _03727_;
	wire _03728_;
	wire _03729_;
	wire _03730_;
	wire _03731_;
	wire _03732_;
	wire _03733_;
	wire _03734_;
	wire _03735_;
	wire _03736_;
	wire _03737_;
	wire _03738_;
	wire _03739_;
	wire _03740_;
	wire _03741_;
	wire _03742_;
	wire _03743_;
	wire _03744_;
	wire _03745_;
	wire _03746_;
	wire _03747_;
	wire _03748_;
	wire _03749_;
	wire _03750_;
	wire _03751_;
	wire _03752_;
	wire _03753_;
	wire _03754_;
	wire _03755_;
	wire _03756_;
	wire _03757_;
	wire _03758_;
	wire _03759_;
	wire _03760_;
	wire _03761_;
	wire _03762_;
	wire _03763_;
	wire _03764_;
	wire _03765_;
	wire _03766_;
	wire _03767_;
	wire _03768_;
	wire _03769_;
	wire _03770_;
	wire _03771_;
	wire _03772_;
	wire _03773_;
	wire _03774_;
	wire _03775_;
	wire _03776_;
	wire _03777_;
	wire _03778_;
	wire _03779_;
	wire _03780_;
	wire _03781_;
	wire _03782_;
	wire _03783_;
	wire _03784_;
	wire _03785_;
	wire _03786_;
	wire _03787_;
	wire _03788_;
	wire _03789_;
	wire _03790_;
	wire _03791_;
	wire _03792_;
	wire _03793_;
	wire _03794_;
	wire _03795_;
	wire _03796_;
	wire _03797_;
	wire _03798_;
	wire _03799_;
	wire _03800_;
	wire _03801_;
	wire _03802_;
	wire _03803_;
	wire _03804_;
	wire _03805_;
	wire _03806_;
	wire _03807_;
	wire _03808_;
	wire _03809_;
	wire _03810_;
	wire _03811_;
	wire _03812_;
	wire _03813_;
	wire _03814_;
	wire _03815_;
	wire _03816_;
	wire _03817_;
	wire _03818_;
	wire _03819_;
	wire _03820_;
	wire _03821_;
	wire _03822_;
	wire _03823_;
	wire _03824_;
	wire _03825_;
	wire _03826_;
	wire _03827_;
	wire _03828_;
	wire _03829_;
	wire _03830_;
	wire _03831_;
	wire _03832_;
	wire _03833_;
	wire _03834_;
	wire _03835_;
	wire _03836_;
	wire _03837_;
	wire _03838_;
	wire _03839_;
	wire _03840_;
	wire _03841_;
	wire _03842_;
	wire _03843_;
	wire _03844_;
	wire _03845_;
	wire _03846_;
	wire _03847_;
	wire _03848_;
	wire _03849_;
	wire _03850_;
	wire _03851_;
	wire _03852_;
	wire _03853_;
	wire _03854_;
	wire _03855_;
	wire _03856_;
	wire _03857_;
	wire _03858_;
	wire _03859_;
	wire _03860_;
	wire _03861_;
	wire _03862_;
	wire _03863_;
	wire _03864_;
	wire _03865_;
	wire _03866_;
	wire _03867_;
	wire _03868_;
	wire _03869_;
	wire _03870_;
	wire _03871_;
	wire _03872_;
	wire _03873_;
	wire _03874_;
	wire _03875_;
	wire _03876_;
	wire _03877_;
	wire _03878_;
	wire _03879_;
	wire _03880_;
	wire _03881_;
	wire _03882_;
	wire _03883_;
	wire _03884_;
	wire _03885_;
	wire _03886_;
	wire _03887_;
	wire _03888_;
	wire _03889_;
	wire _03890_;
	wire _03891_;
	wire _03892_;
	wire _03893_;
	wire _03894_;
	wire _03895_;
	wire _03896_;
	wire _03897_;
	wire _03898_;
	wire _03899_;
	wire _03900_;
	wire _03901_;
	wire _03902_;
	wire _03903_;
	wire _03904_;
	wire _03905_;
	wire _03906_;
	wire _03907_;
	wire _03908_;
	wire _03909_;
	wire _03910_;
	wire _03911_;
	wire _03912_;
	wire _03913_;
	wire _03914_;
	wire _03915_;
	wire _03916_;
	wire _03917_;
	wire _03918_;
	wire _03919_;
	wire _03920_;
	wire _03921_;
	wire _03922_;
	wire _03923_;
	wire _03924_;
	wire _03925_;
	wire _03926_;
	wire _03927_;
	wire _03928_;
	wire _03929_;
	wire _03930_;
	wire _03931_;
	wire _03932_;
	wire _03933_;
	wire _03934_;
	wire _03935_;
	wire _03936_;
	wire _03937_;
	wire _03938_;
	wire _03939_;
	wire _03940_;
	wire _03941_;
	wire _03942_;
	wire _03943_;
	wire _03944_;
	wire _03945_;
	wire _03946_;
	wire _03947_;
	wire _03948_;
	wire _03949_;
	wire _03950_;
	wire _03951_;
	wire _03952_;
	wire _03953_;
	wire _03954_;
	wire _03955_;
	wire _03956_;
	wire _03957_;
	wire _03958_;
	wire _03959_;
	wire _03960_;
	wire _03961_;
	wire _03962_;
	wire _03963_;
	wire _03964_;
	wire _03965_;
	wire _03966_;
	wire _03967_;
	wire _03968_;
	wire _03969_;
	wire _03970_;
	wire _03971_;
	wire _03972_;
	wire _03973_;
	wire _03974_;
	wire _03975_;
	wire _03976_;
	wire _03977_;
	wire _03978_;
	wire _03979_;
	wire _03980_;
	wire _03981_;
	wire _03982_;
	wire _03983_;
	wire _03984_;
	wire _03985_;
	wire _03986_;
	wire _03987_;
	wire _03988_;
	wire _03989_;
	wire _03990_;
	wire _03991_;
	wire _03992_;
	wire _03993_;
	wire _03994_;
	wire _03995_;
	wire _03996_;
	wire _03997_;
	wire _03998_;
	wire _03999_;
	wire _04000_;
	wire _04001_;
	wire _04002_;
	wire _04003_;
	wire _04004_;
	wire _04005_;
	wire _04006_;
	wire _04007_;
	wire _04008_;
	wire _04009_;
	wire _04010_;
	wire _04011_;
	wire _04012_;
	wire _04013_;
	wire _04014_;
	wire _04015_;
	wire _04016_;
	wire _04017_;
	wire _04018_;
	wire _04019_;
	wire _04020_;
	wire _04021_;
	wire _04022_;
	wire _04023_;
	wire _04024_;
	wire _04025_;
	wire _04026_;
	wire _04027_;
	wire _04028_;
	wire _04029_;
	wire _04030_;
	wire _04031_;
	wire _04032_;
	wire _04033_;
	wire _04034_;
	wire _04035_;
	wire _04036_;
	wire _04037_;
	wire _04038_;
	wire _04039_;
	wire _04040_;
	wire _04041_;
	wire _04042_;
	wire _04043_;
	wire _04044_;
	wire _04045_;
	wire _04046_;
	wire _04047_;
	wire _04048_;
	wire _04049_;
	wire _04050_;
	wire _04051_;
	wire _04052_;
	wire _04053_;
	wire _04054_;
	wire _04055_;
	wire _04056_;
	wire _04057_;
	wire _04058_;
	wire _04059_;
	wire _04060_;
	wire _04061_;
	wire _04062_;
	wire _04063_;
	wire _04064_;
	wire _04065_;
	wire _04066_;
	wire _04067_;
	wire _04068_;
	wire _04069_;
	wire _04070_;
	wire _04071_;
	wire _04072_;
	wire _04073_;
	wire _04074_;
	wire _04075_;
	wire _04076_;
	wire _04077_;
	wire _04078_;
	wire _04079_;
	wire _04080_;
	wire _04081_;
	wire _04082_;
	wire _04083_;
	wire _04084_;
	wire _04085_;
	wire _04086_;
	wire _04087_;
	wire _04088_;
	wire _04089_;
	wire _04090_;
	wire _04091_;
	wire _04092_;
	wire _04093_;
	wire _04094_;
	wire _04095_;
	wire _04096_;
	wire _04097_;
	wire _04098_;
	wire _04099_;
	wire _04100_;
	wire _04101_;
	wire _04102_;
	wire _04103_;
	wire _04104_;
	wire _04105_;
	wire _04106_;
	wire _04107_;
	wire _04108_;
	wire _04109_;
	wire _04110_;
	wire _04111_;
	wire _04112_;
	wire _04113_;
	wire _04114_;
	wire _04115_;
	wire _04116_;
	wire _04117_;
	wire _04118_;
	wire _04119_;
	wire _04120_;
	wire _04121_;
	wire _04122_;
	wire _04123_;
	wire _04124_;
	wire _04125_;
	wire _04126_;
	wire _04127_;
	wire _04128_;
	wire _04129_;
	wire _04130_;
	wire _04131_;
	wire _04132_;
	wire _04133_;
	wire _04134_;
	wire _04135_;
	wire _04136_;
	wire _04137_;
	wire _04138_;
	wire _04139_;
	wire _04140_;
	wire _04141_;
	wire _04142_;
	wire _04143_;
	wire _04144_;
	wire _04145_;
	wire _04146_;
	wire _04147_;
	wire _04148_;
	wire _04149_;
	wire _04150_;
	wire _04151_;
	wire _04152_;
	wire _04153_;
	wire _04154_;
	wire _04155_;
	wire _04156_;
	wire _04157_;
	wire _04158_;
	wire _04159_;
	wire _04160_;
	wire _04161_;
	wire _04162_;
	wire _04163_;
	wire _04164_;
	wire _04165_;
	wire _04166_;
	wire _04167_;
	wire _04168_;
	wire _04169_;
	wire _04170_;
	wire _04171_;
	wire _04172_;
	wire _04173_;
	wire _04174_;
	wire _04175_;
	wire _04176_;
	wire _04177_;
	wire _04178_;
	wire _04179_;
	wire _04180_;
	wire _04181_;
	wire _04182_;
	wire _04183_;
	wire _04184_;
	wire _04185_;
	wire _04186_;
	wire _04187_;
	wire _04188_;
	wire _04189_;
	wire _04190_;
	wire _04191_;
	wire _04192_;
	wire _04193_;
	wire _04194_;
	wire _04195_;
	wire _04196_;
	wire _04197_;
	wire _04198_;
	wire _04199_;
	wire _04200_;
	wire _04201_;
	wire _04202_;
	wire _04203_;
	wire _04204_;
	wire _04205_;
	wire _04206_;
	wire _04207_;
	wire _04208_;
	wire _04209_;
	wire _04210_;
	wire _04211_;
	wire _04212_;
	wire _04213_;
	wire _04214_;
	wire _04215_;
	wire _04216_;
	wire _04217_;
	wire _04218_;
	wire _04219_;
	wire _04220_;
	wire _04221_;
	wire _04222_;
	wire _04223_;
	wire _04224_;
	wire _04225_;
	wire _04226_;
	wire _04227_;
	wire _04228_;
	wire _04229_;
	wire _04230_;
	wire _04231_;
	wire _04232_;
	wire _04233_;
	wire _04234_;
	wire _04235_;
	wire _04236_;
	wire _04237_;
	wire _04238_;
	wire _04239_;
	wire _04240_;
	wire _04241_;
	wire _04242_;
	wire _04243_;
	wire _04244_;
	wire _04245_;
	wire _04246_;
	wire _04247_;
	wire _04248_;
	wire _04249_;
	wire _04250_;
	wire _04251_;
	wire _04252_;
	wire _04253_;
	wire _04254_;
	wire _04255_;
	wire _04256_;
	wire _04257_;
	wire _04258_;
	wire _04259_;
	wire _04260_;
	wire _04261_;
	wire _04262_;
	wire _04263_;
	wire _04264_;
	wire _04265_;
	wire _04266_;
	wire _04267_;
	wire _04268_;
	wire _04269_;
	wire _04270_;
	wire _04271_;
	wire _04272_;
	wire _04273_;
	wire _04274_;
	wire _04275_;
	wire _04276_;
	wire _04277_;
	wire _04278_;
	wire _04279_;
	wire _04280_;
	wire _04281_;
	wire _04282_;
	wire _04283_;
	wire _04284_;
	wire _04285_;
	wire _04286_;
	wire _04287_;
	wire _04288_;
	wire _04289_;
	wire _04290_;
	wire _04291_;
	wire _04292_;
	wire _04293_;
	wire _04294_;
	wire _04295_;
	wire _04296_;
	wire _04297_;
	wire _04298_;
	wire _04299_;
	wire _04300_;
	wire _04301_;
	wire _04302_;
	wire _04303_;
	wire _04304_;
	wire _04305_;
	wire _04306_;
	wire _04307_;
	wire _04308_;
	wire _04309_;
	wire _04310_;
	wire _04311_;
	wire _04312_;
	wire _04313_;
	wire _04314_;
	wire _04315_;
	wire _04316_;
	wire _04317_;
	wire _04318_;
	wire _04319_;
	wire _04320_;
	wire _04321_;
	wire _04322_;
	wire _04323_;
	wire _04324_;
	wire _04325_;
	wire _04326_;
	wire _04327_;
	wire _04328_;
	wire _04329_;
	wire _04330_;
	wire _04331_;
	wire _04332_;
	wire _04333_;
	wire _04334_;
	wire _04335_;
	wire _04336_;
	wire _04337_;
	wire _04338_;
	wire _04339_;
	wire _04340_;
	wire _04341_;
	wire _04342_;
	wire _04343_;
	wire _04344_;
	wire _04345_;
	wire _04346_;
	wire _04347_;
	wire _04348_;
	wire _04349_;
	wire _04350_;
	wire _04351_;
	wire _04352_;
	wire _04353_;
	wire _04354_;
	wire _04355_;
	wire _04356_;
	wire _04357_;
	wire _04358_;
	wire _04359_;
	wire _04360_;
	wire _04361_;
	wire _04362_;
	wire _04363_;
	wire _04364_;
	wire _04365_;
	wire _04366_;
	wire _04367_;
	wire _04368_;
	wire _04369_;
	wire _04370_;
	wire _04371_;
	wire _04372_;
	wire _04373_;
	wire _04374_;
	wire _04375_;
	wire _04376_;
	wire _04377_;
	wire _04378_;
	wire _04379_;
	wire _04380_;
	wire _04381_;
	wire _04382_;
	wire _04383_;
	wire _04384_;
	wire _04385_;
	wire _04386_;
	wire _04387_;
	wire _04388_;
	wire _04389_;
	wire _04390_;
	wire _04391_;
	wire _04392_;
	wire _04393_;
	wire _04394_;
	wire _04395_;
	wire _04396_;
	wire _04397_;
	wire _04398_;
	wire _04399_;
	wire _04400_;
	wire _04401_;
	wire _04402_;
	wire _04403_;
	wire _04404_;
	wire _04405_;
	wire _04406_;
	wire _04407_;
	wire _04408_;
	wire _04409_;
	wire _04410_;
	wire _04411_;
	wire _04412_;
	wire _04413_;
	wire _04414_;
	wire _04415_;
	wire _04416_;
	wire _04417_;
	wire _04418_;
	wire _04419_;
	wire _04420_;
	wire _04421_;
	wire _04422_;
	wire _04423_;
	wire _04424_;
	wire _04425_;
	wire _04426_;
	wire _04427_;
	wire _04428_;
	wire _04429_;
	wire _04430_;
	wire _04431_;
	wire _04432_;
	wire _04433_;
	wire _04434_;
	wire _04435_;
	wire _04436_;
	wire _04437_;
	wire _04438_;
	wire _04439_;
	wire _04440_;
	wire _04441_;
	wire _04442_;
	wire _04443_;
	wire _04444_;
	wire _04445_;
	wire _04446_;
	wire _04447_;
	wire _04448_;
	wire _04449_;
	wire _04450_;
	wire _04451_;
	wire _04452_;
	wire _04453_;
	wire _04454_;
	wire _04455_;
	wire _04456_;
	wire _04457_;
	wire _04458_;
	wire _04459_;
	wire _04460_;
	wire _04461_;
	wire _04462_;
	wire _04463_;
	wire _04464_;
	wire _04465_;
	wire _04466_;
	wire _04467_;
	wire _04468_;
	wire _04469_;
	wire _04470_;
	wire _04471_;
	wire _04472_;
	wire _04473_;
	wire _04474_;
	wire _04475_;
	wire _04476_;
	wire _04477_;
	wire _04478_;
	wire _04479_;
	wire _04480_;
	wire _04481_;
	wire _04482_;
	wire _04483_;
	wire _04484_;
	wire _04485_;
	wire _04486_;
	wire _04487_;
	wire _04488_;
	wire _04489_;
	wire _04490_;
	wire _04491_;
	wire _04492_;
	wire _04493_;
	wire _04494_;
	wire _04495_;
	wire _04496_;
	wire _04497_;
	wire _04498_;
	wire _04499_;
	wire _04500_;
	wire _04501_;
	wire _04502_;
	wire _04503_;
	wire _04504_;
	wire _04505_;
	wire _04506_;
	wire _04507_;
	wire _04508_;
	wire _04509_;
	wire _04510_;
	wire _04511_;
	wire _04512_;
	wire _04513_;
	wire _04514_;
	wire _04515_;
	wire _04516_;
	wire _04517_;
	wire _04518_;
	wire _04519_;
	wire _04520_;
	wire _04521_;
	wire _04522_;
	wire _04523_;
	wire _04524_;
	wire _04525_;
	wire _04526_;
	wire _04527_;
	wire _04528_;
	wire _04529_;
	wire _04530_;
	wire _04531_;
	wire _04532_;
	wire _04533_;
	wire _04534_;
	wire _04535_;
	wire _04536_;
	wire _04537_;
	wire _04538_;
	wire _04539_;
	wire _04540_;
	wire _04541_;
	wire _04542_;
	wire _04543_;
	wire _04544_;
	wire _04545_;
	wire _04546_;
	wire _04547_;
	wire _04548_;
	wire _04549_;
	wire _04550_;
	wire _04551_;
	wire _04552_;
	wire _04553_;
	wire _04554_;
	wire _04555_;
	wire _04556_;
	wire _04557_;
	wire _04558_;
	wire _04559_;
	wire _04560_;
	wire _04561_;
	wire _04562_;
	wire _04563_;
	wire _04564_;
	wire _04565_;
	wire _04566_;
	wire _04567_;
	wire _04568_;
	wire _04569_;
	wire _04570_;
	wire _04571_;
	wire _04572_;
	wire _04573_;
	wire _04574_;
	wire _04575_;
	wire _04576_;
	wire _04577_;
	wire _04578_;
	wire _04579_;
	wire _04580_;
	wire _04581_;
	wire _04582_;
	wire _04583_;
	wire _04584_;
	wire _04585_;
	wire _04586_;
	wire _04587_;
	wire _04588_;
	wire _04589_;
	wire _04590_;
	wire _04591_;
	wire _04592_;
	wire _04593_;
	wire _04594_;
	wire _04595_;
	wire _04596_;
	wire _04597_;
	wire _04598_;
	wire _04599_;
	wire _04600_;
	wire _04601_;
	wire _04602_;
	wire _04603_;
	wire _04604_;
	wire _04605_;
	wire _04606_;
	wire _04607_;
	wire _04608_;
	wire _04609_;
	wire _04610_;
	wire _04611_;
	wire _04612_;
	wire _04613_;
	wire _04614_;
	wire _04615_;
	wire _04616_;
	wire _04617_;
	wire _04618_;
	wire _04619_;
	wire _04620_;
	wire _04621_;
	wire _04622_;
	wire _04623_;
	wire _04624_;
	wire _04625_;
	wire _04626_;
	wire _04627_;
	wire _04628_;
	wire _04629_;
	wire _04630_;
	wire _04631_;
	wire _04632_;
	wire _04633_;
	wire _04634_;
	wire _04635_;
	wire _04636_;
	wire _04637_;
	wire _04638_;
	wire _04639_;
	wire _04640_;
	wire _04641_;
	wire _04642_;
	wire _04643_;
	wire _04644_;
	wire _04645_;
	wire _04646_;
	wire _04647_;
	wire _04648_;
	wire _04649_;
	wire _04650_;
	wire _04651_;
	wire _04652_;
	wire _04653_;
	wire _04654_;
	wire _04655_;
	wire _04656_;
	wire _04657_;
	wire _04658_;
	wire _04659_;
	wire _04660_;
	wire _04661_;
	wire _04662_;
	wire _04663_;
	wire _04664_;
	wire _04665_;
	wire _04666_;
	wire _04667_;
	wire _04668_;
	wire _04669_;
	wire _04670_;
	wire _04671_;
	wire _04672_;
	wire _04673_;
	wire _04674_;
	wire _04675_;
	wire _04676_;
	wire _04677_;
	wire _04678_;
	wire _04679_;
	wire _04680_;
	wire _04681_;
	wire _04682_;
	wire _04683_;
	wire _04684_;
	wire _04685_;
	wire _04686_;
	wire _04687_;
	wire _04688_;
	wire _04689_;
	wire _04690_;
	wire _04691_;
	wire _04692_;
	wire _04693_;
	wire _04694_;
	wire _04695_;
	wire _04696_;
	wire _04697_;
	wire _04698_;
	wire _04699_;
	wire _04700_;
	wire _04701_;
	wire _04702_;
	wire _04703_;
	wire _04704_;
	wire _04705_;
	wire _04706_;
	wire _04707_;
	wire _04708_;
	wire _04709_;
	wire _04710_;
	wire _04711_;
	wire _04712_;
	wire _04713_;
	wire _04714_;
	wire _04715_;
	wire _04716_;
	wire _04717_;
	wire _04718_;
	wire _04719_;
	wire _04720_;
	wire _04721_;
	wire _04722_;
	wire _04723_;
	wire _04724_;
	wire _04725_;
	wire _04726_;
	wire _04727_;
	wire _04728_;
	wire _04729_;
	wire _04730_;
	wire _04731_;
	wire _04732_;
	wire _04733_;
	wire _04734_;
	wire _04735_;
	wire _04736_;
	wire _04737_;
	wire _04738_;
	wire _04739_;
	wire _04740_;
	wire _04741_;
	wire _04742_;
	wire _04743_;
	wire _04744_;
	wire _04745_;
	wire _04746_;
	wire _04747_;
	wire _04748_;
	wire _04749_;
	wire _04750_;
	wire _04751_;
	wire _04752_;
	wire _04753_;
	wire _04754_;
	wire _04755_;
	wire _04756_;
	wire _04757_;
	wire _04758_;
	wire _04759_;
	wire _04760_;
	wire _04761_;
	wire _04762_;
	wire _04763_;
	wire _04764_;
	wire _04765_;
	wire _04766_;
	wire _04767_;
	wire _04768_;
	wire _04769_;
	wire _04770_;
	wire _04771_;
	wire _04772_;
	wire _04773_;
	wire _04774_;
	wire _04775_;
	wire _04776_;
	wire _04777_;
	wire _04778_;
	wire _04779_;
	wire _04780_;
	wire _04781_;
	wire _04782_;
	wire _04783_;
	wire _04784_;
	wire _04785_;
	wire _04786_;
	wire _04787_;
	wire _04788_;
	wire _04789_;
	wire _04790_;
	wire _04791_;
	wire _04792_;
	wire _04793_;
	wire _04794_;
	wire _04795_;
	wire _04796_;
	wire _04797_;
	wire _04798_;
	wire _04799_;
	wire _04800_;
	wire _04801_;
	wire _04802_;
	wire _04803_;
	wire _04804_;
	wire _04805_;
	wire _04806_;
	wire _04807_;
	wire _04808_;
	wire _04809_;
	wire _04810_;
	wire _04811_;
	wire _04812_;
	wire _04813_;
	wire _04814_;
	wire _04815_;
	wire _04816_;
	wire _04817_;
	wire _04818_;
	wire _04819_;
	wire _04820_;
	wire _04821_;
	wire _04822_;
	wire _04823_;
	wire _04824_;
	wire _04825_;
	wire _04826_;
	wire _04827_;
	wire _04828_;
	wire _04829_;
	wire _04830_;
	wire _04831_;
	wire _04832_;
	wire _04833_;
	wire _04834_;
	wire _04835_;
	wire _04836_;
	wire _04837_;
	wire _04838_;
	wire _04839_;
	wire _04840_;
	wire _04841_;
	wire _04842_;
	wire _04843_;
	wire _04844_;
	wire _04845_;
	wire _04846_;
	wire _04847_;
	wire _04848_;
	wire _04849_;
	wire _04850_;
	wire _04851_;
	wire _04852_;
	wire _04853_;
	wire _04854_;
	wire _04855_;
	wire _04856_;
	wire _04857_;
	wire _04858_;
	wire _04859_;
	wire _04860_;
	wire _04861_;
	wire _04862_;
	wire _04863_;
	wire _04864_;
	wire _04865_;
	wire _04866_;
	wire _04867_;
	wire _04868_;
	wire _04869_;
	wire _04870_;
	wire _04871_;
	wire _04872_;
	wire _04873_;
	wire _04874_;
	wire _04875_;
	wire _04876_;
	wire _04877_;
	wire _04878_;
	wire _04879_;
	wire _04880_;
	wire _04881_;
	wire _04882_;
	wire _04883_;
	wire _04884_;
	wire _04885_;
	wire _04886_;
	wire _04887_;
	wire _04888_;
	wire _04889_;
	wire _04890_;
	wire _04891_;
	wire _04892_;
	wire _04893_;
	wire _04894_;
	wire _04895_;
	wire _04896_;
	wire _04897_;
	wire _04898_;
	wire _04899_;
	wire _04900_;
	wire _04901_;
	wire _04902_;
	wire _04903_;
	wire _04904_;
	wire _04905_;
	wire _04906_;
	wire _04907_;
	wire _04908_;
	wire _04909_;
	wire _04910_;
	wire _04911_;
	wire _04912_;
	wire _04913_;
	wire _04914_;
	wire _04915_;
	wire _04916_;
	wire _04917_;
	wire _04918_;
	wire _04919_;
	wire _04920_;
	wire _04921_;
	wire _04922_;
	wire _04923_;
	wire _04924_;
	wire _04925_;
	wire _04926_;
	wire _04927_;
	wire _04928_;
	wire _04929_;
	wire _04930_;
	wire _04931_;
	wire _04932_;
	wire _04933_;
	wire _04934_;
	wire _04935_;
	wire _04936_;
	wire _04937_;
	wire _04938_;
	wire _04939_;
	wire _04940_;
	wire _04941_;
	wire _04942_;
	wire _04943_;
	wire _04944_;
	wire _04945_;
	wire _04946_;
	wire _04947_;
	wire _04948_;
	wire _04949_;
	wire _04950_;
	wire _04951_;
	wire _04952_;
	wire _04953_;
	wire _04954_;
	wire _04955_;
	wire _04956_;
	wire _04957_;
	wire _04958_;
	wire _04959_;
	wire _04960_;
	wire _04961_;
	wire _04962_;
	wire _04963_;
	wire _04964_;
	wire _04965_;
	wire _04966_;
	wire _04967_;
	wire _04968_;
	wire _04969_;
	wire _04970_;
	wire _04971_;
	wire _04972_;
	wire _04973_;
	wire _04974_;
	wire _04975_;
	wire _04976_;
	wire _04977_;
	wire _04978_;
	wire _04979_;
	wire _04980_;
	wire _04981_;
	wire _04982_;
	wire _04983_;
	wire _04984_;
	wire _04985_;
	wire _04986_;
	wire _04987_;
	wire _04988_;
	wire _04989_;
	wire _04990_;
	wire _04991_;
	wire _04992_;
	wire _04993_;
	wire _04994_;
	wire _04995_;
	wire _04996_;
	wire _04997_;
	wire _04998_;
	wire _04999_;
	wire _05000_;
	wire _05001_;
	wire _05002_;
	wire _05003_;
	wire _05004_;
	wire _05005_;
	wire _05006_;
	wire _05007_;
	wire _05008_;
	wire _05009_;
	wire _05010_;
	wire _05011_;
	wire _05012_;
	wire _05013_;
	wire _05014_;
	wire _05015_;
	wire _05016_;
	wire _05017_;
	wire _05018_;
	wire _05019_;
	wire _05020_;
	wire _05021_;
	wire _05022_;
	wire _05023_;
	wire _05024_;
	wire _05025_;
	wire _05026_;
	wire _05027_;
	wire _05028_;
	wire _05029_;
	wire _05030_;
	wire _05031_;
	wire _05032_;
	wire _05033_;
	wire _05034_;
	wire _05035_;
	wire _05036_;
	wire _05037_;
	wire _05038_;
	wire _05039_;
	wire _05040_;
	wire _05041_;
	wire _05042_;
	wire _05043_;
	wire _05044_;
	wire _05045_;
	wire _05046_;
	wire _05047_;
	wire _05048_;
	wire _05049_;
	wire _05050_;
	wire _05051_;
	wire _05052_;
	wire _05053_;
	wire _05054_;
	wire _05055_;
	wire _05056_;
	wire _05057_;
	wire _05058_;
	wire _05059_;
	wire _05060_;
	wire _05061_;
	wire _05062_;
	wire _05063_;
	wire _05064_;
	wire _05065_;
	wire _05066_;
	wire _05067_;
	wire _05068_;
	wire _05069_;
	wire _05070_;
	wire _05071_;
	wire _05072_;
	wire _05073_;
	wire _05074_;
	wire _05075_;
	wire _05076_;
	wire _05077_;
	wire _05078_;
	wire _05079_;
	wire _05080_;
	wire _05081_;
	wire _05082_;
	wire _05083_;
	wire _05084_;
	wire _05085_;
	wire _05086_;
	wire _05087_;
	wire _05088_;
	wire _05089_;
	wire _05090_;
	wire _05091_;
	wire _05092_;
	wire _05093_;
	wire _05094_;
	wire _05095_;
	wire _05096_;
	wire _05097_;
	wire _05098_;
	wire _05099_;
	wire _05100_;
	wire _05101_;
	wire _05102_;
	wire _05103_;
	wire _05104_;
	wire _05105_;
	wire _05106_;
	wire _05107_;
	wire _05108_;
	wire _05109_;
	wire _05110_;
	wire _05111_;
	wire _05112_;
	wire _05113_;
	wire _05114_;
	wire _05115_;
	wire _05116_;
	wire _05117_;
	wire _05118_;
	wire _05119_;
	wire _05120_;
	wire _05121_;
	wire _05122_;
	wire _05123_;
	wire _05124_;
	wire _05125_;
	wire _05126_;
	wire _05127_;
	wire _05128_;
	wire _05129_;
	wire _05130_;
	wire _05131_;
	wire _05132_;
	wire _05133_;
	wire _05134_;
	wire _05135_;
	wire _05136_;
	wire _05137_;
	wire _05138_;
	wire _05139_;
	wire _05140_;
	wire _05141_;
	wire _05142_;
	wire _05143_;
	wire _05144_;
	wire _05145_;
	wire _05146_;
	wire _05147_;
	wire _05148_;
	wire _05149_;
	wire _05150_;
	wire _05151_;
	wire _05152_;
	wire _05153_;
	wire _05154_;
	wire _05155_;
	wire _05156_;
	wire _05157_;
	wire _05158_;
	wire _05159_;
	wire _05160_;
	wire _05161_;
	wire _05162_;
	wire _05163_;
	wire _05164_;
	wire _05165_;
	wire _05166_;
	wire _05167_;
	wire _05168_;
	wire _05169_;
	wire _05170_;
	wire _05171_;
	wire _05172_;
	wire _05173_;
	wire _05174_;
	wire _05175_;
	wire _05176_;
	wire _05177_;
	wire _05178_;
	wire _05179_;
	wire _05180_;
	wire _05181_;
	wire _05182_;
	wire _05183_;
	wire _05184_;
	wire _05185_;
	wire _05186_;
	wire _05187_;
	wire _05188_;
	wire _05189_;
	wire _05190_;
	wire _05191_;
	wire _05192_;
	wire _05193_;
	wire _05194_;
	wire _05195_;
	wire _05196_;
	wire _05197_;
	wire _05198_;
	wire _05199_;
	wire _05200_;
	wire _05201_;
	wire _05202_;
	wire _05203_;
	wire _05204_;
	wire _05205_;
	wire _05206_;
	wire _05207_;
	wire _05208_;
	wire _05209_;
	wire _05210_;
	wire _05211_;
	wire _05212_;
	wire _05213_;
	wire _05214_;
	wire _05215_;
	wire _05216_;
	wire _05217_;
	wire _05218_;
	wire _05219_;
	wire _05220_;
	wire _05221_;
	wire _05222_;
	wire _05223_;
	wire _05224_;
	wire _05225_;
	wire _05226_;
	wire _05227_;
	wire _05228_;
	wire _05229_;
	wire _05230_;
	wire _05231_;
	wire _05232_;
	wire _05233_;
	wire _05234_;
	wire _05235_;
	wire _05236_;
	wire _05237_;
	wire _05238_;
	wire _05239_;
	wire _05240_;
	wire _05241_;
	wire _05242_;
	wire _05243_;
	wire _05244_;
	wire _05245_;
	wire _05246_;
	wire _05247_;
	wire _05248_;
	wire _05249_;
	wire _05250_;
	wire _05251_;
	wire _05252_;
	wire _05253_;
	wire _05254_;
	wire _05255_;
	wire _05256_;
	wire _05257_;
	wire _05258_;
	wire _05259_;
	wire _05260_;
	wire _05261_;
	wire _05262_;
	wire _05263_;
	wire _05264_;
	wire _05265_;
	wire _05266_;
	wire _05267_;
	wire _05268_;
	wire _05269_;
	wire _05270_;
	wire _05271_;
	wire _05272_;
	wire _05273_;
	wire _05274_;
	wire _05275_;
	wire _05276_;
	wire _05277_;
	wire _05278_;
	wire _05279_;
	wire _05280_;
	wire _05281_;
	wire _05282_;
	wire _05283_;
	wire _05284_;
	wire _05285_;
	wire _05286_;
	wire _05287_;
	wire _05288_;
	wire _05289_;
	wire _05290_;
	wire _05291_;
	wire _05292_;
	wire _05293_;
	wire _05294_;
	wire _05295_;
	wire _05296_;
	wire _05297_;
	wire _05298_;
	wire _05299_;
	wire _05300_;
	wire _05301_;
	wire _05302_;
	wire _05303_;
	wire _05304_;
	wire _05305_;
	wire _05306_;
	wire _05307_;
	wire _05308_;
	wire _05309_;
	wire _05310_;
	wire _05311_;
	wire _05312_;
	wire _05313_;
	wire _05314_;
	wire _05315_;
	wire _05316_;
	wire _05317_;
	wire _05318_;
	wire _05319_;
	wire _05320_;
	wire _05321_;
	wire _05322_;
	wire _05323_;
	wire _05324_;
	wire _05325_;
	wire _05326_;
	wire _05327_;
	wire _05328_;
	wire _05329_;
	wire _05330_;
	wire _05331_;
	wire _05332_;
	wire _05333_;
	wire _05334_;
	wire _05335_;
	wire _05336_;
	wire _05337_;
	wire _05338_;
	wire _05339_;
	wire _05340_;
	wire _05341_;
	wire _05342_;
	wire _05343_;
	wire _05344_;
	wire _05345_;
	wire _05346_;
	wire _05347_;
	wire _05348_;
	wire _05349_;
	wire _05350_;
	wire _05351_;
	wire _05352_;
	wire _05353_;
	wire _05354_;
	wire _05355_;
	wire _05356_;
	wire _05357_;
	wire _05358_;
	wire _05359_;
	wire _05360_;
	wire _05361_;
	wire _05362_;
	wire _05363_;
	wire _05364_;
	wire _05365_;
	wire _05366_;
	wire _05367_;
	wire _05368_;
	wire _05369_;
	wire _05370_;
	wire _05371_;
	wire _05372_;
	wire _05373_;
	wire _05374_;
	wire _05375_;
	wire _05376_;
	wire _05377_;
	wire _05378_;
	wire _05379_;
	wire _05380_;
	wire _05381_;
	wire _05382_;
	wire _05383_;
	wire _05384_;
	wire _05385_;
	wire _05386_;
	wire _05387_;
	wire _05388_;
	wire _05389_;
	wire _05390_;
	wire _05391_;
	wire _05392_;
	wire _05393_;
	wire _05394_;
	wire _05395_;
	wire _05396_;
	wire _05397_;
	wire _05398_;
	wire _05399_;
	wire _05400_;
	wire _05401_;
	wire _05402_;
	wire _05403_;
	wire _05404_;
	wire _05405_;
	wire _05406_;
	wire _05407_;
	wire _05408_;
	wire _05409_;
	wire _05410_;
	wire _05411_;
	wire _05412_;
	wire _05413_;
	wire _05414_;
	wire _05415_;
	wire _05416_;
	wire _05417_;
	wire _05418_;
	wire _05419_;
	wire _05420_;
	wire _05421_;
	wire _05422_;
	wire _05423_;
	wire _05424_;
	wire _05425_;
	wire _05426_;
	wire _05427_;
	wire _05428_;
	wire _05429_;
	wire _05430_;
	wire _05431_;
	wire _05432_;
	wire _05433_;
	wire _05434_;
	wire _05435_;
	wire _05436_;
	wire _05437_;
	wire _05438_;
	wire _05439_;
	wire _05440_;
	wire _05441_;
	wire _05442_;
	wire _05443_;
	wire _05444_;
	wire _05445_;
	wire _05446_;
	wire _05447_;
	wire _05448_;
	wire _05449_;
	wire _05450_;
	wire _05451_;
	wire _05452_;
	wire _05453_;
	wire _05454_;
	wire _05455_;
	wire _05456_;
	wire _05457_;
	wire _05458_;
	wire _05459_;
	wire _05460_;
	wire _05461_;
	wire _05462_;
	wire _05463_;
	wire _05464_;
	wire _05465_;
	wire _05466_;
	wire _05467_;
	wire _05468_;
	wire _05469_;
	wire _05470_;
	wire _05471_;
	wire _05472_;
	wire _05473_;
	wire _05474_;
	wire _05475_;
	wire _05476_;
	wire _05477_;
	wire _05478_;
	wire _05479_;
	wire _05480_;
	wire _05481_;
	wire _05482_;
	wire _05483_;
	wire _05484_;
	wire _05485_;
	wire _05486_;
	wire _05487_;
	wire _05488_;
	wire _05489_;
	wire _05490_;
	wire _05491_;
	wire _05492_;
	wire _05493_;
	wire _05494_;
	wire _05495_;
	wire _05496_;
	wire _05497_;
	wire _05498_;
	wire _05499_;
	wire _05500_;
	wire _05501_;
	wire _05502_;
	wire _05503_;
	wire _05504_;
	wire _05505_;
	wire _05506_;
	wire _05507_;
	wire _05508_;
	wire _05509_;
	wire _05510_;
	wire _05511_;
	wire _05512_;
	wire _05513_;
	wire _05514_;
	wire _05515_;
	wire _05516_;
	wire _05517_;
	wire _05518_;
	wire _05519_;
	wire _05520_;
	wire _05521_;
	wire _05522_;
	wire _05523_;
	wire _05524_;
	wire _05525_;
	wire _05526_;
	wire _05527_;
	wire _05528_;
	wire _05529_;
	wire _05530_;
	wire _05531_;
	wire _05532_;
	wire _05533_;
	wire _05534_;
	wire _05535_;
	wire _05536_;
	wire _05537_;
	wire _05538_;
	wire _05539_;
	wire _05540_;
	wire _05541_;
	wire _05542_;
	wire _05543_;
	wire _05544_;
	wire _05545_;
	wire _05546_;
	wire _05547_;
	wire _05548_;
	wire _05549_;
	wire _05550_;
	wire _05551_;
	wire _05552_;
	wire _05553_;
	wire _05554_;
	wire _05555_;
	wire _05556_;
	wire _05557_;
	wire _05558_;
	wire _05559_;
	wire _05560_;
	wire _05561_;
	wire _05562_;
	wire _05563_;
	wire _05564_;
	wire _05565_;
	wire _05566_;
	wire _05567_;
	wire _05568_;
	wire _05569_;
	wire _05570_;
	wire _05571_;
	wire _05572_;
	wire _05573_;
	wire _05574_;
	wire _05575_;
	wire _05576_;
	wire _05577_;
	wire _05578_;
	wire _05579_;
	wire _05580_;
	wire _05581_;
	wire _05582_;
	wire _05583_;
	wire _05584_;
	wire _05585_;
	wire _05586_;
	wire _05587_;
	wire _05588_;
	wire _05589_;
	wire _05590_;
	wire _05591_;
	wire _05592_;
	wire _05593_;
	wire _05594_;
	wire _05595_;
	wire _05596_;
	wire _05597_;
	wire _05598_;
	wire _05599_;
	wire _05600_;
	wire _05601_;
	wire _05602_;
	wire _05603_;
	wire _05604_;
	wire _05605_;
	wire _05606_;
	wire _05607_;
	wire _05608_;
	wire _05609_;
	wire _05610_;
	wire _05611_;
	wire _05612_;
	wire _05613_;
	wire _05614_;
	wire _05615_;
	wire _05616_;
	wire _05617_;
	wire _05618_;
	wire _05619_;
	wire _05620_;
	wire _05621_;
	wire _05622_;
	wire _05623_;
	wire _05624_;
	wire _05625_;
	wire _05626_;
	wire _05627_;
	wire _05628_;
	wire _05629_;
	wire _05630_;
	wire _05631_;
	wire _05632_;
	wire _05633_;
	wire _05634_;
	wire _05635_;
	wire _05636_;
	wire _05637_;
	wire _05638_;
	wire _05639_;
	wire _05640_;
	wire _05641_;
	wire _05642_;
	wire _05643_;
	wire _05644_;
	wire _05645_;
	wire _05646_;
	wire _05647_;
	wire _05648_;
	wire _05649_;
	wire _05650_;
	wire _05651_;
	wire _05652_;
	wire _05653_;
	wire _05654_;
	wire _05655_;
	wire _05656_;
	wire _05657_;
	wire _05658_;
	wire _05659_;
	wire _05660_;
	wire _05661_;
	wire _05662_;
	wire _05663_;
	wire _05664_;
	wire _05665_;
	wire _05666_;
	wire _05667_;
	wire _05668_;
	wire _05669_;
	wire _05670_;
	wire _05671_;
	wire _05672_;
	wire _05673_;
	wire _05674_;
	wire _05675_;
	wire _05676_;
	wire _05677_;
	wire _05678_;
	wire _05679_;
	wire _05680_;
	wire _05681_;
	wire _05682_;
	wire _05683_;
	wire _05684_;
	wire _05685_;
	wire _05686_;
	wire _05687_;
	wire _05688_;
	wire _05689_;
	wire _05690_;
	wire _05691_;
	wire _05692_;
	wire _05693_;
	wire _05694_;
	wire _05695_;
	wire _05696_;
	wire _05697_;
	wire _05698_;
	wire _05699_;
	wire _05700_;
	wire _05701_;
	wire _05702_;
	wire _05703_;
	wire _05704_;
	wire _05705_;
	wire _05706_;
	wire _05707_;
	wire _05708_;
	wire _05709_;
	wire _05710_;
	wire _05711_;
	wire _05712_;
	wire _05713_;
	wire _05714_;
	wire _05715_;
	wire _05716_;
	wire _05717_;
	wire _05718_;
	wire _05719_;
	wire _05720_;
	wire _05721_;
	wire _05722_;
	wire _05723_;
	wire _05724_;
	wire _05725_;
	wire _05726_;
	wire _05727_;
	wire _05728_;
	wire _05729_;
	wire _05730_;
	wire _05731_;
	wire _05732_;
	wire _05733_;
	wire _05734_;
	wire _05735_;
	wire _05736_;
	wire _05737_;
	wire _05738_;
	wire _05739_;
	wire _05740_;
	wire _05741_;
	wire _05742_;
	wire _05743_;
	wire _05744_;
	wire _05745_;
	wire _05746_;
	wire _05747_;
	wire _05748_;
	wire _05749_;
	wire _05750_;
	wire _05751_;
	wire _05752_;
	wire _05753_;
	wire _05754_;
	wire _05755_;
	wire _05756_;
	wire _05757_;
	wire _05758_;
	wire _05759_;
	wire _05760_;
	wire _05761_;
	wire _05762_;
	wire _05763_;
	wire _05764_;
	wire _05765_;
	wire _05766_;
	wire _05767_;
	wire _05768_;
	wire _05769_;
	wire _05770_;
	wire _05771_;
	wire _05772_;
	wire _05773_;
	wire _05774_;
	wire _05775_;
	wire _05776_;
	wire _05777_;
	wire _05778_;
	wire _05779_;
	wire _05780_;
	wire _05781_;
	wire _05782_;
	wire _05783_;
	wire _05784_;
	wire _05785_;
	wire _05786_;
	wire _05787_;
	wire _05788_;
	wire _05789_;
	wire _05790_;
	wire _05791_;
	wire _05792_;
	wire _05793_;
	wire _05794_;
	wire _05795_;
	wire _05796_;
	wire _05797_;
	wire _05798_;
	wire _05799_;
	wire _05800_;
	wire _05801_;
	wire _05802_;
	wire _05803_;
	wire _05804_;
	wire _05805_;
	wire _05806_;
	wire _05807_;
	wire _05808_;
	wire _05809_;
	wire _05810_;
	wire _05811_;
	wire _05812_;
	wire _05813_;
	wire _05814_;
	wire _05815_;
	wire _05816_;
	wire _05817_;
	wire _05818_;
	wire _05819_;
	wire _05820_;
	wire _05821_;
	wire _05822_;
	wire _05823_;
	wire _05824_;
	wire _05825_;
	wire _05826_;
	wire _05827_;
	wire _05828_;
	wire _05829_;
	wire _05830_;
	wire _05831_;
	wire _05832_;
	wire _05833_;
	wire _05834_;
	wire _05835_;
	wire _05836_;
	wire _05837_;
	wire _05838_;
	wire _05839_;
	wire _05840_;
	wire _05841_;
	wire _05842_;
	wire _05843_;
	wire _05844_;
	wire _05845_;
	wire _05846_;
	wire _05847_;
	wire _05848_;
	wire _05849_;
	wire _05850_;
	wire _05851_;
	wire _05852_;
	wire _05853_;
	wire _05854_;
	wire _05855_;
	wire _05856_;
	wire _05857_;
	wire _05858_;
	wire _05859_;
	wire _05860_;
	wire _05861_;
	wire _05862_;
	wire _05863_;
	wire _05864_;
	wire _05865_;
	wire _05866_;
	wire _05867_;
	wire _05868_;
	wire _05869_;
	wire _05870_;
	wire _05871_;
	wire _05872_;
	wire _05873_;
	wire _05874_;
	wire _05875_;
	wire _05876_;
	wire _05877_;
	wire _05878_;
	wire _05879_;
	wire _05880_;
	wire _05881_;
	wire _05882_;
	wire _05883_;
	wire _05884_;
	wire _05885_;
	wire _05886_;
	wire _05887_;
	wire _05888_;
	wire _05889_;
	wire _05890_;
	wire _05891_;
	wire _05892_;
	wire _05893_;
	wire _05894_;
	wire _05895_;
	wire _05896_;
	wire _05897_;
	wire _05898_;
	wire _05899_;
	wire _05900_;
	wire _05901_;
	wire _05902_;
	wire _05903_;
	wire _05904_;
	wire _05905_;
	wire _05906_;
	wire _05907_;
	wire _05908_;
	wire _05909_;
	wire _05910_;
	wire _05911_;
	wire _05912_;
	wire _05913_;
	wire _05914_;
	wire _05915_;
	wire _05916_;
	wire _05917_;
	wire _05918_;
	wire _05919_;
	wire _05920_;
	wire _05921_;
	wire _05922_;
	wire _05923_;
	wire _05924_;
	wire _05925_;
	wire _05926_;
	wire _05927_;
	wire _05928_;
	wire _05929_;
	wire _05930_;
	wire _05931_;
	wire _05932_;
	wire _05933_;
	wire _05934_;
	wire _05935_;
	wire _05936_;
	wire _05937_;
	wire _05938_;
	wire _05939_;
	wire _05940_;
	wire _05941_;
	wire _05942_;
	wire _05943_;
	wire _05944_;
	wire _05945_;
	wire _05946_;
	wire _05947_;
	wire _05948_;
	wire _05949_;
	wire _05950_;
	wire _05951_;
	wire _05952_;
	wire _05953_;
	wire _05954_;
	wire _05955_;
	wire _05956_;
	wire _05957_;
	wire _05958_;
	wire _05959_;
	wire _05960_;
	wire _05961_;
	wire _05962_;
	wire _05963_;
	wire _05964_;
	wire _05965_;
	wire _05966_;
	wire _05967_;
	wire _05968_;
	wire _05969_;
	wire _05970_;
	wire _05971_;
	wire _05972_;
	wire _05973_;
	wire _05974_;
	wire _05975_;
	wire _05976_;
	wire _05977_;
	wire _05978_;
	wire _05979_;
	wire _05980_;
	wire _05981_;
	wire _05982_;
	wire _05983_;
	wire _05984_;
	wire _05985_;
	wire _05986_;
	wire _05987_;
	wire _05988_;
	wire _05989_;
	wire _05990_;
	wire _05991_;
	wire _05992_;
	wire _05993_;
	wire _05994_;
	wire _05995_;
	wire _05996_;
	wire _05997_;
	wire _05998_;
	wire _05999_;
	wire _06000_;
	wire _06001_;
	wire _06002_;
	wire _06003_;
	wire _06004_;
	wire _06005_;
	wire _06006_;
	wire _06007_;
	wire _06008_;
	wire _06009_;
	wire _06010_;
	wire _06011_;
	wire _06012_;
	wire _06013_;
	wire _06014_;
	wire _06015_;
	wire _06016_;
	wire _06017_;
	wire _06018_;
	wire _06019_;
	wire _06020_;
	wire _06021_;
	wire _06022_;
	wire _06023_;
	wire _06024_;
	wire _06025_;
	wire _06026_;
	wire _06027_;
	wire _06028_;
	wire _06029_;
	wire _06030_;
	wire _06031_;
	wire _06032_;
	wire _06033_;
	wire _06034_;
	wire _06035_;
	wire _06036_;
	wire _06037_;
	wire _06038_;
	wire _06039_;
	wire _06040_;
	wire _06041_;
	wire _06042_;
	wire _06043_;
	wire _06044_;
	wire _06045_;
	wire _06046_;
	wire _06047_;
	wire _06048_;
	wire _06049_;
	wire _06050_;
	wire _06051_;
	wire _06052_;
	wire _06053_;
	wire _06054_;
	wire _06055_;
	wire _06056_;
	wire _06057_;
	wire _06058_;
	wire _06059_;
	wire _06060_;
	wire _06061_;
	wire _06062_;
	wire _06063_;
	wire _06064_;
	wire _06065_;
	wire _06066_;
	wire _06067_;
	wire _06068_;
	wire _06069_;
	wire _06070_;
	wire _06071_;
	wire _06072_;
	wire _06073_;
	wire _06074_;
	wire _06075_;
	wire _06076_;
	wire _06077_;
	wire _06078_;
	wire _06079_;
	wire _06080_;
	wire _06081_;
	wire _06082_;
	wire _06083_;
	wire _06084_;
	wire _06085_;
	wire _06086_;
	wire _06087_;
	wire _06088_;
	wire _06089_;
	wire _06090_;
	wire _06091_;
	wire _06092_;
	wire _06093_;
	wire _06094_;
	wire _06095_;
	wire _06096_;
	wire _06097_;
	wire _06098_;
	wire _06099_;
	wire _06100_;
	wire _06101_;
	wire _06102_;
	wire _06103_;
	wire _06104_;
	wire _06105_;
	wire _06106_;
	wire _06107_;
	wire _06108_;
	wire _06109_;
	wire _06110_;
	wire _06111_;
	wire _06112_;
	wire _06113_;
	wire _06114_;
	wire _06115_;
	wire _06116_;
	wire _06117_;
	wire _06118_;
	wire _06119_;
	wire _06120_;
	wire _06121_;
	wire _06122_;
	wire _06123_;
	wire _06124_;
	wire _06125_;
	wire _06126_;
	wire _06127_;
	wire _06128_;
	wire _06129_;
	wire _06130_;
	wire _06131_;
	wire _06132_;
	wire _06133_;
	wire _06134_;
	wire _06135_;
	wire _06136_;
	wire _06137_;
	wire _06138_;
	wire _06139_;
	wire _06140_;
	wire _06141_;
	wire _06142_;
	wire _06143_;
	wire _06144_;
	wire _06145_;
	wire _06146_;
	wire _06147_;
	wire _06148_;
	wire _06149_;
	wire _06150_;
	wire _06151_;
	wire _06152_;
	wire _06153_;
	wire _06154_;
	wire _06155_;
	wire _06156_;
	wire _06157_;
	wire _06158_;
	wire _06159_;
	wire _06160_;
	wire _06161_;
	wire _06162_;
	wire _06163_;
	wire _06164_;
	wire _06165_;
	wire _06166_;
	wire _06167_;
	wire _06168_;
	wire _06169_;
	wire _06170_;
	wire _06171_;
	wire _06172_;
	wire _06173_;
	wire _06174_;
	wire _06175_;
	wire _06176_;
	wire _06177_;
	wire _06178_;
	wire _06179_;
	wire _06180_;
	wire _06181_;
	wire _06182_;
	wire _06183_;
	wire _06184_;
	wire _06185_;
	wire _06186_;
	wire _06187_;
	wire _06188_;
	wire _06189_;
	wire _06190_;
	wire _06191_;
	wire _06192_;
	wire _06193_;
	wire _06194_;
	wire _06195_;
	wire _06196_;
	wire _06197_;
	wire _06198_;
	wire _06199_;
	wire _06200_;
	wire _06201_;
	wire _06202_;
	wire _06203_;
	wire _06204_;
	wire _06205_;
	wire _06206_;
	wire _06207_;
	wire _06208_;
	wire _06209_;
	wire _06210_;
	wire _06211_;
	wire _06212_;
	wire _06213_;
	wire _06214_;
	wire _06215_;
	wire _06216_;
	wire _06217_;
	wire _06218_;
	wire _06219_;
	wire _06220_;
	wire _06221_;
	wire _06222_;
	wire _06223_;
	wire _06224_;
	wire _06225_;
	wire _06226_;
	wire _06227_;
	wire _06228_;
	wire _06229_;
	wire _06230_;
	wire _06231_;
	wire _06232_;
	wire _06233_;
	wire _06234_;
	wire _06235_;
	wire _06236_;
	wire _06237_;
	wire _06238_;
	wire _06239_;
	wire _06240_;
	wire _06241_;
	wire _06242_;
	wire _06243_;
	wire _06244_;
	wire _06245_;
	wire _06246_;
	wire _06247_;
	wire _06248_;
	wire _06249_;
	wire _06250_;
	wire _06251_;
	wire _06252_;
	wire _06253_;
	wire _06254_;
	wire _06255_;
	wire _06256_;
	wire _06257_;
	wire _06258_;
	wire _06259_;
	wire _06260_;
	wire _06261_;
	wire _06262_;
	wire _06263_;
	wire _06264_;
	wire _06265_;
	wire _06266_;
	wire _06267_;
	wire _06268_;
	wire _06269_;
	wire _06270_;
	wire _06271_;
	wire _06272_;
	wire _06273_;
	wire _06274_;
	wire _06275_;
	wire _06276_;
	wire _06277_;
	wire _06278_;
	wire _06279_;
	wire _06280_;
	wire _06281_;
	wire _06282_;
	wire _06283_;
	wire _06284_;
	wire _06285_;
	wire _06286_;
	wire _06287_;
	wire _06288_;
	wire _06289_;
	wire _06290_;
	wire _06291_;
	wire _06292_;
	wire _06293_;
	wire _06294_;
	wire _06295_;
	wire _06296_;
	wire _06297_;
	wire _06298_;
	wire _06299_;
	wire _06300_;
	wire _06301_;
	wire _06302_;
	wire _06303_;
	wire _06304_;
	wire _06305_;
	wire _06306_;
	wire _06307_;
	wire _06308_;
	wire _06309_;
	wire _06310_;
	wire _06311_;
	wire _06312_;
	wire _06313_;
	wire _06314_;
	wire _06315_;
	wire _06316_;
	wire _06317_;
	wire _06318_;
	wire _06319_;
	wire _06320_;
	wire _06321_;
	wire _06322_;
	wire _06323_;
	wire _06324_;
	wire _06325_;
	wire _06326_;
	wire _06327_;
	wire _06328_;
	wire _06329_;
	wire _06330_;
	wire _06331_;
	wire _06332_;
	wire _06333_;
	wire _06334_;
	wire _06335_;
	wire _06336_;
	wire _06337_;
	wire _06338_;
	wire _06339_;
	wire _06340_;
	wire _06341_;
	wire _06342_;
	wire _06343_;
	wire _06344_;
	wire _06345_;
	wire _06346_;
	wire _06347_;
	wire _06348_;
	wire _06349_;
	wire _06350_;
	wire _06351_;
	wire _06352_;
	wire _06353_;
	wire _06354_;
	wire _06355_;
	wire _06356_;
	wire _06357_;
	wire _06358_;
	wire _06359_;
	wire _06360_;
	wire _06361_;
	wire _06362_;
	wire _06363_;
	wire _06364_;
	wire _06365_;
	wire _06366_;
	wire _06367_;
	wire _06368_;
	wire _06369_;
	wire _06370_;
	wire _06371_;
	wire _06372_;
	wire _06373_;
	wire _06374_;
	wire _06375_;
	wire _06376_;
	wire _06377_;
	wire _06378_;
	wire _06379_;
	wire _06380_;
	wire _06381_;
	wire _06382_;
	wire _06383_;
	wire _06384_;
	wire _06385_;
	wire _06386_;
	wire _06387_;
	wire _06388_;
	wire _06389_;
	wire _06390_;
	wire _06391_;
	wire _06392_;
	wire _06393_;
	wire _06394_;
	wire _06395_;
	wire _06396_;
	wire _06397_;
	wire _06398_;
	wire _06399_;
	wire _06400_;
	wire _06401_;
	wire _06402_;
	wire _06403_;
	wire _06404_;
	wire _06405_;
	wire _06406_;
	wire _06407_;
	wire _06408_;
	wire _06409_;
	wire _06410_;
	wire _06411_;
	wire _06412_;
	wire _06413_;
	wire _06414_;
	wire _06415_;
	wire _06416_;
	wire _06417_;
	wire _06418_;
	wire _06419_;
	wire _06420_;
	wire _06421_;
	wire _06422_;
	wire _06423_;
	wire _06424_;
	wire _06425_;
	wire _06426_;
	wire _06427_;
	wire _06428_;
	wire _06429_;
	wire _06430_;
	wire _06431_;
	wire _06432_;
	wire _06433_;
	wire _06434_;
	wire _06435_;
	wire _06436_;
	wire _06437_;
	wire _06438_;
	wire _06439_;
	wire _06440_;
	wire _06441_;
	wire _06442_;
	wire _06443_;
	wire _06444_;
	wire _06445_;
	wire _06446_;
	wire _06447_;
	wire _06448_;
	wire _06449_;
	wire _06450_;
	wire _06451_;
	wire _06452_;
	wire _06453_;
	wire _06454_;
	wire _06455_;
	wire _06456_;
	wire _06457_;
	wire _06458_;
	wire _06459_;
	wire _06460_;
	wire _06461_;
	wire _06462_;
	wire _06463_;
	wire _06464_;
	wire _06465_;
	wire _06466_;
	input wire [13:0] io_in;
	output wire [13:0] io_out;
	wire \mchip.clock ;
	wire [11:0] \mchip.io_in ;
	wire [11:0] \mchip.io_out ;
	wire \mchip.reset ;
	wire \mchip.wrapper.clock ;
	reg \mchip.wrapper.currState ;
	wire [15:0] \mchip.wrapper.de.KEY ;
	wire [7:0] \mchip.wrapper.de.P1 ;
	wire [15:0] \mchip.wrapper.de.intxt ;
	wire [7:0] \mchip.wrapper.de.p1start ;
	wire [7:0] \mchip.wrapper.de.p2start ;
	wire [7:0] \mchip.wrapper.de.p3start ;
	wire [7:0] \mchip.wrapper.de.p4start ;
	wire [7:0] \mchip.wrapper.de.p5start ;
	wire [7:0] \mchip.wrapper.de.p6start ;
	wire [7:0] \mchip.wrapper.de.p7start ;
	wire [7:0] \mchip.wrapper.de.p8start ;
	wire [7:0] \mchip.wrapper.de.s11 ;
	wire [7:0] \mchip.wrapper.de.sub1.s1 ;
	wire [7:0] \mchip.wrapper.de.sub17.s1 ;
	wire [7:0] \mchip.wrapper.de.sub25.s1 ;
	wire [7:0] \mchip.wrapper.de.sub29.s1 ;
	wire [7:0] \mchip.wrapper.de.sub37.s1 ;
	wire [7:0] \mchip.wrapper.de.sub45.s1 ;
	wire [7:0] \mchip.wrapper.de.sub5.s1 ;
	wire [7:0] \mchip.wrapper.de.sub9.s1 ;
	wire [15:0] \mchip.wrapper.de.temp8 ;
	wire [3:0] \mchip.wrapper.display_sel ;
	wire [15:0] \mchip.wrapper.en.KEY ;
	wire [7:0] \mchip.wrapper.en.P1 ;
	wire [15:0] \mchip.wrapper.en.intxt ;
	wire [7:0] \mchip.wrapper.en.p1start ;
	wire [7:0] \mchip.wrapper.en.p2start ;
	wire [7:0] \mchip.wrapper.en.p3start ;
	wire [7:0] \mchip.wrapper.en.p4start ;
	wire [7:0] \mchip.wrapper.en.p5start ;
	wire [7:0] \mchip.wrapper.en.p6start ;
	wire [7:0] \mchip.wrapper.en.p7start ;
	wire [7:0] \mchip.wrapper.en.p8start ;
	wire [7:0] \mchip.wrapper.en.s11 ;
	wire [7:0] \mchip.wrapper.en.sub1.s1 ;
	wire [1:0] \mchip.wrapper.en.sub1.sel ;
	wire [7:0] \mchip.wrapper.en.sub17.s1 ;
	wire [1:0] \mchip.wrapper.en.sub2.sel ;
	wire [7:0] \mchip.wrapper.en.sub25.s1 ;
	wire [7:0] \mchip.wrapper.en.sub29.s1 ;
	wire [1:0] \mchip.wrapper.en.sub3.sel ;
	wire [7:0] \mchip.wrapper.en.sub37.s1 ;
	wire [1:0] \mchip.wrapper.en.sub4.sel ;
	wire [7:0] \mchip.wrapper.en.sub45.s1 ;
	wire [7:0] \mchip.wrapper.en.sub5.s1 ;
	wire [7:0] \mchip.wrapper.en.sub9.s1 ;
	wire [7:0] \mchip.wrapper.hex_out ;
	wire [3:0] \mchip.wrapper.i1.hexdigit ;
	wire [7:0] \mchip.wrapper.i1.seg ;
	wire [7:0] \mchip.wrapper.i10.seg ;
	wire [7:0] \mchip.wrapper.i11.seg ;
	wire [7:0] \mchip.wrapper.i12.seg ;
	wire [7:0] \mchip.wrapper.i13.seg ;
	wire [7:0] \mchip.wrapper.i14.seg ;
	wire [7:0] \mchip.wrapper.i15.seg ;
	wire [7:0] \mchip.wrapper.i16.seg ;
	wire [3:0] \mchip.wrapper.i2.hexdigit ;
	wire [7:0] \mchip.wrapper.i2.seg ;
	wire [3:0] \mchip.wrapper.i3.hexdigit ;
	wire [7:0] \mchip.wrapper.i3.seg ;
	wire [3:0] \mchip.wrapper.i4.hexdigit ;
	wire [7:0] \mchip.wrapper.i4.seg ;
	wire [3:0] \mchip.wrapper.i5.hexdigit ;
	wire [7:0] \mchip.wrapper.i5.seg ;
	wire [3:0] \mchip.wrapper.i6.hexdigit ;
	wire [7:0] \mchip.wrapper.i6.seg ;
	wire [3:0] \mchip.wrapper.i7.hexdigit ;
	wire [7:0] \mchip.wrapper.i7.seg ;
	wire [3:0] \mchip.wrapper.i8.hexdigit ;
	wire [7:0] \mchip.wrapper.i8.seg ;
	wire [7:0] \mchip.wrapper.i9.seg ;
	wire \mchip.wrapper.in_bit ;
	wire [15:0] \mchip.wrapper.intxt ;
	reg [15:0] \mchip.wrapper.intxtReg.Q ;
	wire \mchip.wrapper.intxtReg.clock ;
	wire \mchip.wrapper.intxtReg.en ;
	wire \mchip.wrapper.intxtReg.left ;
	wire \mchip.wrapper.intxtReg.serial ;
	wire [7:0] \mchip.wrapper.intxt_hex1 ;
	wire [7:0] \mchip.wrapper.intxt_hex2 ;
	wire [7:0] \mchip.wrapper.intxt_hex3 ;
	wire [7:0] \mchip.wrapper.intxt_hex4 ;
	wire [15:0] \mchip.wrapper.key ;
	reg [15:0] \mchip.wrapper.keyReg.Q ;
	wire \mchip.wrapper.keyReg.clock ;
	wire \mchip.wrapper.keyReg.en ;
	wire \mchip.wrapper.keyReg.left ;
	wire \mchip.wrapper.keyReg.serial ;
	wire [7:0] \mchip.wrapper.key_hex1 ;
	wire [7:0] \mchip.wrapper.key_hex2 ;
	wire [7:0] \mchip.wrapper.key_hex3 ;
	wire [7:0] \mchip.wrapper.key_hex4 ;
	wire [1:0] \mchip.wrapper.mode_sel ;
	wire \mchip.wrapper.nextState ;
	wire [7:0] \mchip.wrapper.outtxt_de_hex1 ;
	wire [7:0] \mchip.wrapper.outtxt_de_hex2 ;
	wire [7:0] \mchip.wrapper.outtxt_de_hex3 ;
	wire [7:0] \mchip.wrapper.outtxt_de_hex4 ;
	wire [7:0] \mchip.wrapper.outtxt_hex1 ;
	wire [7:0] \mchip.wrapper.outtxt_hex2 ;
	wire [7:0] \mchip.wrapper.outtxt_hex3 ;
	wire [7:0] \mchip.wrapper.outtxt_hex4 ;
	wire \mchip.wrapper.ready ;
	wire \mchip.wrapper.reset ;
	assign _04591_ = io_in[2] & ~io_in[3];
	assign _04701_ = ~(io_in[4] | io_in[5]);
	assign _04811_ = _04701_ & _04591_;
	assign _04922_ = \mchip.wrapper.intxtReg.Q [5] & \mchip.wrapper.intxtReg.Q [4];
	assign _05033_ = ~(\mchip.wrapper.intxtReg.Q [7] & \mchip.wrapper.intxtReg.Q [6]);
	assign _05141_ = _04922_ & ~_05033_;
	assign _05250_ = \mchip.wrapper.intxtReg.Q [4] | ~\mchip.wrapper.intxtReg.Q [5];
	assign _05360_ = ~(_05250_ | _05033_);
	assign _05471_ = \mchip.wrapper.intxtReg.Q [5] | ~\mchip.wrapper.intxtReg.Q [4];
	assign _05581_ = ~(_05471_ | _05033_);
	assign _05691_ = ~_05581_;
	assign _05802_ = \mchip.wrapper.intxtReg.Q [7] | ~\mchip.wrapper.intxtReg.Q [6];
	assign _05912_ = ~(_05802_ | _05250_);
	assign _06022_ = ~_05912_;
	assign _06101_ = ~(_05802_ | _05471_);
	assign _06112_ = \mchip.wrapper.intxtReg.Q [7] | \mchip.wrapper.intxtReg.Q [6];
	assign _06121_ = _06112_ | _05471_;
	assign _06132_ = \mchip.wrapper.intxtReg.Q [5] | \mchip.wrapper.intxtReg.Q [4];
	assign _06143_ = _06132_ | _06112_;
	assign _06153_ = _06143_ | ~_06121_;
	assign _06164_ = ~(_06112_ | _05250_);
	assign _06175_ = _06153_ & ~_06164_;
	assign _06185_ = _04922_ & ~_06112_;
	assign _06196_ = _06185_ | ~_06175_;
	assign _06207_ = ~(_06132_ | _05802_);
	assign _06217_ = _06196_ & ~_06207_;
	assign _06228_ = _06217_ | _06101_;
	assign _06239_ = _06022_ & ~_06228_;
	assign _06250_ = _04922_ & ~_05802_;
	assign _06261_ = _06239_ & ~_06250_;
	assign _06271_ = \mchip.wrapper.intxtReg.Q [6] | ~\mchip.wrapper.intxtReg.Q [7];
	assign _06281_ = ~(_06271_ | _06132_);
	assign _06291_ = _06261_ & ~_06281_;
	assign _06302_ = ~(_06271_ | _05471_);
	assign _06313_ = _06291_ & ~_06302_;
	assign _06324_ = ~(_06271_ | _05250_);
	assign _06335_ = _06313_ & ~_06324_;
	assign _06346_ = _04922_ & ~_06271_;
	assign _06357_ = _06346_ | _06335_;
	assign _06368_ = ~(_06132_ | _05033_);
	assign _06379_ = ~_06368_;
	assign _06390_ = _06379_ & _06357_;
	assign _06401_ = _05691_ & ~_06390_;
	assign _06412_ = _06401_ | _05360_;
	assign _06423_ = _06412_ | _05141_;
	assign _06433_ = _04811_ & ~_06423_;
	assign _06444_ = io_in[3] & ~io_in[2];
	assign _06455_ = _06444_ & _04701_;
	assign _06466_ = \mchip.wrapper.intxtReg.Q [8] & \mchip.wrapper.intxtReg.Q [9];
	assign _00010_ = ~(\mchip.wrapper.intxtReg.Q [10] & \mchip.wrapper.intxtReg.Q [11]);
	assign _00021_ = _06466_ & ~_00010_;
	assign _00032_ = \mchip.wrapper.intxtReg.Q [9] & ~\mchip.wrapper.intxtReg.Q [8];
	assign _00043_ = _00032_ & ~_00010_;
	assign _00054_ = \mchip.wrapper.intxtReg.Q [8] & ~\mchip.wrapper.intxtReg.Q [9];
	assign _00065_ = _00054_ & ~_00010_;
	assign _00076_ = ~_00065_;
	assign _00087_ = \mchip.wrapper.intxtReg.Q [10] & ~\mchip.wrapper.intxtReg.Q [11];
	assign _00098_ = _00087_ & _00032_;
	assign _00109_ = ~_00098_;
	assign _00120_ = _00087_ & _00054_;
	assign _00131_ = ~(\mchip.wrapper.intxtReg.Q [10] | \mchip.wrapper.intxtReg.Q [11]);
	assign _00142_ = _00131_ & _00054_;
	assign _00153_ = ~(\mchip.wrapper.intxtReg.Q [8] | \mchip.wrapper.intxtReg.Q [9]);
	assign _00164_ = _00153_ & _00131_;
	assign _00175_ = _00164_ & ~_00142_;
	assign _00186_ = _00131_ & _00032_;
	assign _00197_ = ~_00186_;
	assign _00208_ = _00197_ & ~_00175_;
	assign _00219_ = _00131_ & _06466_;
	assign _00230_ = ~_00219_;
	assign _00241_ = ~(_00230_ & _00208_);
	assign _00252_ = _00153_ & _00087_;
	assign _00263_ = _00241_ & ~_00252_;
	assign _00274_ = _00263_ | _00120_;
	assign _00285_ = _00109_ & ~_00274_;
	assign _00296_ = _00087_ & _06466_;
	assign _00307_ = _00285_ & ~_00296_;
	assign _00318_ = \mchip.wrapper.intxtReg.Q [11] & ~\mchip.wrapper.intxtReg.Q [10];
	assign _00329_ = _00318_ & _00153_;
	assign _00339_ = _00307_ & ~_00329_;
	assign _00350_ = _00318_ & _00054_;
	assign _00361_ = _00339_ & ~_00350_;
	assign _00372_ = _00318_ & _00032_;
	assign _00383_ = _00361_ & ~_00372_;
	assign _00394_ = _00318_ & _06466_;
	assign _00405_ = _00394_ | _00383_;
	assign _00415_ = _00153_ & ~_00010_;
	assign _00426_ = ~_00415_;
	assign _00437_ = _00426_ & _00405_;
	assign _00448_ = _00076_ & ~_00437_;
	assign _00459_ = _00448_ | _00043_;
	assign _00470_ = _00459_ | _00021_;
	assign _00481_ = _06455_ & ~_00470_;
	assign _00492_ = io_in[2] & io_in[3];
	assign _00503_ = _00492_ & _04701_;
	assign _00514_ = \mchip.wrapper.intxtReg.Q [14] & \mchip.wrapper.intxtReg.Q [15];
	assign _00525_ = ~(\mchip.wrapper.intxtReg.Q [12] & \mchip.wrapper.intxtReg.Q [13]);
	assign _00536_ = _00514_ & ~_00525_;
	assign _00547_ = \mchip.wrapper.intxtReg.Q [13] & ~\mchip.wrapper.intxtReg.Q [12];
	assign _00558_ = _00547_ & _00514_;
	assign _00569_ = \mchip.wrapper.intxtReg.Q [12] & ~\mchip.wrapper.intxtReg.Q [13];
	assign _00580_ = _00569_ & _00514_;
	assign _00591_ = ~_00580_;
	assign _00602_ = \mchip.wrapper.intxtReg.Q [15] | ~\mchip.wrapper.intxtReg.Q [14];
	assign _00613_ = _00547_ & ~_00602_;
	assign _00624_ = ~_00613_;
	assign _00635_ = _00569_ & ~_00602_;
	assign _00646_ = ~(\mchip.wrapper.intxtReg.Q [14] | \mchip.wrapper.intxtReg.Q [15]);
	assign _00657_ = _00646_ & _00569_;
	assign _00668_ = ~(\mchip.wrapper.intxtReg.Q [12] | \mchip.wrapper.intxtReg.Q [13]);
	assign _00679_ = _00668_ & _00646_;
	assign _00690_ = _00679_ & ~_00657_;
	assign _00701_ = _00646_ & _00547_;
	assign _00712_ = ~_00701_;
	assign _00723_ = _00712_ & ~_00690_;
	assign _00734_ = _00646_ & ~_00525_;
	assign _00745_ = ~_00734_;
	assign _00756_ = ~(_00745_ & _00723_);
	assign _00767_ = _00668_ & ~_00602_;
	assign _00778_ = _00756_ & ~_00767_;
	assign _00789_ = _00778_ | _00635_;
	assign _00800_ = _00624_ & ~_00789_;
	assign _00811_ = ~(_00602_ | _00525_);
	assign _00822_ = _00800_ & ~_00811_;
	assign _00833_ = \mchip.wrapper.intxtReg.Q [15] & ~\mchip.wrapper.intxtReg.Q [14];
	assign _00844_ = _00833_ & _00668_;
	assign _00855_ = _00822_ & ~_00844_;
	assign _00866_ = _00833_ & _00569_;
	assign _00877_ = _00855_ & ~_00866_;
	assign _00888_ = _00833_ & _00547_;
	assign _00899_ = _00877_ & ~_00888_;
	assign _00910_ = _00833_ & ~_00525_;
	assign _00921_ = _00910_ | _00899_;
	assign _00932_ = _00668_ & _00514_;
	assign _00943_ = ~_00932_;
	assign _00954_ = _00943_ & _00921_;
	assign _00965_ = _00591_ & ~_00954_;
	assign _00976_ = _00965_ | _00558_;
	assign _00987_ = _00976_ | _00536_;
	assign _00998_ = _00503_ & ~_00987_;
	assign _01009_ = _00998_ | _00481_;
	assign _01020_ = _01009_ | _06433_;
	assign _01031_ = ~(io_in[2] | io_in[3]);
	assign _01042_ = io_in[5] | ~io_in[4];
	assign _01053_ = _01031_ & ~_01042_;
	assign _01064_ = \mchip.wrapper.keyReg.Q [1] & \mchip.wrapper.keyReg.Q [0];
	assign _01075_ = ~(\mchip.wrapper.keyReg.Q [3] & \mchip.wrapper.keyReg.Q [2]);
	assign _01086_ = _01064_ & ~_01075_;
	assign _01097_ = \mchip.wrapper.keyReg.Q [0] | ~\mchip.wrapper.keyReg.Q [1];
	assign _01108_ = ~(_01097_ | _01075_);
	assign _01119_ = \mchip.wrapper.keyReg.Q [1] | ~\mchip.wrapper.keyReg.Q [0];
	assign _01130_ = ~(_01119_ | _01075_);
	assign _01141_ = ~_01130_;
	assign _01152_ = \mchip.wrapper.keyReg.Q [3] | ~\mchip.wrapper.keyReg.Q [2];
	assign _01163_ = ~(_01152_ | _01097_);
	assign _01174_ = ~_01163_;
	assign _01185_ = ~(_01152_ | _01119_);
	assign _01196_ = \mchip.wrapper.keyReg.Q [3] | \mchip.wrapper.keyReg.Q [2];
	assign _01207_ = _01196_ | _01119_;
	assign _01218_ = \mchip.wrapper.keyReg.Q [1] | \mchip.wrapper.keyReg.Q [0];
	assign _01229_ = _01218_ | _01196_;
	assign _01240_ = _01229_ | ~_01207_;
	assign _01251_ = ~(_01196_ | _01097_);
	assign _01262_ = _01240_ & ~_01251_;
	assign _01273_ = _01064_ & ~_01196_;
	assign _01284_ = _01273_ | ~_01262_;
	assign _01295_ = ~(_01218_ | _01152_);
	assign _01306_ = _01284_ & ~_01295_;
	assign _01317_ = _01306_ | _01185_;
	assign _01328_ = _01174_ & ~_01317_;
	assign _01339_ = _01064_ & ~_01152_;
	assign _01350_ = _01328_ & ~_01339_;
	assign _01361_ = \mchip.wrapper.keyReg.Q [2] | ~\mchip.wrapper.keyReg.Q [3];
	assign _01372_ = ~(_01361_ | _01218_);
	assign _01383_ = _01350_ & ~_01372_;
	assign _01394_ = ~(_01361_ | _01119_);
	assign _01405_ = _01383_ & ~_01394_;
	assign _01416_ = ~(_01361_ | _01097_);
	assign _01427_ = _01405_ & ~_01416_;
	assign _01438_ = _01064_ & ~_01361_;
	assign _01449_ = _01438_ | _01427_;
	assign _01460_ = ~(_01218_ | _01075_);
	assign _01471_ = ~_01460_;
	assign _01482_ = _01471_ & _01449_;
	assign _01493_ = _01141_ & ~_01482_;
	assign _01504_ = _01493_ | _01108_;
	assign _01515_ = _01504_ | _01086_;
	assign _01526_ = _01053_ & ~_01515_;
	assign _01537_ = _04591_ & ~_01042_;
	assign _01548_ = \mchip.wrapper.keyReg.Q [5] & \mchip.wrapper.keyReg.Q [4];
	assign _01559_ = ~(\mchip.wrapper.keyReg.Q [7] & \mchip.wrapper.keyReg.Q [6]);
	assign _01570_ = _01548_ & ~_01559_;
	assign _01581_ = \mchip.wrapper.keyReg.Q [4] | ~\mchip.wrapper.keyReg.Q [5];
	assign _01592_ = ~(_01581_ | _01559_);
	assign _01603_ = \mchip.wrapper.keyReg.Q [5] | ~\mchip.wrapper.keyReg.Q [4];
	assign _01614_ = ~(_01603_ | _01559_);
	assign _01625_ = ~_01614_;
	assign _01636_ = \mchip.wrapper.keyReg.Q [7] | ~\mchip.wrapper.keyReg.Q [6];
	assign _01647_ = ~(_01636_ | _01581_);
	assign _01657_ = ~_01647_;
	assign _01668_ = ~(_01636_ | _01603_);
	assign _01679_ = \mchip.wrapper.keyReg.Q [7] | \mchip.wrapper.keyReg.Q [6];
	assign _01690_ = ~(_01679_ | _01603_);
	assign _01701_ = \mchip.wrapper.keyReg.Q [5] | \mchip.wrapper.keyReg.Q [4];
	assign _01712_ = ~(_01701_ | _01679_);
	assign _01723_ = _01690_ | ~_01712_;
	assign _01734_ = ~(_01679_ | _01581_);
	assign _01745_ = _01723_ & ~_01734_;
	assign _01756_ = _01548_ & ~_01679_;
	assign _01767_ = _01756_ | ~_01745_;
	assign _01778_ = ~(_01701_ | _01636_);
	assign _01789_ = _01767_ & ~_01778_;
	assign _01800_ = _01789_ | _01668_;
	assign _01811_ = _01657_ & ~_01800_;
	assign _01822_ = _01548_ & ~_01636_;
	assign _01833_ = _01811_ & ~_01822_;
	assign _01844_ = \mchip.wrapper.keyReg.Q [6] | ~\mchip.wrapper.keyReg.Q [7];
	assign _01855_ = ~(_01844_ | _01701_);
	assign _01866_ = _01833_ & ~_01855_;
	assign _01877_ = ~(_01844_ | _01603_);
	assign _01888_ = _01866_ & ~_01877_;
	assign _01899_ = ~(_01844_ | _01581_);
	assign _01910_ = _01888_ & ~_01899_;
	assign _01921_ = _01548_ & ~_01844_;
	assign _01932_ = _01921_ | _01910_;
	assign _01943_ = ~(_01701_ | _01559_);
	assign _01954_ = ~_01943_;
	assign _01965_ = _01954_ & _01932_;
	assign _01976_ = _01625_ & ~_01965_;
	assign _01987_ = _01976_ | _01592_;
	assign _01997_ = _01987_ | _01570_;
	assign _02007_ = _01537_ & ~_01997_;
	assign _02018_ = _02007_ | _01526_;
	assign _02028_ = _06444_ & ~_01042_;
	assign _02039_ = \mchip.wrapper.keyReg.Q [9] & \mchip.wrapper.keyReg.Q [8];
	assign _02050_ = ~(\mchip.wrapper.keyReg.Q [11] & \mchip.wrapper.keyReg.Q [10]);
	assign _02059_ = _02039_ & ~_02050_;
	assign _02069_ = \mchip.wrapper.keyReg.Q [8] | ~\mchip.wrapper.keyReg.Q [9];
	assign _02079_ = ~(_02069_ | _02050_);
	assign _02089_ = \mchip.wrapper.keyReg.Q [9] | ~\mchip.wrapper.keyReg.Q [8];
	assign _02099_ = ~(_02089_ | _02050_);
	assign _02110_ = ~_02099_;
	assign _02121_ = \mchip.wrapper.keyReg.Q [11] | ~\mchip.wrapper.keyReg.Q [10];
	assign _02130_ = ~(_02121_ | _02069_);
	assign _02141_ = ~_02130_;
	assign _02152_ = ~(_02121_ | _02089_);
	assign _02163_ = \mchip.wrapper.keyReg.Q [11] | \mchip.wrapper.keyReg.Q [10];
	assign _02174_ = _02163_ | _02089_;
	assign _02185_ = \mchip.wrapper.keyReg.Q [9] | \mchip.wrapper.keyReg.Q [8];
	assign _02196_ = _02185_ | _02163_;
	assign _02205_ = _02196_ | ~_02174_;
	assign _02216_ = ~(_02163_ | _02069_);
	assign _02227_ = _02205_ & ~_02216_;
	assign _02238_ = _02039_ & ~_02163_;
	assign _02249_ = _02238_ | ~_02227_;
	assign _02260_ = ~(_02185_ | _02121_);
	assign _02271_ = _02249_ & ~_02260_;
	assign _02282_ = _02271_ | _02152_;
	assign _02293_ = _02141_ & ~_02282_;
	assign _02304_ = _02039_ & ~_02121_;
	assign _02315_ = _02293_ & ~_02304_;
	assign _02326_ = \mchip.wrapper.keyReg.Q [10] | ~\mchip.wrapper.keyReg.Q [11];
	assign _02337_ = ~(_02326_ | _02185_);
	assign _02348_ = _02315_ & ~_02337_;
	assign _02359_ = ~(_02326_ | _02089_);
	assign _02370_ = _02348_ & ~_02359_;
	assign _02381_ = ~(_02326_ | _02069_);
	assign _02392_ = _02370_ & ~_02381_;
	assign _02403_ = _02039_ & ~_02326_;
	assign _02414_ = _02403_ | _02392_;
	assign _02425_ = ~(_02185_ | _02050_);
	assign _02436_ = ~_02425_;
	assign _02447_ = _02436_ & _02414_;
	assign _02458_ = _02110_ & ~_02447_;
	assign _02469_ = _02458_ | _02079_;
	assign _02480_ = _02469_ | _02059_;
	assign _02491_ = _02028_ & ~_02480_;
	assign _02502_ = _00492_ & ~_01042_;
	assign _02513_ = \mchip.wrapper.keyReg.Q [13] & \mchip.wrapper.keyReg.Q [12];
	assign _02524_ = ~(\mchip.wrapper.keyReg.Q [15] & \mchip.wrapper.keyReg.Q [14]);
	assign _02535_ = _02513_ & ~_02524_;
	assign _02546_ = \mchip.wrapper.keyReg.Q [12] | ~\mchip.wrapper.keyReg.Q [13];
	assign _02557_ = ~(_02546_ | _02524_);
	assign _02568_ = \mchip.wrapper.keyReg.Q [13] | ~\mchip.wrapper.keyReg.Q [12];
	assign _02579_ = ~(_02568_ | _02524_);
	assign _02590_ = ~_02579_;
	assign _02601_ = \mchip.wrapper.keyReg.Q [15] | ~\mchip.wrapper.keyReg.Q [14];
	assign _02612_ = ~(_02601_ | _02546_);
	assign _02623_ = ~_02612_;
	assign _02634_ = ~(_02601_ | _02568_);
	assign _02645_ = \mchip.wrapper.keyReg.Q [15] | \mchip.wrapper.keyReg.Q [14];
	assign _02656_ = ~(_02645_ | _02568_);
	assign _02667_ = \mchip.wrapper.keyReg.Q [13] | \mchip.wrapper.keyReg.Q [12];
	assign _02678_ = ~(_02667_ | _02645_);
	assign _02689_ = _02656_ | ~_02678_;
	assign _02700_ = ~(_02645_ | _02546_);
	assign _02711_ = _02689_ & ~_02700_;
	assign _02722_ = _02513_ & ~_02645_;
	assign _02733_ = _02722_ | ~_02711_;
	assign _02744_ = ~(_02667_ | _02601_);
	assign _02755_ = _02733_ & ~_02744_;
	assign _02766_ = _02755_ | _02634_;
	assign _02777_ = _02623_ & ~_02766_;
	assign _02788_ = _02513_ & ~_02601_;
	assign _02799_ = _02777_ & ~_02788_;
	assign _02810_ = \mchip.wrapper.keyReg.Q [14] | ~\mchip.wrapper.keyReg.Q [15];
	assign _02821_ = ~(_02810_ | _02667_);
	assign _02832_ = _02799_ & ~_02821_;
	assign _02843_ = ~(_02810_ | _02568_);
	assign _02854_ = _02832_ & ~_02843_;
	assign _02865_ = ~(_02810_ | _02546_);
	assign _02876_ = _02854_ & ~_02865_;
	assign _02887_ = _02513_ & ~_02810_;
	assign _02898_ = _02887_ | _02876_;
	assign _02909_ = ~(_02667_ | _02524_);
	assign _02920_ = ~_02909_;
	assign _02931_ = _02920_ & _02898_;
	assign _02942_ = _02590_ & ~_02931_;
	assign _02953_ = _02942_ | _02557_;
	assign _02964_ = _02953_ | _02535_;
	assign _02975_ = _02502_ & ~_02964_;
	assign _02986_ = _02975_ | _02491_;
	assign _02997_ = _02986_ | _02018_;
	assign _03008_ = _02997_ | _01020_;
	assign _03019_ = io_in[4] | ~io_in[5];
	assign _03030_ = _01031_ & ~_03019_;
	assign _03041_ = ~\mchip.wrapper.keyReg.Q [1];
	assign _03052_ = ~(\mchip.wrapper.keyReg.Q [9] ^ \mchip.wrapper.keyReg.Q [1]);
	assign _03063_ = _03052_ ^ \mchip.wrapper.keyReg.Q [1];
	assign _03074_ = _03063_ ^ \mchip.wrapper.keyReg.Q [9];
	assign _03085_ = \mchip.wrapper.keyReg.Q [14] ^ \mchip.wrapper.keyReg.Q [6];
	assign _03096_ = ~_03085_;
	assign _03107_ = ~\mchip.wrapper.keyReg.Q [6];
	assign _03118_ = ~\mchip.wrapper.keyReg.Q [14];
	assign _03129_ = _03085_ ^ \mchip.wrapper.keyReg.Q [6];
	assign _03140_ = _03129_ ^ _03118_;
	assign _03151_ = ~\mchip.wrapper.keyReg.Q [15];
	assign _03162_ = \mchip.wrapper.keyReg.Q [7] ^ \mchip.wrapper.keyReg.Q [15];
	assign _03173_ = _03162_ ^ \mchip.wrapper.keyReg.Q [7];
	assign _03184_ = _03173_ ^ _03151_;
	assign _03195_ = ~\mchip.wrapper.keyReg.Q [7];
	assign _03206_ = _03162_ ^ _03195_;
	assign _03217_ = _03206_ ^ \mchip.wrapper.keyReg.Q [15];
	assign _03228_ = ~(\mchip.wrapper.keyReg.Q [7] ^ \mchip.wrapper.keyReg.Q [15]);
	assign _03239_ = _03228_ ^ \mchip.wrapper.keyReg.Q [7];
	assign _03250_ = _03239_ ^ _03151_;
	assign _03261_ = ~_03217_;
	assign _03272_ = _03250_ ^ \mchip.wrapper.intxtReg.Q [7];
	assign _03283_ = ~(\mchip.wrapper.keyReg.Q [14] ^ \mchip.wrapper.keyReg.Q [6]);
	assign _03294_ = _03283_ ^ \mchip.wrapper.keyReg.Q [6];
	assign _03305_ = _03294_ ^ _03118_;
	assign _03316_ = _03305_ ^ \mchip.wrapper.intxtReg.Q [6];
	assign _03327_ = ~(_03316_ & _03272_);
	assign _03338_ = _03327_ | _03217_;
	assign _03349_ = _03272_ & ~_03316_;
	assign _03360_ = _03349_ & _03206_;
	assign _03371_ = _03338_ & ~_03360_;
	assign _03382_ = ~_03162_;
	assign _03393_ = _03316_ & ~_03272_;
	assign _03404_ = _03393_ & ~_03382_;
	assign _03415_ = _03371_ & ~_03404_;
	assign _03426_ = ~(_03316_ | _03272_);
	assign _03437_ = (_03426_ ? _03195_ : _03415_);
	assign _03448_ = ~\mchip.wrapper.keyReg.Q [13];
	assign _03459_ = \mchip.wrapper.keyReg.Q [13] ^ \mchip.wrapper.keyReg.Q [5];
	assign _03470_ = _03459_ ^ \mchip.wrapper.keyReg.Q [5];
	assign _03481_ = _03470_ ^ _03448_;
	assign _03492_ = ~(_03481_ ^ \mchip.wrapper.intxtReg.Q [5]);
	assign _03503_ = ~(\mchip.wrapper.keyReg.Q [4] ^ \mchip.wrapper.keyReg.Q [12]);
	assign _03514_ = _03503_ ^ \mchip.wrapper.keyReg.Q [4];
	assign _03525_ = _03514_ ^ \mchip.wrapper.keyReg.Q [12];
	assign _03536_ = ~(_03525_ ^ \mchip.wrapper.intxtReg.Q [4]);
	assign _03547_ = ~(_03536_ & _03492_);
	assign _03568_ = _03184_ | _03547_;
	assign _03579_ = ~_03173_;
	assign _03590_ = _03492_ & ~_03536_;
	assign _03601_ = _03590_ & ~_03579_;
	assign _03612_ = _03568_ & ~_03601_;
	assign _03623_ = _03536_ & ~_03492_;
	assign _03634_ = _03623_ & ~_03382_;
	assign _03645_ = _03612_ & ~_03634_;
	assign _03656_ = _03536_ | _03492_;
	assign _03667_ = _03217_ ^ \mchip.wrapper.keyReg.Q [7];
	assign _03678_ = (_03656_ ? _03645_ : _03667_);
	assign _03689_ = ~(\mchip.wrapper.keyReg.Q [10] ^ \mchip.wrapper.keyReg.Q [2]);
	assign _03700_ = _03689_ ^ \mchip.wrapper.keyReg.Q [2];
	assign _03711_ = _03700_ ^ \mchip.wrapper.keyReg.Q [10];
	assign _03722_ = ~(_03711_ ^ \mchip.wrapper.intxtReg.Q [2]);
	assign _03733_ = ~\mchip.wrapper.keyReg.Q [3];
	assign _03744_ = ~(\mchip.wrapper.keyReg.Q [3] ^ \mchip.wrapper.keyReg.Q [11]);
	assign _03755_ = _03744_ ^ _03733_;
	assign _03766_ = _03755_ ^ \mchip.wrapper.keyReg.Q [11];
	assign _03777_ = ~(_03766_ ^ \mchip.wrapper.intxtReg.Q [3]);
	assign _03788_ = _03777_ | _03722_;
	assign _03799_ = _03239_ ^ \mchip.wrapper.keyReg.Q [15];
	assign _03810_ = ~_03799_;
	assign _03821_ = _03810_ | _03788_;
	assign _03832_ = ~_03239_;
	assign _03843_ = _03722_ & ~_03777_;
	assign _03854_ = _03843_ & ~_03832_;
	assign _03865_ = _03821_ & ~_03854_;
	assign _03876_ = ~_03228_;
	assign _03887_ = _03777_ & ~_03722_;
	assign _03898_ = _03887_ & ~_03876_;
	assign _03909_ = _03865_ & ~_03898_;
	assign _03920_ = ~(_03777_ & _03722_);
	assign _00996_ = _03184_ ^ _03195_;
	assign _03941_ = (_03920_ ? _03909_ : _00996_);
	assign _03952_ = ~(\mchip.wrapper.keyReg.Q [8] ^ \mchip.wrapper.keyReg.Q [0]);
	assign _03963_ = _03952_ ^ \mchip.wrapper.keyReg.Q [0];
	assign _00086_ = _03963_ ^ \mchip.wrapper.keyReg.Q [8];
	assign _03984_ = _00086_ ^ \mchip.wrapper.intxtReg.Q [0];
	assign _04015_ = _03074_ ^ \mchip.wrapper.intxtReg.Q [1];
	assign _04026_ = _04015_ | _03984_;
	assign _04067_ = _03810_ | _04026_;
	assign _04078_ = _03984_ & ~_04015_;
	assign _04089_ = _04078_ & ~_03239_;
	assign _04100_ = _04067_ & ~_04089_;
	assign _04111_ = ~\mchip.wrapper.keyReg.Q [8];
	assign _04122_ = _03963_ ^ _04111_;
	assign _04133_ = _04122_ ^ \mchip.wrapper.intxtReg.Q [0];
	assign _04144_ = ~\mchip.wrapper.keyReg.Q [9];
	assign _00051_ = _03063_ ^ _04144_;
	assign _04165_ = _00051_ ^ \mchip.wrapper.intxtReg.Q [1];
	assign _04176_ = _04133_ & ~_04165_;
	assign _04187_ = _04176_ & ~_03228_;
	assign _04198_ = _04100_ & ~_04187_;
	assign _04209_ = _03984_ & ~_04165_;
	assign _04230_ = _03799_ ^ \mchip.wrapper.keyReg.Q [7];
	assign _04241_ = ~_04230_;
	assign _04252_ = (_04209_ ? _04241_ : _04198_);
	assign _04263_ = ~(\mchip.wrapper.keyReg.Q [15] ^ \mchip.wrapper.intxtReg.Q [15]);
	assign _04274_ = _04263_ ^ _04252_;
	assign _04285_ = _04274_ ^ _03941_;
	assign _04296_ = _04285_ ^ _03678_;
	assign _04307_ = _04296_ ^ _03437_;
	assign _04318_ = _04307_ ^ _03228_;
	assign _04329_ = _03327_ | _03140_;
	assign _04340_ = _03349_ & _03129_;
	assign _04351_ = _04329_ & ~_04340_;
	assign _04362_ = _03393_ & ~_03096_;
	assign _04373_ = _04351_ & ~_04362_;
	assign _04384_ = (_03426_ ? _03107_ : _04373_);
	assign _04405_ = _03305_ | _03547_;
	assign _04416_ = _03590_ & ~_03294_;
	assign _04427_ = _04405_ & ~_04416_;
	assign _04438_ = ~_03283_;
	assign _04449_ = _03623_ & ~_04438_;
	assign _04460_ = _04427_ & ~_04449_;
	assign _04471_ = _03140_ ^ \mchip.wrapper.keyReg.Q [6];
	assign _04481_ = (_03656_ ? _04460_ : _04471_);
	assign _04492_ = _03305_ | _03788_;
	assign _04503_ = ~_03294_;
	assign _04514_ = _03843_ & ~_04503_;
	assign _04525_ = _04492_ & ~_04514_;
	assign _04536_ = _03887_ & ~_04438_;
	assign _04547_ = _04525_ & ~_04536_;
	assign _04558_ = _03305_ ^ \mchip.wrapper.keyReg.Q [6];
	assign _04569_ = (_03920_ ? _04547_ : _04558_);
	assign _01835_ = ~_03305_;
	assign _04590_ = _04026_ | _01835_;
	assign _04602_ = _04078_ & ~_04503_;
	assign _04613_ = _04590_ & ~_04602_;
	assign _04624_ = _04176_ & ~_04438_;
	assign _04635_ = _04613_ & ~_04624_;
	assign _04646_ = (_04209_ ? _04558_ : _04635_);
	assign _04657_ = _03294_ ^ \mchip.wrapper.intxtReg.Q [14];
	assign _04667_ = _04657_ ^ _04646_;
	assign _04678_ = _04667_ ^ _04569_;
	assign _04689_ = _04678_ ^ _04481_;
	assign _04700_ = _04689_ ^ _04384_;
	assign _04712_ = _04700_ ^ _03283_;
	assign _04723_ = ~(_04712_ & _04318_);
	assign _04734_ = _04723_ | ~_03261_;
	assign _04745_ = _04318_ & ~_04712_;
	assign _04756_ = _04745_ & _03206_;
	assign _04767_ = _04734_ & ~_04756_;
	assign _04778_ = _04712_ & ~_04318_;
	assign _04788_ = _04778_ & ~_03382_;
	assign _04799_ = _04767_ & ~_04788_;
	assign _04810_ = ~(_04712_ | _04318_);
	assign _04822_ = (_04810_ ? _03195_ : _04799_);
	assign _04833_ = ~\mchip.wrapper.keyReg.Q [5];
	assign _04844_ = _03481_ | _03327_;
	assign _04855_ = ~_03470_;
	assign _04866_ = _03349_ & ~_04855_;
	assign _04877_ = _04844_ & ~_04866_;
	assign _04888_ = ~_03459_;
	assign _04899_ = _03393_ & ~_04888_;
	assign _04910_ = _04877_ & ~_04899_;
	assign _04921_ = (_03426_ ? _04833_ : _04910_);
	assign _04933_ = ~(\mchip.wrapper.keyReg.Q [13] ^ \mchip.wrapper.keyReg.Q [5]);
	assign _04944_ = _04933_ ^ \mchip.wrapper.keyReg.Q [5];
	assign _04955_ = _04944_ ^ \mchip.wrapper.keyReg.Q [13];
	assign _04966_ = _04955_ | _03547_;
	assign _04977_ = _03590_ & ~_04944_;
	assign _04988_ = _04966_ & ~_04977_;
	assign _04999_ = ~_04933_;
	assign _05010_ = _03623_ & ~_04999_;
	assign _05021_ = _04988_ & ~_05010_;
	assign _05032_ = _03481_ ^ \mchip.wrapper.keyReg.Q [5];
	assign _05044_ = (_03656_ ? _05021_ : _05032_);
	assign _02450_ = ~_04955_;
	assign _05075_ = _02450_ | _03788_;
	assign _05086_ = _03843_ & ~_04944_;
	assign _05096_ = _05075_ & ~_05086_;
	assign _05107_ = _03887_ & ~_04999_;
	assign _05118_ = _05096_ & ~_05107_;
	assign _05129_ = _04955_ ^ _04833_;
	assign _05140_ = (_03920_ ? _05118_ : _05129_);
	assign _05152_ = _03470_ ^ \mchip.wrapper.keyReg.Q [13];
	assign _05163_ = _05152_ | _04026_;
	assign _05174_ = _04078_ & ~_03470_;
	assign _05185_ = _05163_ & ~_05174_;
	assign _05196_ = _04176_ & ~_04888_;
	assign _05207_ = _05185_ & ~_05196_;
	assign _01735_ = ~_05129_;
	assign _05238_ = (_04209_ ? _01735_ : _05207_);
	assign _05249_ = _03470_ ^ \mchip.wrapper.intxtReg.Q [13];
	assign _05261_ = _05249_ ^ _05238_;
	assign _05272_ = _05261_ ^ _05140_;
	assign _05283_ = _05272_ ^ _05044_;
	assign _05293_ = _05283_ ^ _04921_;
	assign _05304_ = _05293_ ^ _03459_;
	assign _05315_ = ~\mchip.wrapper.keyReg.Q [12];
	assign _05326_ = \mchip.wrapper.keyReg.Q [4] ^ \mchip.wrapper.keyReg.Q [12];
	assign _05337_ = _05326_ ^ \mchip.wrapper.keyReg.Q [4];
	assign _05348_ = _05337_ ^ _05315_;
	assign _05359_ = _05348_ | _03327_;
	assign _05371_ = ~_05337_;
	assign _05382_ = _03349_ & ~_05371_;
	assign _05393_ = _05359_ & ~_05382_;
	assign _05404_ = ~_05326_;
	assign _05415_ = _03393_ & ~_05404_;
	assign _05426_ = _05393_ & ~_05415_;
	assign _05437_ = (_03426_ ? \mchip.wrapper.keyReg.Q [4] : _05426_);
	assign _05448_ = _03547_ | _03525_;
	assign _05459_ = _03590_ & ~_03514_;
	assign _05470_ = _05448_ & ~_05459_;
	assign _05482_ = ~_03503_;
	assign _05493_ = _03623_ & ~_05482_;
	assign _05504_ = _05470_ & ~_05493_;
	assign _05515_ = _05348_ ^ \mchip.wrapper.keyReg.Q [4];
	assign _05526_ = (_03656_ ? _05504_ : _05515_);
	assign _05537_ = _05337_ ^ \mchip.wrapper.keyReg.Q [12];
	assign _05548_ = _05537_ | _03788_;
	assign _05558_ = _03843_ & ~_05337_;
	assign _05569_ = _05548_ & ~_05558_;
	assign _05580_ = _03887_ & ~_05404_;
	assign _05592_ = _05569_ & ~_05580_;
	assign _01110_ = _03525_ ^ \mchip.wrapper.keyReg.Q [4];
	assign _05613_ = (_03920_ ? _05592_ : _01110_);
	assign _05624_ = ~\mchip.wrapper.keyReg.Q [4];
	assign _05635_ = _03503_ ^ _05624_;
	assign _05646_ = _05635_ ^ _05315_;
	assign _05657_ = _05646_ | _04026_;
	assign _05668_ = _04078_ & ~_05635_;
	assign _05679_ = _05657_ & ~_05668_;
	assign _05690_ = _04176_ & ~_03503_;
	assign _05702_ = _05679_ & ~_05690_;
	assign _05713_ = _05537_ ^ \mchip.wrapper.keyReg.Q [4];
	assign _05724_ = (_04209_ ? _05713_ : _05702_);
	assign _05735_ = _03514_ ^ \mchip.wrapper.intxtReg.Q [12];
	assign _05746_ = _05735_ ^ _05724_;
	assign _05757_ = _05746_ ^ _05613_;
	assign _05768_ = _05757_ ^ _05526_;
	assign _05779_ = _05768_ ^ _05437_;
	assign _05790_ = _05779_ ^ _03503_;
	assign _05801_ = ~(_05790_ & _05304_);
	assign _05813_ = _05801_ | _03184_;
	assign _05824_ = _05304_ & ~_05790_;
	assign _05835_ = _05824_ & ~_03579_;
	assign _05845_ = _05813_ & ~_05835_;
	assign _05856_ = _05790_ & ~_05304_;
	assign _05867_ = _05856_ & ~_03382_;
	assign _05878_ = _05845_ & ~_05867_;
	assign _05889_ = ~(_05790_ | _05304_);
	assign _05900_ = (_05889_ ? _03667_ : _05878_);
	assign _05911_ = ~_03744_;
	assign _05923_ = ~\mchip.wrapper.keyReg.Q [11];
	assign _05934_ = _03755_ ^ _05923_;
	assign _05945_ = ~_05934_;
	assign _05956_ = _05945_ | _03327_;
	assign _00271_ = ~_03755_;
	assign _05977_ = _03349_ & ~_00271_;
	assign _05988_ = _05956_ & ~_05977_;
	assign _05999_ = _03393_ & ~_05911_;
	assign _06010_ = _05988_ & ~_05999_;
	assign _06021_ = (_03426_ ? _03733_ : _06010_);
	assign _06063_ = _05945_ | _03547_;
	assign _06074_ = _03590_ & ~_03755_;
	assign _06085_ = _06063_ & ~_06074_;
	assign _06094_ = _03623_ & ~_05911_;
	assign _06098_ = _06085_ & ~_06094_;
	assign _06099_ = _05934_ ^ _03733_;
	assign _06100_ = (_03656_ ? _06098_ : _06099_);
	assign _06102_ = _05945_ | _03788_;
	assign _06103_ = _03843_ & ~_03755_;
	assign _06104_ = _06102_ & ~_06103_;
	assign _06105_ = _03887_ & ~_03744_;
	assign _06106_ = _06104_ & ~_06105_;
	assign _06107_ = _05934_ ^ \mchip.wrapper.keyReg.Q [3];
	assign _06108_ = ~_06107_;
	assign _06109_ = (_03920_ ? _06106_ : _06108_);
	assign _06110_ = \mchip.wrapper.keyReg.Q [3] ^ \mchip.wrapper.keyReg.Q [11];
	assign _06111_ = _06110_ ^ _03733_;
	assign _06113_ = _06111_ ^ _05923_;
	assign _06114_ = _06113_ | _04026_;
	assign _06115_ = ~_06111_;
	assign _06116_ = _04078_ & ~_06115_;
	assign _06117_ = _06114_ & ~_06116_;
	assign _06118_ = _04176_ & ~_06110_;
	assign _06119_ = _06117_ & ~_06118_;
	assign _02616_ = ~_06099_;
	assign _06120_ = (_04209_ ? _02616_ : _06119_);
	assign _06122_ = \mchip.wrapper.keyReg.Q [11] ^ \mchip.wrapper.intxtReg.Q [11];
	assign _06123_ = _06122_ ^ _06120_;
	assign _06124_ = _06123_ ^ _06109_;
	assign _06125_ = _06124_ ^ _06100_;
	assign _06126_ = _06125_ ^ _06021_;
	assign _06127_ = _06126_ ^ _05911_;
	assign _06128_ = ~_03689_;
	assign _06129_ = ~\mchip.wrapper.keyReg.Q [2];
	assign _06130_ = \mchip.wrapper.keyReg.Q [10] ^ \mchip.wrapper.keyReg.Q [2];
	assign _06131_ = _06130_ ^ \mchip.wrapper.keyReg.Q [2];
	assign _06133_ = _06131_ ^ \mchip.wrapper.keyReg.Q [10];
	assign _06134_ = ~_06133_;
	assign _06135_ = _06134_ | _03327_;
	assign _06136_ = ~_06131_;
	assign _06137_ = _03349_ & ~_06136_;
	assign _06138_ = _06135_ & ~_06137_;
	assign _06139_ = ~_06130_;
	assign _06140_ = _03393_ & ~_06139_;
	assign _06141_ = _06138_ & ~_06140_;
	assign _06142_ = (_03426_ ? _06129_ : _06141_);
	assign _06144_ = ~\mchip.wrapper.keyReg.Q [10];
	assign _06145_ = _06131_ ^ _06144_;
	assign _06146_ = ~_06145_;
	assign _06147_ = _06146_ | _03547_;
	assign _06148_ = _03590_ & ~_06136_;
	assign _06149_ = _06147_ & ~_06148_;
	assign _06150_ = _03623_ & ~_06139_;
	assign _06151_ = _06149_ & ~_06150_;
	assign _01188_ = _06133_ ^ _06129_;
	assign _06152_ = (_03656_ ? _06151_ : _01188_);
	assign _06154_ = _06134_ | _03788_;
	assign _06155_ = _03843_ & ~_06136_;
	assign _06156_ = _06154_ & ~_06155_;
	assign _06157_ = _03887_ & ~_06139_;
	assign _06158_ = _06156_ & ~_06157_;
	assign _06159_ = _06145_ ^ _06129_;
	assign _06160_ = ~_06159_;
	assign _06161_ = (_03920_ ? _06158_ : _06160_);
	assign _06162_ = _06130_ ^ _06129_;
	assign _06163_ = _06162_ ^ _06144_;
	assign _06165_ = _06163_ | _04026_;
	assign _06166_ = ~_06162_;
	assign _06167_ = _04078_ & ~_06166_;
	assign _06168_ = _06165_ & ~_06167_;
	assign _06169_ = _04176_ & ~_06130_;
	assign _06170_ = _06168_ & ~_06169_;
	assign _06171_ = (_04209_ ? _01188_ : _06170_);
	assign _06172_ = _03700_ ^ \mchip.wrapper.intxtReg.Q [10];
	assign _06173_ = _06172_ ^ _06171_;
	assign _06174_ = _06173_ ^ _06161_;
	assign _06176_ = _06174_ ^ _06152_;
	assign _06177_ = _06176_ ^ _06142_;
	assign _06178_ = _06177_ ^ _06128_;
	assign _06179_ = _06178_ | _06127_;
	assign _06180_ = _06179_ | _03810_;
	assign _06181_ = _06177_ ^ _03689_;
	assign _06182_ = _06127_ | _06181_;
	assign _06183_ = _03239_ & ~_06182_;
	assign _06184_ = _06180_ & ~_06183_;
	assign _06186_ = ~(_06127_ & _06181_);
	assign _06187_ = _03228_ & ~_06186_;
	assign _06188_ = _06184_ & ~_06187_;
	assign _06189_ = _06127_ & ~_06181_;
	assign _06190_ = (_06189_ ? _00996_ : _06188_);
	assign _06191_ = ~_03052_;
	assign _06192_ = ~_03074_;
	assign _06193_ = _03327_ | _06192_;
	assign _06194_ = _03349_ & ~_03063_;
	assign _06195_ = _06193_ & ~_06194_;
	assign _06197_ = _03393_ & ~_06191_;
	assign _06198_ = _06195_ & ~_06197_;
	assign _06199_ = (_03426_ ? \mchip.wrapper.keyReg.Q [1] : _06198_);
	assign _06200_ = \mchip.wrapper.keyReg.Q [9] ^ \mchip.wrapper.keyReg.Q [1];
	assign _06201_ = _06200_ ^ \mchip.wrapper.keyReg.Q [1];
	assign _06202_ = _06201_ ^ \mchip.wrapper.keyReg.Q [9];
	assign _06203_ = _06202_ | _03547_;
	assign _06204_ = _03590_ & ~_06201_;
	assign _06205_ = _06203_ & ~_06204_;
	assign _06206_ = ~_06200_;
	assign _06208_ = _03623_ & ~_06206_;
	assign _06209_ = _06205_ & ~_06208_;
	assign _06210_ = _03074_ ^ _03041_;
	assign _06211_ = ~_06210_;
	assign _06212_ = (_03656_ ? _06209_ : _06211_);
	assign _06213_ = _03074_ | _03788_;
	assign _00344_ = ~_03063_;
	assign _06214_ = _03843_ & ~_00344_;
	assign _06215_ = _06213_ & ~_06214_;
	assign _06216_ = _03887_ & ~_06191_;
	assign _06218_ = _06215_ & ~_06216_;
	assign _06219_ = _06202_ ^ _03041_;
	assign _06220_ = ~_06219_;
	assign _06221_ = (_03920_ ? _06218_ : _06220_);
	assign _06222_ = _06200_ ^ _03041_;
	assign _06223_ = _06222_ ^ _04144_;
	assign _06224_ = _06223_ | _04026_;
	assign _06225_ = ~_06222_;
	assign _06226_ = _04078_ & ~_06225_;
	assign _06227_ = _06224_ & ~_06226_;
	assign _06229_ = _04176_ & ~_06200_;
	assign _06230_ = _06227_ & ~_06229_;
	assign _06231_ = _00051_ ^ _03041_;
	assign _06232_ = (_04209_ ? _06231_ : _06230_);
	assign _06233_ = _03063_ ^ \mchip.wrapper.intxtReg.Q [9];
	assign _06234_ = _06233_ ^ _06232_;
	assign _06235_ = _06234_ ^ _06221_;
	assign _06236_ = _06235_ ^ _06212_;
	assign _06237_ = _06236_ ^ _06199_;
	assign _06238_ = _06237_ ^ _06191_;
	assign _06240_ = ~_03952_;
	assign _06241_ = \mchip.wrapper.keyReg.Q [8] ^ \mchip.wrapper.keyReg.Q [0];
	assign _06242_ = _06241_ ^ \mchip.wrapper.keyReg.Q [0];
	assign _06243_ = _06242_ ^ _04111_;
	assign _06244_ = _06243_ | _03327_;
	assign _06245_ = ~_06242_;
	assign _06246_ = _03349_ & ~_06245_;
	assign _06247_ = _06244_ & ~_06246_;
	assign _06248_ = ~_06241_;
	assign _06249_ = _03393_ & ~_06248_;
	assign _06251_ = _06247_ & ~_06249_;
	assign _06252_ = (_03426_ ? \mchip.wrapper.keyReg.Q [0] : _06251_);
	assign _06253_ = _00086_ | _03547_;
	assign _06254_ = _03590_ & ~_03963_;
	assign _06255_ = _06253_ & ~_06254_;
	assign _06256_ = _03623_ & ~_06240_;
	assign _06257_ = _06255_ & ~_06256_;
	assign _06258_ = _06243_ ^ \mchip.wrapper.keyReg.Q [0];
	assign _06259_ = ~_06258_;
	assign _06260_ = (_03656_ ? _06257_ : _06259_);
	assign _06262_ = ~\mchip.wrapper.keyReg.Q [0];
	assign _06263_ = _06241_ ^ _06262_;
	assign _06264_ = _06263_ ^ \mchip.wrapper.keyReg.Q [8];
	assign _02279_ = ~_06264_;
	assign _06265_ = _02279_ | _03788_;
	assign _06266_ = ~_06263_;
	assign _06267_ = _03843_ & ~_06266_;
	assign _06268_ = _06265_ & ~_06267_;
	assign _06269_ = _03887_ & ~_06241_;
	assign _06270_ = _06268_ & ~_06269_;
	assign _06272_ = _04122_ ^ \mchip.wrapper.keyReg.Q [0];
	assign _06273_ = ~_06272_;
	assign _06274_ = (_03920_ ? _06270_ : _06273_);
	assign _06275_ = _06264_ | _04026_;
	assign _06276_ = _04078_ & ~_06263_;
	assign _06277_ = _06275_ & ~_06276_;
	assign _06278_ = _04176_ & ~_06241_;
	assign _06279_ = _06277_ & ~_06278_;
	assign _06280_ = _06264_ ^ \mchip.wrapper.keyReg.Q [0];
	assign _06282_ = (_04209_ ? _06280_ : _06279_);
	assign _06283_ = _03963_ ^ \mchip.wrapper.intxtReg.Q [8];
	assign _06284_ = _06283_ ^ _06282_;
	assign _06285_ = _06284_ ^ _06274_;
	assign _06286_ = _06285_ ^ _06260_;
	assign _06287_ = _06286_ ^ _06252_;
	assign _06288_ = _06287_ ^ _06240_;
	assign _06289_ = _06288_ | _06238_;
	assign _06290_ = _06289_ | _03810_;
	assign _06292_ = _06237_ ^ _03052_;
	assign _06293_ = ~(_06292_ & _06288_);
	assign _06294_ = _03832_ & ~_06293_;
	assign _06295_ = _06290_ & ~_06294_;
	assign _06296_ = _06292_ | _06288_;
	assign _06297_ = _03876_ & ~_06296_;
	assign _06298_ = _06295_ & ~_06297_;
	assign _06299_ = _06288_ & ~_06292_;
	assign _06300_ = (_06299_ ? _04241_ : _06298_);
	assign _06301_ = \mchip.wrapper.intxtReg.Q [7] ^ \mchip.wrapper.keyReg.Q [7];
	assign _06303_ = _06301_ ^ _06300_;
	assign _06304_ = _06303_ ^ _06190_;
	assign _06305_ = _06304_ ^ _05900_;
	assign _06306_ = _06305_ ^ _04822_;
	assign _06307_ = _06306_ ^ _03184_;
	assign _06308_ = ~_03140_;
	assign _06309_ = _06308_ & ~_04723_;
	assign _06310_ = _04745_ & _03129_;
	assign _06311_ = ~(_06310_ | _06309_);
	assign _06312_ = _04778_ & ~_03096_;
	assign _06314_ = _06311_ & ~_06312_;
	assign _06315_ = (_04810_ ? _03107_ : _06314_);
	assign _06316_ = _05801_ | _03305_;
	assign _06317_ = _05824_ & ~_03294_;
	assign _06318_ = _06316_ & ~_06317_;
	assign _06319_ = _05856_ & ~_04438_;
	assign _06320_ = _06318_ & ~_06319_;
	assign _06321_ = (_05889_ ? _04471_ : _06320_);
	assign _06322_ = _06179_ | _03305_;
	assign _06323_ = _03294_ & ~_06182_;
	assign _06325_ = _06322_ & ~_06323_;
	assign _06326_ = _03283_ & ~_06186_;
	assign _06327_ = _06325_ & ~_06326_;
	assign _06328_ = (_06189_ ? _04558_ : _06327_);
	assign _06329_ = _06289_ | _01835_;
	assign _06330_ = _03294_ & ~_06293_;
	assign _06331_ = _06329_ & ~_06330_;
	assign _06332_ = _03283_ & ~_06296_;
	assign _06333_ = _06331_ & ~_06332_;
	assign _06334_ = (_06299_ ? _04558_ : _06333_);
	assign _06336_ = ~(\mchip.wrapper.intxtReg.Q [6] ^ \mchip.wrapper.keyReg.Q [6]);
	assign _06337_ = _06336_ ^ _06334_;
	assign _06338_ = _06337_ ^ _06328_;
	assign _06339_ = _06338_ ^ _06321_;
	assign _06340_ = _06339_ ^ _06315_;
	assign _06341_ = _03085_ ^ _03107_;
	assign _06342_ = _06341_ ^ \mchip.wrapper.keyReg.Q [14];
	assign _06343_ = _06342_ ^ _06340_;
	assign _06344_ = ~(_06343_ & _06307_);
	assign _06345_ = _06344_ | _03217_;
	assign _06347_ = _06343_ | ~_06307_;
	assign _06348_ = _03206_ & ~_06347_;
	assign _06349_ = _06345_ & ~_06348_;
	assign _06350_ = _06307_ | ~_06343_;
	assign _06351_ = _03162_ & ~_06350_;
	assign _06352_ = _06349_ & ~_06351_;
	assign _06353_ = ~(_06343_ | _06307_);
	assign _06354_ = (_06353_ ? _03195_ : _06352_);
	assign _06355_ = ~_03481_;
	assign _06356_ = _06355_ & ~_04723_;
	assign _06358_ = _04745_ & ~_04855_;
	assign _06359_ = ~(_06358_ | _06356_);
	assign _06360_ = _04778_ & ~_04888_;
	assign _06361_ = _06359_ & ~_06360_;
	assign _06362_ = (_04810_ ? _04833_ : _06361_);
	assign _06363_ = _05801_ | _04955_;
	assign _06364_ = _05824_ & ~_04944_;
	assign _06365_ = _06363_ & ~_06364_;
	assign _06366_ = _05856_ & ~_04999_;
	assign _06367_ = _06365_ & ~_06366_;
	assign _06369_ = (_05889_ ? _05032_ : _06367_);
	assign _06370_ = _06179_ | _02450_;
	assign _06371_ = ~_04944_;
	assign _06372_ = _06371_ & ~_06182_;
	assign _06373_ = _06370_ & ~_06372_;
	assign _06374_ = _04933_ & ~_06186_;
	assign _06375_ = _06373_ & ~_06374_;
	assign _06376_ = (_06189_ ? _05129_ : _06375_);
	assign _06377_ = _06289_ | _05152_;
	assign _06378_ = _04855_ & ~_06293_;
	assign _06380_ = _06377_ & ~_06378_;
	assign _06381_ = _03459_ & ~_06296_;
	assign _06382_ = _06380_ & ~_06381_;
	assign _06383_ = (_06299_ ? _01735_ : _06382_);
	assign _06384_ = ~(\mchip.wrapper.intxtReg.Q [5] ^ \mchip.wrapper.keyReg.Q [5]);
	assign _06385_ = _06384_ ^ _06383_;
	assign _06386_ = _06385_ ^ _06376_;
	assign _06387_ = _06386_ ^ _06369_;
	assign _06388_ = _06387_ ^ _06362_;
	assign _06389_ = _03459_ ^ _04833_;
	assign _06391_ = _06389_ ^ \mchip.wrapper.keyReg.Q [13];
	assign _06392_ = _06391_ ^ _06388_;
	assign _06393_ = ~_05348_;
	assign _06394_ = _06393_ & ~_04723_;
	assign _06395_ = _04745_ & ~_05371_;
	assign _06396_ = ~(_06395_ | _06394_);
	assign _06397_ = _04778_ & ~_05404_;
	assign _06398_ = _06396_ & ~_06397_;
	assign _06399_ = (_04810_ ? \mchip.wrapper.keyReg.Q [4] : _06398_);
	assign _06400_ = _05801_ | _03525_;
	assign _06402_ = _05824_ & ~_03514_;
	assign _06403_ = _06400_ & ~_06402_;
	assign _06404_ = _05856_ & ~_05482_;
	assign _06405_ = _06403_ & ~_06404_;
	assign _06406_ = (_05889_ ? _05515_ : _06405_);
	assign _06407_ = _06179_ | _05537_;
	assign _06408_ = _05371_ & ~_06182_;
	assign _06409_ = _06407_ & ~_06408_;
	assign _06410_ = _05326_ & ~_06186_;
	assign _06411_ = _06409_ & ~_06410_;
	assign _06413_ = (_06189_ ? _01110_ : _06411_);
	assign _06414_ = _06289_ | _05646_;
	assign _06415_ = ~_05635_;
	assign _06416_ = _06415_ & ~_06293_;
	assign _06417_ = _06414_ & ~_06416_;
	assign _06418_ = _05482_ & ~_06296_;
	assign _06419_ = _06417_ & ~_06418_;
	assign _06420_ = (_06299_ ? _05713_ : _06419_);
	assign _06421_ = ~(\mchip.wrapper.intxtReg.Q [4] ^ \mchip.wrapper.keyReg.Q [4]);
	assign _06422_ = _06421_ ^ _06420_;
	assign _06424_ = _06422_ ^ _06413_;
	assign _06425_ = _06424_ ^ _06406_;
	assign _06426_ = _06425_ ^ _06399_;
	assign _06427_ = _03525_ ^ _06426_;
	assign _06428_ = ~(_06427_ & _06392_);
	assign _06429_ = _06428_ | _03184_;
	assign _06430_ = _06427_ | ~_06392_;
	assign _06431_ = _03173_ & ~_06430_;
	assign _06432_ = _06429_ & ~_06431_;
	assign _06434_ = _06392_ | ~_06427_;
	assign _06435_ = _03162_ & ~_06434_;
	assign _06436_ = _06432_ & ~_06435_;
	assign _06437_ = ~(_06427_ | _06392_);
	assign _06438_ = (_06437_ ? _03667_ : _06436_);
	assign _06439_ = _05945_ | _04723_;
	assign _06440_ = _04745_ & ~_00271_;
	assign _06441_ = _06439_ & ~_06440_;
	assign _06442_ = _04778_ & ~_05911_;
	assign _06443_ = _06441_ & ~_06442_;
	assign _06445_ = (_04810_ ? _03733_ : _06443_);
	assign _06446_ = _05945_ | _05801_;
	assign _06447_ = _05824_ & ~_03755_;
	assign _06448_ = _06446_ & ~_06447_;
	assign _06449_ = _05856_ & ~_05911_;
	assign _06450_ = _06448_ & ~_06449_;
	assign _06451_ = (_05889_ ? _06099_ : _06450_);
	assign _06452_ = _06179_ | _05945_;
	assign _06453_ = _00271_ & ~_06182_;
	assign _06454_ = _06452_ & ~_06453_;
	assign _06456_ = _05911_ & ~_06186_;
	assign _06457_ = _06454_ & ~_06456_;
	assign _06458_ = (_06189_ ? _06108_ : _06457_);
	assign _06459_ = _06289_ | _06113_;
	assign _06460_ = _06111_ & ~_06293_;
	assign _06461_ = _06459_ & ~_06460_;
	assign _06462_ = ~_06110_;
	assign _06463_ = _06462_ & ~_06296_;
	assign _06464_ = _06461_ & ~_06463_;
	assign _06465_ = (_06299_ ? _02616_ : _06464_);
	assign _00000_ = _06099_ ^ _03777_;
	assign _00001_ = _00000_ ^ _06465_;
	assign _00002_ = _00001_ ^ _06458_;
	assign _00003_ = _00002_ ^ _06451_;
	assign _00004_ = _00003_ ^ _06445_;
	assign _00005_ = _00004_ ^ _05945_;
	assign _00006_ = _06134_ | _04723_;
	assign _00007_ = _04745_ & ~_06136_;
	assign _00008_ = _00006_ & ~_00007_;
	assign _00009_ = _04778_ & ~_06139_;
	assign _00011_ = _00008_ & ~_00009_;
	assign _00012_ = (_04810_ ? _06129_ : _00011_);
	assign _00013_ = _06146_ | _05801_;
	assign _00014_ = _05824_ & ~_06136_;
	assign _00015_ = _00013_ & ~_00014_;
	assign _00016_ = _05856_ & ~_06139_;
	assign _00017_ = _00015_ & ~_00016_;
	assign _00018_ = (_05889_ ? _01188_ : _00017_);
	assign _00019_ = _06179_ | _06134_;
	assign _00020_ = _06131_ & ~_06182_;
	assign _00022_ = _00019_ & ~_00020_;
	assign _00023_ = _06130_ & ~_06186_;
	assign _00024_ = _00022_ & ~_00023_;
	assign _00025_ = (_06189_ ? _06160_ : _00024_);
	assign _00026_ = _06289_ | _06163_;
	assign _00027_ = _06162_ & ~_06293_;
	assign _00028_ = _00026_ & ~_00027_;
	assign _00029_ = _06139_ & ~_06296_;
	assign _00030_ = _00028_ & ~_00029_;
	assign _00031_ = (_06299_ ? _01188_ : _00030_);
	assign _00033_ = \mchip.wrapper.keyReg.Q [2] ^ \mchip.wrapper.intxtReg.Q [2];
	assign _00034_ = _00033_ ^ _00031_;
	assign _00035_ = _00034_ ^ _00025_;
	assign _00036_ = _00035_ ^ _00018_;
	assign _00037_ = _00036_ ^ _00012_;
	assign _00038_ = _00037_ ^ _06134_;
	assign _00039_ = _00038_ | _00005_;
	assign _00040_ = _00039_ | _03810_;
	assign _00041_ = _00004_ ^ _05934_;
	assign _00042_ = ~(_00041_ & _00038_);
	assign _00044_ = _03239_ & ~_00042_;
	assign _00045_ = _00040_ & ~_00044_;
	assign _00046_ = _00041_ | _00038_;
	assign _00047_ = _03228_ & ~_00046_;
	assign _00048_ = _00045_ & ~_00047_;
	assign _00049_ = _00038_ & ~_00041_;
	assign _00050_ = (_00049_ ? _00996_ : _00048_);
	assign _00052_ = ~_00051_;
	assign _00053_ = _04723_ | ~_03074_;
	assign _00055_ = _04745_ & ~_03063_;
	assign _00056_ = _00053_ & ~_00055_;
	assign _00057_ = _04778_ & ~_06191_;
	assign _00058_ = _00056_ & ~_00057_;
	assign _00059_ = (_04810_ ? \mchip.wrapper.keyReg.Q [1] : _00058_);
	assign _00060_ = _06202_ | _05801_;
	assign _00061_ = _05824_ & ~_06201_;
	assign _00062_ = _00060_ & ~_00061_;
	assign _00063_ = _05856_ & ~_06206_;
	assign _00064_ = _00062_ & ~_00063_;
	assign _00066_ = (_05889_ ? _06211_ : _00064_);
	assign _00067_ = _06179_ | _03074_;
	assign _00068_ = _03063_ & ~_06182_;
	assign _00069_ = _00067_ & ~_00068_;
	assign _00070_ = _03052_ & ~_06186_;
	assign _00071_ = _00069_ & ~_00070_;
	assign _00072_ = (_06189_ ? _06220_ : _00071_);
	assign _00073_ = _06289_ | _06223_;
	assign _00074_ = _06222_ & ~_06293_;
	assign _00075_ = _00073_ & ~_00074_;
	assign _00077_ = _06206_ & ~_06296_;
	assign _00078_ = _00075_ & ~_00077_;
	assign _00079_ = (_06299_ ? _06231_ : _00078_);
	assign _00080_ = \mchip.wrapper.keyReg.Q [1] ^ \mchip.wrapper.intxtReg.Q [1];
	assign _00081_ = _00080_ ^ _00079_;
	assign _00082_ = _00081_ ^ _00072_;
	assign _00083_ = _00082_ ^ _00066_;
	assign _00084_ = _00083_ ^ _00059_;
	assign _00085_ = _00084_ ^ _00052_;
	assign _00088_ = ~_00086_;
	assign _00089_ = ~_06243_;
	assign _00090_ = _04723_ | ~_00089_;
	assign _00091_ = _04745_ & ~_06245_;
	assign _00092_ = _00090_ & ~_00091_;
	assign _00093_ = _04778_ & ~_06248_;
	assign _00094_ = _00092_ & ~_00093_;
	assign _00095_ = (_04810_ ? \mchip.wrapper.keyReg.Q [0] : _00094_);
	assign _00096_ = _05801_ | _00086_;
	assign _00097_ = _05824_ & ~_03963_;
	assign _00099_ = _00096_ & ~_00097_;
	assign _00100_ = _05856_ & ~_06240_;
	assign _00101_ = _00099_ & ~_00100_;
	assign _00102_ = (_05889_ ? _06259_ : _00101_);
	assign _00103_ = _02279_ | _06179_;
	assign _00104_ = _06263_ & ~_06182_;
	assign _00105_ = _00103_ & ~_00104_;
	assign _00106_ = _06248_ & ~_06186_;
	assign _00107_ = _00105_ & ~_00106_;
	assign _00108_ = (_06189_ ? _06273_ : _00107_);
	assign _00110_ = _06289_ | _06264_;
	assign _00111_ = _06266_ & ~_06293_;
	assign _00112_ = _00110_ & ~_00111_;
	assign _00113_ = _06248_ & ~_06296_;
	assign _00114_ = _00112_ & ~_00113_;
	assign _00115_ = (_06299_ ? _06280_ : _00114_);
	assign _00116_ = \mchip.wrapper.keyReg.Q [0] ^ \mchip.wrapper.intxtReg.Q [0];
	assign _00117_ = _00116_ ^ _00115_;
	assign _00118_ = _00117_ ^ _00108_;
	assign _00119_ = _00118_ ^ _00102_;
	assign _00121_ = _00119_ ^ _00095_;
	assign _00122_ = _00121_ ^ _00088_;
	assign _00123_ = _00122_ | _00085_;
	assign _00124_ = _00123_ | _03810_;
	assign _00125_ = _00084_ ^ _00051_;
	assign _00126_ = ~(_00125_ & _00122_);
	assign _00127_ = _03832_ & ~_00126_;
	assign _00128_ = _00124_ & ~_00127_;
	assign _00129_ = _00125_ | _00122_;
	assign _00130_ = _03876_ & ~_00129_;
	assign _00132_ = _00128_ & ~_00130_;
	assign _00133_ = _00122_ & ~_00125_;
	assign _00134_ = (_00133_ ? _04241_ : _00132_);
	assign _00135_ = _04318_ ^ _03173_;
	assign _00136_ = _00135_ ^ _00134_;
	assign _00137_ = _00136_ ^ _00050_;
	assign _00138_ = _00137_ ^ _06438_;
	assign _00139_ = _00138_ ^ _06354_;
	assign _00140_ = _00139_ ^ _03162_;
	assign _00141_ = _06344_ | _03140_;
	assign _00143_ = _03129_ & ~_06347_;
	assign _00144_ = _00141_ & ~_00143_;
	assign _00145_ = _03085_ & ~_06350_;
	assign _00146_ = _00144_ & ~_00145_;
	assign _00147_ = (_06353_ ? _03107_ : _00146_);
	assign _00148_ = _06428_ | _03305_;
	assign _00149_ = _04503_ & ~_06430_;
	assign _00150_ = _00148_ & ~_00149_;
	assign _00151_ = _03283_ & ~_06434_;
	assign _00152_ = _00150_ & ~_00151_;
	assign _00154_ = (_06437_ ? _04471_ : _00152_);
	assign _00155_ = _00039_ | _03305_;
	assign _00156_ = _03294_ & ~_00042_;
	assign _00157_ = _00155_ & ~_00156_;
	assign _00158_ = _03283_ & ~_00046_;
	assign _00159_ = _00157_ & ~_00158_;
	assign _00160_ = (_00049_ ? _04558_ : _00159_);
	assign _00161_ = _00123_ | _01835_;
	assign _00162_ = _03294_ & ~_00126_;
	assign _00163_ = _00161_ & ~_00162_;
	assign _00165_ = _03283_ & ~_00129_;
	assign _00166_ = _00163_ & ~_00165_;
	assign _00167_ = (_00133_ ? _04558_ : _00166_);
	assign _00168_ = _06341_ ^ _04712_;
	assign _00169_ = _00168_ ^ _00167_;
	assign _00170_ = _00169_ ^ _00160_;
	assign _00171_ = _00170_ ^ _00154_;
	assign _00172_ = _00171_ ^ _00147_;
	assign _00173_ = _00172_ ^ _03085_;
	assign _00174_ = ~(_00173_ & _00140_);
	assign _00176_ = _00174_ | _03217_;
	assign _00177_ = _00173_ | ~_00140_;
	assign _00178_ = _03206_ & ~_00177_;
	assign _00179_ = _00176_ & ~_00178_;
	assign _00180_ = _00140_ | ~_00173_;
	assign _00181_ = _03162_ & ~_00180_;
	assign _00182_ = _00179_ & ~_00181_;
	assign _00183_ = ~(_00173_ | _00140_);
	assign _00184_ = (_00183_ ? _03195_ : _00182_);
	assign _00185_ = _06344_ | _03481_;
	assign _00187_ = _03470_ & ~_06347_;
	assign _00188_ = _00185_ & ~_00187_;
	assign _00189_ = _03459_ & ~_06350_;
	assign _00190_ = _00188_ & ~_00189_;
	assign _00191_ = (_06353_ ? _04833_ : _00190_);
	assign _00192_ = _06428_ | _04955_;
	assign _00193_ = _06371_ & ~_06430_;
	assign _00194_ = _00192_ & ~_00193_;
	assign _00195_ = _04933_ & ~_06434_;
	assign _00196_ = _00194_ & ~_00195_;
	assign _00198_ = (_06437_ ? _05032_ : _00196_);
	assign _00199_ = _00039_ | _02450_;
	assign _00200_ = _06371_ & ~_00042_;
	assign _00201_ = _00199_ & ~_00200_;
	assign _00202_ = _04933_ & ~_00046_;
	assign _00203_ = _00201_ & ~_00202_;
	assign _00204_ = (_00049_ ? _05129_ : _00203_);
	assign _00205_ = _00123_ | _05152_;
	assign _00206_ = _04855_ & ~_00126_;
	assign _00207_ = _00205_ & ~_00206_;
	assign _00209_ = _03459_ & ~_00129_;
	assign _00210_ = _00207_ & ~_00209_;
	assign _00211_ = (_00133_ ? _01735_ : _00210_);
	assign _00212_ = _06389_ ^ _05304_;
	assign _00213_ = _00212_ ^ _00211_;
	assign _00214_ = _00213_ ^ _00204_;
	assign _00215_ = _00214_ ^ _00198_;
	assign _00216_ = _00215_ ^ _00191_;
	assign _00217_ = _00216_ ^ _03459_;
	assign _00218_ = _06344_ | _05348_;
	assign _00220_ = _05337_ & ~_06347_;
	assign _00221_ = _00218_ & ~_00220_;
	assign _00222_ = _05326_ & ~_06350_;
	assign _00223_ = _00221_ & ~_00222_;
	assign _00224_ = (_06353_ ? \mchip.wrapper.keyReg.Q [4] : _00223_);
	assign _00225_ = _06428_ | _03525_;
	assign _00226_ = ~_03514_;
	assign _00227_ = _00226_ & ~_06430_;
	assign _00228_ = _00225_ & ~_00227_;
	assign _00229_ = _03503_ & ~_06434_;
	assign _00231_ = _00228_ & ~_00229_;
	assign _00232_ = (_06437_ ? _05515_ : _00231_);
	assign _00233_ = _00039_ | _05537_;
	assign _00234_ = _05371_ & ~_00042_;
	assign _00235_ = _00233_ & ~_00234_;
	assign _00236_ = _05326_ & ~_00046_;
	assign _00237_ = _00235_ & ~_00236_;
	assign _00238_ = (_00049_ ? _01110_ : _00237_);
	assign _00239_ = _00123_ | _05646_;
	assign _00240_ = _06415_ & ~_00126_;
	assign _00242_ = _00239_ & ~_00240_;
	assign _00243_ = _05482_ & ~_00129_;
	assign _00244_ = _00242_ & ~_00243_;
	assign _00245_ = (_00133_ ? _05713_ : _00244_);
	assign _00246_ = _05790_ ^ _03514_;
	assign _00247_ = _00246_ ^ _00245_;
	assign _00248_ = _00247_ ^ _00238_;
	assign _00249_ = _00248_ ^ _00232_;
	assign _00250_ = _00249_ ^ _00224_;
	assign _00251_ = _00250_ ^ _03503_;
	assign _00253_ = ~(_00251_ & _00217_);
	assign _00254_ = _00253_ | _03184_;
	assign _00255_ = _00251_ | ~_00217_;
	assign _00256_ = _03173_ & ~_00255_;
	assign _00257_ = _00254_ & ~_00256_;
	assign _00258_ = _00217_ | ~_00251_;
	assign _00259_ = _03162_ & ~_00258_;
	assign _00260_ = _00257_ & ~_00259_;
	assign _00261_ = ~(_00251_ | _00217_);
	assign _00262_ = (_00261_ ? _03667_ : _00260_);
	assign _00264_ = _06344_ | _05945_;
	assign _00265_ = _03755_ & ~_06347_;
	assign _00266_ = _00264_ & ~_00265_;
	assign _00267_ = _03744_ & ~_06350_;
	assign _00268_ = _00266_ & ~_00267_;
	assign _00269_ = (_06353_ ? _03733_ : _00268_);
	assign _00270_ = _06428_ | _05945_;
	assign _00272_ = _00271_ & ~_06430_;
	assign _00273_ = _00270_ & ~_00272_;
	assign _00275_ = _03744_ & ~_06434_;
	assign _00276_ = _00273_ & ~_00275_;
	assign _00277_ = (_06437_ ? _06099_ : _00276_);
	assign _00278_ = _00039_ | _05945_;
	assign _00279_ = _00271_ & ~_00042_;
	assign _00280_ = _00278_ & ~_00279_;
	assign _00281_ = _05911_ & ~_00046_;
	assign _00282_ = _00280_ & ~_00281_;
	assign _00283_ = (_00049_ ? _06108_ : _00282_);
	assign _00284_ = _00123_ | _06113_;
	assign _00286_ = _06111_ & ~_00126_;
	assign _00287_ = _00284_ & ~_00286_;
	assign _00288_ = _06462_ & ~_00129_;
	assign _00289_ = _00287_ & ~_00288_;
	assign _00290_ = (_00133_ ? _02616_ : _00289_);
	assign _00291_ = _06127_ ^ _00271_;
	assign _00292_ = _00291_ ^ _00290_;
	assign _00293_ = _00292_ ^ _00283_;
	assign _00294_ = _00293_ ^ _00277_;
	assign _00295_ = _00294_ ^ _00269_;
	assign _00297_ = _00295_ ^ _05911_;
	assign _00298_ = _06344_ | _06134_;
	assign _00299_ = _06131_ & ~_06347_;
	assign _00300_ = _00298_ & ~_00299_;
	assign _00301_ = _06130_ & ~_06350_;
	assign _00302_ = _00300_ & ~_00301_;
	assign _00303_ = (_06353_ ? _06129_ : _00302_);
	assign _00304_ = _06428_ | _06146_;
	assign _00305_ = _06131_ & ~_06430_;
	assign _00306_ = _00304_ & ~_00305_;
	assign _00308_ = _06130_ & ~_06434_;
	assign _00309_ = _00306_ & ~_00308_;
	assign _00310_ = (_06437_ ? _01188_ : _00309_);
	assign _00311_ = _00039_ | _06134_;
	assign _00312_ = _06131_ & ~_00042_;
	assign _00313_ = _00311_ & ~_00312_;
	assign _00314_ = _06130_ & ~_00046_;
	assign _00315_ = _00313_ & ~_00314_;
	assign _00316_ = (_00049_ ? _06160_ : _00315_);
	assign _00317_ = _00123_ | _06163_;
	assign _00319_ = _06162_ & ~_00126_;
	assign _00320_ = _00317_ & ~_00319_;
	assign _00321_ = _06139_ & ~_00129_;
	assign _00322_ = _00320_ & ~_00321_;
	assign _00323_ = (_00133_ ? _01188_ : _00322_);
	assign _00324_ = _06181_ ^ _06131_;
	assign _00325_ = _00324_ ^ _00323_;
	assign _00326_ = _00325_ ^ _00316_;
	assign _00327_ = _00326_ ^ _00310_;
	assign _00328_ = _00327_ ^ _00303_;
	assign _00330_ = _00328_ ^ _06139_;
	assign _00331_ = _00330_ | _00297_;
	assign _00332_ = _00331_ | _03810_;
	assign _00333_ = _00328_ ^ _06130_;
	assign _00334_ = _00297_ | _00333_;
	assign _00335_ = _03239_ & ~_00334_;
	assign _00336_ = _00332_ & ~_00335_;
	assign _00337_ = ~(_00297_ & _00333_);
	assign _00338_ = _03228_ & ~_00337_;
	assign _00340_ = _00336_ & ~_00338_;
	assign _00341_ = _00297_ & ~_00333_;
	assign _00342_ = (_00341_ ? _00996_ : _00340_);
	assign _00343_ = _06344_ | _06192_;
	assign _00345_ = _00344_ & ~_06347_;
	assign _00346_ = _00343_ & ~_00345_;
	assign _00347_ = _03052_ & ~_06350_;
	assign _00348_ = _00346_ & ~_00347_;
	assign _00349_ = (_06353_ ? \mchip.wrapper.keyReg.Q [1] : _00348_);
	assign _00351_ = _06428_ | _06202_;
	assign _00352_ = ~_06201_;
	assign _00353_ = _00352_ & ~_06430_;
	assign _00354_ = _00351_ & ~_00353_;
	assign _00355_ = _06200_ & ~_06434_;
	assign _00356_ = _00354_ & ~_00355_;
	assign _00357_ = (_06437_ ? _06211_ : _00356_);
	assign _00358_ = _00039_ | _03074_;
	assign _00359_ = _03063_ & ~_00042_;
	assign _00360_ = _00358_ & ~_00359_;
	assign _00362_ = _03052_ & ~_00046_;
	assign _00363_ = _00360_ & ~_00362_;
	assign _00364_ = (_00049_ ? _06220_ : _00363_);
	assign _00365_ = _00123_ | _06223_;
	assign _00366_ = _06222_ & ~_00126_;
	assign _00367_ = _00365_ & ~_00366_;
	assign _00368_ = _06206_ & ~_00129_;
	assign _00369_ = _00367_ & ~_00368_;
	assign _00370_ = (_00133_ ? _06231_ : _00369_);
	assign _00371_ = _06238_ ^ _03063_;
	assign _00373_ = _00371_ ^ _00370_;
	assign _00374_ = _00373_ ^ _00364_;
	assign _00375_ = _00374_ ^ _00357_;
	assign _00376_ = _00375_ ^ _00349_;
	assign _00377_ = _00376_ ^ _06191_;
	assign _00378_ = _06344_ | _06243_;
	assign _00379_ = _06242_ & ~_06347_;
	assign _00380_ = _00378_ & ~_00379_;
	assign _00381_ = _06241_ & ~_06350_;
	assign _00382_ = _00380_ & ~_00381_;
	assign _00384_ = (_06353_ ? \mchip.wrapper.keyReg.Q [0] : _00382_);
	assign _00385_ = _06428_ | _00086_;
	assign _00386_ = ~_03963_;
	assign _00387_ = _00386_ & ~_06430_;
	assign _00388_ = _00385_ & ~_00387_;
	assign _00389_ = _03952_ & ~_06434_;
	assign _00390_ = _00388_ & ~_00389_;
	assign _00391_ = (_06437_ ? _06259_ : _00390_);
	assign _00392_ = _00039_ | _02279_;
	assign _00393_ = _06263_ & ~_00042_;
	assign _00395_ = _00392_ & ~_00393_;
	assign _00396_ = _06248_ & ~_00046_;
	assign _00397_ = _00395_ & ~_00396_;
	assign _00398_ = (_00049_ ? _06273_ : _00397_);
	assign _00399_ = _00123_ | _06264_;
	assign _00400_ = _06266_ & ~_00126_;
	assign _00401_ = _00399_ & ~_00400_;
	assign _00402_ = _06248_ & ~_00129_;
	assign _00403_ = _00401_ & ~_00402_;
	assign _00404_ = (_00133_ ? _06280_ : _00403_);
	assign _00406_ = _06288_ ^ _00386_;
	assign _00407_ = _00406_ ^ _00404_;
	assign _00408_ = _00407_ ^ _00398_;
	assign _00409_ = _00408_ ^ _00391_;
	assign _00410_ = _00409_ ^ _00384_;
	assign _00411_ = _00410_ ^ _06240_;
	assign _00412_ = _00411_ | _00377_;
	assign _00413_ = _00412_ | _03810_;
	assign _00414_ = _00410_ ^ _03952_;
	assign _00416_ = _00377_ | _00414_;
	assign _00417_ = _03832_ & ~_00416_;
	assign _00418_ = _00413_ & ~_00417_;
	assign _00419_ = _00376_ ^ _03052_;
	assign _00420_ = _00419_ | _00411_;
	assign _00421_ = _03876_ & ~_00420_;
	assign _00422_ = _00418_ & ~_00421_;
	assign _00423_ = _00411_ & ~_00419_;
	assign _00424_ = (_00423_ ? _04241_ : _00422_);
	assign _00425_ = _06307_ ^ \mchip.wrapper.keyReg.Q [7];
	assign _00427_ = _00425_ ^ _00424_;
	assign _00428_ = _00427_ ^ _00342_;
	assign _00429_ = _00428_ ^ _00262_;
	assign _00430_ = _00429_ ^ _00184_;
	assign _00431_ = _00430_ ^ _03250_;
	assign _00432_ = _00174_ | _03140_;
	assign _00433_ = _03129_ & ~_00177_;
	assign _00434_ = _00432_ & ~_00433_;
	assign _00435_ = _03085_ & ~_00180_;
	assign _00436_ = _00434_ & ~_00435_;
	assign _00438_ = (_00183_ ? _03107_ : _00436_);
	assign _00439_ = _00253_ | _03305_;
	assign _00440_ = _04503_ & ~_00255_;
	assign _00441_ = _00439_ & ~_00440_;
	assign _00442_ = _03283_ & ~_00258_;
	assign _00443_ = _00441_ & ~_00442_;
	assign _00444_ = (_00261_ ? _04471_ : _00443_);
	assign _00445_ = _00331_ | _03305_;
	assign _00446_ = _03294_ & ~_00334_;
	assign _00447_ = _00445_ & ~_00446_;
	assign _00449_ = _03283_ & ~_00337_;
	assign _00450_ = _00447_ & ~_00449_;
	assign _00451_ = (_00341_ ? _04558_ : _00450_);
	assign _00452_ = _00412_ | _01835_;
	assign _00453_ = _03294_ & ~_00416_;
	assign _00454_ = _00452_ & ~_00453_;
	assign _00455_ = _03283_ & ~_00420_;
	assign _00456_ = _00454_ & ~_00455_;
	assign _00457_ = (_00423_ ? _04558_ : _00456_);
	assign _00458_ = _06343_ ^ \mchip.wrapper.keyReg.Q [6];
	assign _00460_ = _00458_ ^ _00457_;
	assign _00461_ = _00460_ ^ _00451_;
	assign _00462_ = _00461_ ^ _00444_;
	assign _00463_ = _00462_ ^ _00438_;
	assign _00464_ = _00463_ ^ _03305_;
	assign _00465_ = ~(_00464_ & _00431_);
	assign _00466_ = _00465_ | _03217_;
	assign _00467_ = _00464_ | ~_00431_;
	assign _00468_ = _03206_ & ~_00467_;
	assign _00469_ = _00466_ & ~_00468_;
	assign _00471_ = _00431_ | ~_00464_;
	assign _00472_ = _03162_ & ~_00471_;
	assign _00473_ = _00469_ & ~_00472_;
	assign _00474_ = ~(_00464_ | _00431_);
	assign _00475_ = (_00474_ ? _03195_ : _00473_);
	assign _00476_ = _00174_ | _03481_;
	assign _00477_ = _03470_ & ~_00177_;
	assign _00478_ = _00476_ & ~_00477_;
	assign _00479_ = _03459_ & ~_00180_;
	assign _00480_ = _00478_ & ~_00479_;
	assign _00482_ = (_00183_ ? _04833_ : _00480_);
	assign _00483_ = _00253_ | _04955_;
	assign _00484_ = _06371_ & ~_00255_;
	assign _00485_ = _00483_ & ~_00484_;
	assign _00486_ = _04933_ & ~_00258_;
	assign _00487_ = _00485_ & ~_00486_;
	assign _00488_ = (_00261_ ? _05032_ : _00487_);
	assign _00489_ = _00331_ | _02450_;
	assign _00490_ = _06371_ & ~_00334_;
	assign _00491_ = _00489_ & ~_00490_;
	assign _00493_ = _04933_ & ~_00337_;
	assign _00494_ = _00491_ & ~_00493_;
	assign _00495_ = (_00341_ ? _05129_ : _00494_);
	assign _00496_ = _00412_ | _05152_;
	assign _00497_ = _04855_ & ~_00416_;
	assign _00498_ = _00496_ & ~_00497_;
	assign _00499_ = _03459_ & ~_00420_;
	assign _00500_ = _00498_ & ~_00499_;
	assign _00501_ = (_00423_ ? _01735_ : _00500_);
	assign _00502_ = _06392_ ^ _04833_;
	assign _00504_ = _00502_ ^ _00501_;
	assign _00505_ = _00504_ ^ _00495_;
	assign _00506_ = _00505_ ^ _00488_;
	assign _00507_ = _00506_ ^ _00482_;
	assign _00508_ = _00507_ ^ _06355_;
	assign _00509_ = ~_03525_;
	assign _00510_ = _00174_ | _05348_;
	assign _00511_ = _05337_ & ~_00177_;
	assign _00512_ = _00510_ & ~_00511_;
	assign _00513_ = _05326_ & ~_00180_;
	assign _00515_ = _00512_ & ~_00513_;
	assign _00516_ = (_00183_ ? \mchip.wrapper.keyReg.Q [4] : _00515_);
	assign _00517_ = _00253_ | _03525_;
	assign _00518_ = _00226_ & ~_00255_;
	assign _00519_ = _00517_ & ~_00518_;
	assign _00520_ = _03503_ & ~_00258_;
	assign _00521_ = _00519_ & ~_00520_;
	assign _00522_ = (_00261_ ? _05515_ : _00521_);
	assign _00523_ = _00331_ | _05537_;
	assign _00524_ = _05371_ & ~_00334_;
	assign _00526_ = _00523_ & ~_00524_;
	assign _00527_ = _05326_ & ~_00337_;
	assign _00528_ = _00526_ & ~_00527_;
	assign _00529_ = (_00341_ ? _01110_ : _00528_);
	assign _00530_ = _00412_ | _05646_;
	assign _00531_ = _06415_ & ~_00416_;
	assign _00532_ = _00530_ & ~_00531_;
	assign _00533_ = _05482_ & ~_00420_;
	assign _00534_ = _00532_ & ~_00533_;
	assign _00535_ = (_00423_ ? _05713_ : _00534_);
	assign _00537_ = _06427_ ^ \mchip.wrapper.keyReg.Q [4];
	assign _00538_ = _00537_ ^ _00535_;
	assign _00539_ = _00538_ ^ _00529_;
	assign _00540_ = _00539_ ^ _00522_;
	assign _00541_ = _00540_ ^ _00516_;
	assign _00542_ = _00541_ ^ _00509_;
	assign _00543_ = ~(_00542_ & _00508_);
	assign _00544_ = _00543_ | _03184_;
	assign _00545_ = _00542_ | ~_00508_;
	assign _00546_ = _03173_ & ~_00545_;
	assign _00548_ = _00544_ & ~_00546_;
	assign _00549_ = _00508_ | ~_00542_;
	assign _00550_ = _03162_ & ~_00549_;
	assign _00551_ = _00548_ & ~_00550_;
	assign _00552_ = ~(_00542_ | _00508_);
	assign _00553_ = (_00552_ ? _03667_ : _00551_);
	assign _00554_ = ~_03766_;
	assign _00555_ = _00174_ | _05945_;
	assign _00556_ = _03755_ & ~_00177_;
	assign _00557_ = _00555_ & ~_00556_;
	assign _00559_ = _03744_ & ~_00180_;
	assign _00560_ = _00557_ & ~_00559_;
	assign _00561_ = (_00183_ ? _03733_ : _00560_);
	assign _00562_ = _00253_ | _05945_;
	assign _00563_ = _00271_ & ~_00255_;
	assign _00564_ = _00562_ & ~_00563_;
	assign _00565_ = _03744_ & ~_00258_;
	assign _00566_ = _00564_ & ~_00565_;
	assign _00567_ = (_00261_ ? _06099_ : _00566_);
	assign _00568_ = _00331_ | _05945_;
	assign _00570_ = _00271_ & ~_00334_;
	assign _00571_ = _00568_ & ~_00570_;
	assign _00572_ = _05911_ & ~_00337_;
	assign _00573_ = _00571_ & ~_00572_;
	assign _00574_ = (_00341_ ? _06108_ : _00573_);
	assign _00575_ = _00412_ | _06113_;
	assign _00576_ = _06111_ & ~_00416_;
	assign _00577_ = _00575_ & ~_00576_;
	assign _00578_ = _06462_ & ~_00420_;
	assign _00579_ = _00577_ & ~_00578_;
	assign _00581_ = (_00423_ ? _02616_ : _00579_);
	assign _00582_ = _00005_ ^ _03733_;
	assign _00583_ = _00582_ ^ _00581_;
	assign _00584_ = _00583_ ^ _00574_;
	assign _00585_ = _00584_ ^ _00567_;
	assign _00586_ = _00585_ ^ _00561_;
	assign _00587_ = _00586_ ^ _00554_;
	assign _00588_ = ~_03711_;
	assign _00589_ = _00174_ | _06134_;
	assign _00590_ = _06131_ & ~_00177_;
	assign _00592_ = _00589_ & ~_00590_;
	assign _00593_ = _06130_ & ~_00180_;
	assign _00594_ = _00592_ & ~_00593_;
	assign _00595_ = (_00183_ ? _06129_ : _00594_);
	assign _00596_ = _00253_ | _06146_;
	assign _00597_ = _06131_ & ~_00255_;
	assign _00598_ = _00596_ & ~_00597_;
	assign _00599_ = _06130_ & ~_00258_;
	assign _00600_ = _00598_ & ~_00599_;
	assign _00601_ = (_00261_ ? _01188_ : _00600_);
	assign _00603_ = _00331_ | _06134_;
	assign _00604_ = _06131_ & ~_00334_;
	assign _00605_ = _00603_ & ~_00604_;
	assign _00606_ = _06130_ & ~_00337_;
	assign _00607_ = _00605_ & ~_00606_;
	assign _00608_ = (_00341_ ? _06160_ : _00607_);
	assign _00609_ = _00412_ | _06163_;
	assign _00610_ = _06162_ & ~_00416_;
	assign _00611_ = _00609_ & ~_00610_;
	assign _00612_ = _06139_ & ~_00420_;
	assign _00614_ = _00611_ & ~_00612_;
	assign _00615_ = (_00423_ ? _01188_ : _00614_);
	assign _00616_ = _00038_ ^ \mchip.wrapper.keyReg.Q [2];
	assign _00617_ = _00616_ ^ _00615_;
	assign _00618_ = _00617_ ^ _00608_;
	assign _00619_ = _00618_ ^ _00601_;
	assign _00620_ = _00619_ ^ _00595_;
	assign _00621_ = _00620_ ^ _00588_;
	assign _00622_ = _00621_ | _00587_;
	assign _00623_ = _00622_ | _03810_;
	assign _00625_ = _00586_ ^ _03766_;
	assign _00626_ = ~(_00625_ & _00621_);
	assign _00627_ = _03239_ & ~_00626_;
	assign _00628_ = _00623_ & ~_00627_;
	assign _00629_ = _00625_ | _00621_;
	assign _00630_ = _03228_ & ~_00629_;
	assign _00631_ = _00628_ & ~_00630_;
	assign _00632_ = _00621_ & ~_00625_;
	assign _00633_ = (_00632_ ? _00996_ : _00631_);
	assign _00634_ = _00174_ | _06192_;
	assign _00636_ = _00344_ & ~_00177_;
	assign _00637_ = _00634_ & ~_00636_;
	assign _00638_ = _03052_ & ~_00180_;
	assign _00639_ = _00637_ & ~_00638_;
	assign _00640_ = (_00183_ ? \mchip.wrapper.keyReg.Q [1] : _00639_);
	assign _00641_ = _00253_ | _06202_;
	assign _00642_ = _00352_ & ~_00255_;
	assign _00643_ = _00641_ & ~_00642_;
	assign _00644_ = _06200_ & ~_00258_;
	assign _00645_ = _00643_ & ~_00644_;
	assign _00647_ = (_00261_ ? _06211_ : _00645_);
	assign _00648_ = _00331_ | _03074_;
	assign _00649_ = _03063_ & ~_00334_;
	assign _00650_ = _00648_ & ~_00649_;
	assign _00651_ = _03052_ & ~_00337_;
	assign _00652_ = _00650_ & ~_00651_;
	assign _00653_ = (_00341_ ? _06220_ : _00652_);
	assign _00654_ = _00412_ | _06223_;
	assign _00655_ = _06222_ & ~_00416_;
	assign _00656_ = _00654_ & ~_00655_;
	assign _00658_ = _06206_ & ~_00420_;
	assign _00659_ = _00656_ & ~_00658_;
	assign _00660_ = (_00423_ ? _06231_ : _00659_);
	assign _00661_ = _00085_ ^ _03041_;
	assign _00662_ = _00661_ ^ _00660_;
	assign _00663_ = _00662_ ^ _00653_;
	assign _00664_ = _00663_ ^ _00647_;
	assign _00665_ = _00664_ ^ _00640_;
	assign _00666_ = _00665_ ^ _03074_;
	assign _00667_ = _00174_ | _06243_;
	assign _00669_ = _06242_ & ~_00177_;
	assign _00670_ = _00667_ & ~_00669_;
	assign _00671_ = _06241_ & ~_00180_;
	assign _00672_ = _00670_ & ~_00671_;
	assign _00673_ = (_00183_ ? \mchip.wrapper.keyReg.Q [0] : _00672_);
	assign _00674_ = _00253_ | _00086_;
	assign _00675_ = _00386_ & ~_00255_;
	assign _00676_ = _00674_ & ~_00675_;
	assign _00677_ = _03952_ & ~_00258_;
	assign _00678_ = _00676_ & ~_00677_;
	assign _00680_ = (_00261_ ? _06259_ : _00678_);
	assign _00681_ = _00331_ | _02279_;
	assign _00682_ = _06263_ & ~_00334_;
	assign _00683_ = _00681_ & ~_00682_;
	assign _00684_ = _06248_ & ~_00337_;
	assign _00685_ = _00683_ & ~_00684_;
	assign _00686_ = (_00341_ ? _06273_ : _00685_);
	assign _00687_ = _00412_ | _06264_;
	assign _00688_ = _06266_ & ~_00416_;
	assign _00689_ = _00687_ & ~_00688_;
	assign _00691_ = _06248_ & ~_00420_;
	assign _00692_ = _00689_ & ~_00691_;
	assign _00693_ = (_00423_ ? _06280_ : _00692_);
	assign _00694_ = _00122_ ^ _06262_;
	assign _00695_ = _00694_ ^ _00693_;
	assign _00696_ = _00695_ ^ _00686_;
	assign _00697_ = _00696_ ^ _00680_;
	assign _00698_ = _00697_ ^ _00673_;
	assign _00699_ = _00698_ ^ _00086_;
	assign _00700_ = _00699_ | _00666_;
	assign _00702_ = _00700_ | _03810_;
	assign _00703_ = _00665_ ^ _00051_;
	assign _00704_ = ~(_00703_ & _00699_);
	assign _00705_ = _03832_ & ~_00704_;
	assign _00706_ = _00702_ & ~_00705_;
	assign _00707_ = _00703_ | _00699_;
	assign _00708_ = _03876_ & ~_00707_;
	assign _00709_ = _00706_ & ~_00708_;
	assign _00710_ = _00699_ & ~_00703_;
	assign _00711_ = (_00710_ ? _04241_ : _00709_);
	assign _00713_ = _00140_ ^ _03239_;
	assign _00714_ = _00713_ ^ _00711_;
	assign _00715_ = _00714_ ^ _00633_;
	assign _00716_ = _00715_ ^ _00553_;
	assign _00717_ = _00716_ ^ _00475_;
	assign _00718_ = _00717_ ^ _03228_;
	assign _00719_ = _00465_ | _03140_;
	assign _00720_ = _03129_ & ~_00467_;
	assign _00721_ = _00719_ & ~_00720_;
	assign _00722_ = _03085_ & ~_00471_;
	assign _00724_ = _00721_ & ~_00722_;
	assign _00725_ = (_00474_ ? _03107_ : _00724_);
	assign _00726_ = _00543_ | _03305_;
	assign _00727_ = _04503_ & ~_00545_;
	assign _00728_ = _00726_ & ~_00727_;
	assign _00729_ = _03283_ & ~_00549_;
	assign _00730_ = _00728_ & ~_00729_;
	assign _00731_ = (_00552_ ? _04471_ : _00730_);
	assign _00732_ = _00622_ | _03305_;
	assign _00733_ = _03294_ & ~_00626_;
	assign _00735_ = _00732_ & ~_00733_;
	assign _00736_ = _03283_ & ~_00629_;
	assign _00737_ = _00735_ & ~_00736_;
	assign _00738_ = (_00632_ ? _04558_ : _00737_);
	assign _00739_ = _00700_ | _01835_;
	assign _00740_ = _03294_ & ~_00704_;
	assign _00741_ = _00739_ & ~_00740_;
	assign _00742_ = _03283_ & ~_00707_;
	assign _00743_ = _00741_ & ~_00742_;
	assign _00744_ = (_00710_ ? _04558_ : _00743_);
	assign _00746_ = _00173_ ^ _03294_;
	assign _00747_ = _00746_ ^ _00744_;
	assign _00748_ = _00747_ ^ _00738_;
	assign _00749_ = _00748_ ^ _00731_;
	assign _00750_ = _00749_ ^ _00725_;
	assign _00751_ = _00750_ ^ _03283_;
	assign _00752_ = ~(_00751_ & _00718_);
	assign _00753_ = _00752_ | _03217_;
	assign _00754_ = _00751_ | ~_00718_;
	assign _00755_ = _03206_ & ~_00754_;
	assign _00757_ = _00753_ & ~_00755_;
	assign _00758_ = _00718_ | ~_00751_;
	assign _00759_ = _03162_ & ~_00758_;
	assign _00760_ = _00757_ & ~_00759_;
	assign _00761_ = ~(_00751_ | _00718_);
	assign _00762_ = (_00761_ ? _03195_ : _00760_);
	assign _00763_ = _00465_ | _03481_;
	assign _00764_ = _03470_ & ~_00467_;
	assign _00765_ = _00763_ & ~_00764_;
	assign _00766_ = _03459_ & ~_00471_;
	assign _00768_ = _00765_ & ~_00766_;
	assign _00769_ = (_00474_ ? _04833_ : _00768_);
	assign _00770_ = _00543_ | _04955_;
	assign _00771_ = _06371_ & ~_00545_;
	assign _00772_ = _00770_ & ~_00771_;
	assign _00773_ = _04933_ & ~_00549_;
	assign _00774_ = _00772_ & ~_00773_;
	assign _00775_ = (_00552_ ? _05032_ : _00774_);
	assign _00776_ = _00622_ | _02450_;
	assign _00777_ = _06371_ & ~_00626_;
	assign _00779_ = _00776_ & ~_00777_;
	assign _00780_ = _04933_ & ~_00629_;
	assign _00781_ = _00779_ & ~_00780_;
	assign _00782_ = (_00632_ ? _05129_ : _00781_);
	assign _00783_ = _00700_ | _05152_;
	assign _00784_ = _04855_ & ~_00704_;
	assign _00785_ = _00783_ & ~_00784_;
	assign _00786_ = _03459_ & ~_00707_;
	assign _00787_ = _00785_ & ~_00786_;
	assign _00788_ = (_00710_ ? _01735_ : _00787_);
	assign _00790_ = _00217_ ^ _03470_;
	assign _00791_ = _00790_ ^ _00788_;
	assign _00792_ = _00791_ ^ _00782_;
	assign _00793_ = _00792_ ^ _00775_;
	assign _00794_ = _00793_ ^ _00769_;
	assign _00795_ = _00794_ ^ _03459_;
	assign _00796_ = _00465_ | _05348_;
	assign _00797_ = _05337_ & ~_00467_;
	assign _00798_ = _00796_ & ~_00797_;
	assign _00799_ = _05326_ & ~_00471_;
	assign _00801_ = _00798_ & ~_00799_;
	assign _00802_ = (_00474_ ? \mchip.wrapper.keyReg.Q [4] : _00801_);
	assign _00803_ = _00543_ | _03525_;
	assign _00804_ = _00226_ & ~_00545_;
	assign _00805_ = _00803_ & ~_00804_;
	assign _00806_ = _03503_ & ~_00549_;
	assign _00807_ = _00805_ & ~_00806_;
	assign _00808_ = (_00552_ ? _05515_ : _00807_);
	assign _00809_ = _00622_ | _05537_;
	assign _00810_ = _05371_ & ~_00626_;
	assign _00812_ = _00809_ & ~_00810_;
	assign _00813_ = _05326_ & ~_00629_;
	assign _00814_ = _00812_ & ~_00813_;
	assign _00815_ = (_00632_ ? _01110_ : _00814_);
	assign _00816_ = _00700_ | _05646_;
	assign _00817_ = _06415_ & ~_00704_;
	assign _00818_ = _00816_ & ~_00817_;
	assign _00819_ = _05482_ & ~_00707_;
	assign _00820_ = _00818_ & ~_00819_;
	assign _00821_ = (_00710_ ? _05713_ : _00820_);
	assign _00823_ = _00251_ ^ _03514_;
	assign _00824_ = _00823_ ^ _00821_;
	assign _00825_ = _00824_ ^ _00815_;
	assign _00826_ = _00825_ ^ _00808_;
	assign _00827_ = _00826_ ^ _00802_;
	assign _00828_ = _00827_ ^ _03503_;
	assign _00829_ = ~(_00828_ & _00795_);
	assign _00830_ = _00829_ | _03184_;
	assign _00831_ = _00828_ | ~_00795_;
	assign _00832_ = _03173_ & ~_00831_;
	assign _00834_ = _00830_ & ~_00832_;
	assign _00835_ = _00795_ | ~_00828_;
	assign _00836_ = _03162_ & ~_00835_;
	assign _00837_ = _00834_ & ~_00836_;
	assign _00838_ = ~(_00828_ | _00795_);
	assign _00839_ = (_00838_ ? _03667_ : _00837_);
	assign _00840_ = _00465_ | _05945_;
	assign _00841_ = _03755_ & ~_00467_;
	assign _00842_ = _00840_ & ~_00841_;
	assign _00843_ = _03744_ & ~_00471_;
	assign _00845_ = _00842_ & ~_00843_;
	assign _00846_ = (_00474_ ? _03733_ : _00845_);
	assign _00847_ = _00543_ | _05945_;
	assign _00848_ = _00271_ & ~_00545_;
	assign _00849_ = _00847_ & ~_00848_;
	assign _00850_ = _03744_ & ~_00549_;
	assign _00851_ = _00849_ & ~_00850_;
	assign _00852_ = (_00552_ ? _06099_ : _00851_);
	assign _00853_ = _00622_ | _05945_;
	assign _00854_ = _00271_ & ~_00626_;
	assign _00856_ = _00853_ & ~_00854_;
	assign _00857_ = _05911_ & ~_00629_;
	assign _00858_ = _00856_ & ~_00857_;
	assign _00859_ = (_00632_ ? _06108_ : _00858_);
	assign _00860_ = _00700_ | _06113_;
	assign _00861_ = _06111_ & ~_00704_;
	assign _00862_ = _00860_ & ~_00861_;
	assign _00863_ = _06462_ & ~_00707_;
	assign _00864_ = _00862_ & ~_00863_;
	assign _00865_ = (_00710_ ? _02616_ : _00864_);
	assign _00867_ = _00297_ ^ _00271_;
	assign _00868_ = _00867_ ^ _00865_;
	assign _00869_ = _00868_ ^ _00859_;
	assign _00870_ = _00869_ ^ _00852_;
	assign _00871_ = _00870_ ^ _00846_;
	assign _00872_ = _00871_ ^ _05911_;
	assign _00873_ = _00465_ | _06134_;
	assign _00874_ = _06131_ & ~_00467_;
	assign _00875_ = _00873_ & ~_00874_;
	assign _00876_ = _06130_ & ~_00471_;
	assign _00878_ = _00875_ & ~_00876_;
	assign _00879_ = (_00474_ ? _06129_ : _00878_);
	assign _00880_ = _00543_ | _06146_;
	assign _00881_ = _06131_ & ~_00545_;
	assign _00882_ = _00880_ & ~_00881_;
	assign _00883_ = _06130_ & ~_00549_;
	assign _00884_ = _00882_ & ~_00883_;
	assign _00885_ = (_00552_ ? _01188_ : _00884_);
	assign _00886_ = _00622_ | _06134_;
	assign _00887_ = _06131_ & ~_00626_;
	assign _00889_ = _00886_ & ~_00887_;
	assign _00890_ = _06130_ & ~_00629_;
	assign _00891_ = _00889_ & ~_00890_;
	assign _00892_ = (_00632_ ? _06160_ : _00891_);
	assign _00893_ = _00700_ | _06163_;
	assign _00894_ = _06162_ & ~_00704_;
	assign _00895_ = _00893_ & ~_00894_;
	assign _00896_ = _06139_ & ~_00707_;
	assign _00897_ = _00895_ & ~_00896_;
	assign _00898_ = (_00710_ ? _01188_ : _00897_);
	assign _00900_ = _00333_ ^ _03700_;
	assign _00901_ = _00900_ ^ _00898_;
	assign _00902_ = _00901_ ^ _00892_;
	assign _00903_ = _00902_ ^ _00885_;
	assign _00904_ = _00903_ ^ _00879_;
	assign _00905_ = _00904_ ^ _06128_;
	assign _00906_ = _00905_ | _00872_;
	assign _00907_ = _00906_ | _03810_;
	assign _00908_ = _00871_ ^ _03744_;
	assign _00909_ = ~(_00908_ & _00905_);
	assign _00911_ = _03239_ & ~_00909_;
	assign _00912_ = _00907_ & ~_00911_;
	assign _00913_ = _00908_ | _00905_;
	assign _00914_ = _03228_ & ~_00913_;
	assign _00915_ = _00912_ & ~_00914_;
	assign _00916_ = _00905_ & ~_00908_;
	assign _00917_ = (_00916_ ? _00996_ : _00915_);
	assign _00918_ = _00465_ | _06192_;
	assign _00919_ = _00344_ & ~_00467_;
	assign _00920_ = _00918_ & ~_00919_;
	assign _00922_ = _03052_ & ~_00471_;
	assign _00923_ = _00920_ & ~_00922_;
	assign _00924_ = (_00474_ ? \mchip.wrapper.keyReg.Q [1] : _00923_);
	assign _00925_ = _00543_ | _06202_;
	assign _00926_ = _00352_ & ~_00545_;
	assign _00927_ = _00925_ & ~_00926_;
	assign _00928_ = _06200_ & ~_00549_;
	assign _00929_ = _00927_ & ~_00928_;
	assign _00930_ = (_00552_ ? _06211_ : _00929_);
	assign _00931_ = _00622_ | _03074_;
	assign _00933_ = _03063_ & ~_00626_;
	assign _00934_ = _00931_ & ~_00933_;
	assign _00935_ = _03052_ & ~_00629_;
	assign _00936_ = _00934_ & ~_00935_;
	assign _00937_ = (_00632_ ? _06220_ : _00936_);
	assign _00938_ = _00700_ | _06223_;
	assign _00939_ = _06222_ & ~_00704_;
	assign _00940_ = _00938_ & ~_00939_;
	assign _00941_ = _06206_ & ~_00707_;
	assign _00942_ = _00940_ & ~_00941_;
	assign _00944_ = (_00710_ ? _06231_ : _00942_);
	assign _00945_ = _00377_ ^ _00344_;
	assign _00946_ = _00945_ ^ _00944_;
	assign _00947_ = _00946_ ^ _00937_;
	assign _00948_ = _00947_ ^ _00930_;
	assign _00949_ = _00948_ ^ _00924_;
	assign _00950_ = _00949_ ^ _06191_;
	assign _00951_ = _00465_ | _06243_;
	assign _00952_ = _06242_ & ~_00467_;
	assign _00953_ = _00951_ & ~_00952_;
	assign _00955_ = _06241_ & ~_00471_;
	assign _00956_ = _00953_ & ~_00955_;
	assign _00957_ = (_00474_ ? \mchip.wrapper.keyReg.Q [0] : _00956_);
	assign _00958_ = _00543_ | _00086_;
	assign _00959_ = _00386_ & ~_00545_;
	assign _00960_ = _00958_ & ~_00959_;
	assign _00961_ = _03952_ & ~_00549_;
	assign _00962_ = _00960_ & ~_00961_;
	assign _00963_ = (_00552_ ? _06259_ : _00962_);
	assign _00964_ = _00622_ | _02279_;
	assign _00966_ = _06263_ & ~_00626_;
	assign _00967_ = _00964_ & ~_00966_;
	assign _00968_ = _06248_ & ~_00629_;
	assign _00969_ = _00967_ & ~_00968_;
	assign _00970_ = (_00632_ ? _06273_ : _00969_);
	assign _00971_ = _00700_ | _06264_;
	assign _00972_ = _06266_ & ~_00704_;
	assign _00973_ = _00971_ & ~_00972_;
	assign _00974_ = _06248_ & ~_00707_;
	assign _00975_ = _00973_ & ~_00974_;
	assign _00977_ = (_00710_ ? _06280_ : _00975_);
	assign _00978_ = _00414_ ^ _03963_;
	assign _00979_ = _00978_ ^ _00977_;
	assign _00980_ = _00979_ ^ _00970_;
	assign _00981_ = _00980_ ^ _00963_;
	assign _00982_ = _00981_ ^ _00957_;
	assign _00983_ = _00982_ ^ _06240_;
	assign _00984_ = _00983_ | _00950_;
	assign _00985_ = _00984_ | _03810_;
	assign _00986_ = _00949_ ^ _03052_;
	assign _00988_ = ~(_00986_ & _00983_);
	assign _00989_ = _03832_ & ~_00988_;
	assign _00990_ = _00985_ & ~_00989_;
	assign _00991_ = _00986_ | _00983_;
	assign _00992_ = _03876_ & ~_00991_;
	assign _00993_ = _00990_ & ~_00992_;
	assign _00994_ = _00983_ & ~_00986_;
	assign _00995_ = (_00994_ ? _04241_ : _00993_);
	assign _00997_ = _00996_ ^ _00431_;
	assign _00999_ = _00997_ ^ _00995_;
	assign _01000_ = _00999_ ^ _00917_;
	assign _01001_ = _01000_ ^ _00839_;
	assign _01002_ = _01001_ ^ _00762_;
	assign _01003_ = _01002_ ^ _03184_;
	assign _01004_ = _00752_ | _03140_;
	assign _01005_ = _03129_ & ~_00754_;
	assign _01006_ = _01004_ & ~_01005_;
	assign _01007_ = _03085_ & ~_00758_;
	assign _01008_ = _01006_ & ~_01007_;
	assign _01010_ = (_00761_ ? _03107_ : _01008_);
	assign _01011_ = _00829_ | _03305_;
	assign _01012_ = _04503_ & ~_00831_;
	assign _01013_ = _01011_ & ~_01012_;
	assign _01014_ = _03283_ & ~_00835_;
	assign _01015_ = _01013_ & ~_01014_;
	assign _01016_ = (_00838_ ? _04471_ : _01015_);
	assign _01017_ = _00906_ | _03305_;
	assign _01018_ = _03294_ & ~_00909_;
	assign _01019_ = _01017_ & ~_01018_;
	assign _01021_ = _03283_ & ~_00913_;
	assign _01022_ = _01019_ & ~_01021_;
	assign _01023_ = (_00916_ ? _04558_ : _01022_);
	assign _01024_ = _00984_ | _01835_;
	assign _01025_ = _03294_ & ~_00988_;
	assign _01026_ = _01024_ & ~_01025_;
	assign _01027_ = _03283_ & ~_00991_;
	assign _01028_ = _01026_ & ~_01027_;
	assign _01029_ = (_00994_ ? _04558_ : _01028_);
	assign _01030_ = _06342_ ^ \mchip.wrapper.keyReg.Q [6];
	assign _01032_ = _01030_ ^ _00464_;
	assign _01033_ = _01032_ ^ _01029_;
	assign _01034_ = _01033_ ^ _01023_;
	assign _01035_ = _01034_ ^ _01016_;
	assign _01036_ = _01035_ ^ _01010_;
	assign _01037_ = _01036_ ^ _06342_;
	assign _01038_ = ~(_01037_ & _01003_);
	assign _01039_ = _01038_ | _03140_;
	assign _01040_ = _01037_ | ~_01003_;
	assign _01041_ = _03129_ & ~_01040_;
	assign _01043_ = _01039_ & ~_01041_;
	assign _01044_ = _01003_ | ~_01037_;
	assign _01045_ = _03085_ & ~_01044_;
	assign _01046_ = _01043_ & ~_01045_;
	assign _01047_ = ~(_01037_ | _01003_);
	assign _01048_ = (_01047_ ? _03107_ : _01046_);
	assign _01049_ = _00752_ | _03481_;
	assign _01050_ = _03470_ & ~_00754_;
	assign _01051_ = _01049_ & ~_01050_;
	assign _01052_ = _03459_ & ~_00758_;
	assign _01054_ = _01051_ & ~_01052_;
	assign _01055_ = (_00761_ ? _04833_ : _01054_);
	assign _01056_ = _00829_ | _04955_;
	assign _01057_ = _06371_ & ~_00831_;
	assign _01058_ = _01056_ & ~_01057_;
	assign _01059_ = _04933_ & ~_00835_;
	assign _01060_ = _01058_ & ~_01059_;
	assign _01061_ = (_00838_ ? _05032_ : _01060_);
	assign _01062_ = _00906_ | _02450_;
	assign _01063_ = _06371_ & ~_00909_;
	assign _01065_ = _01062_ & ~_01063_;
	assign _01066_ = _04933_ & ~_00913_;
	assign _01067_ = _01065_ & ~_01066_;
	assign _01068_ = (_00916_ ? _05129_ : _01067_);
	assign _01069_ = _00984_ | _05152_;
	assign _01070_ = _04855_ & ~_00988_;
	assign _01071_ = _01069_ & ~_01070_;
	assign _01072_ = _03459_ & ~_00991_;
	assign _01073_ = _01071_ & ~_01072_;
	assign _01074_ = (_00994_ ? _01735_ : _01073_);
	assign _01076_ = _06391_ ^ \mchip.wrapper.keyReg.Q [5];
	assign _01077_ = _01076_ ^ _00508_;
	assign _01078_ = _01077_ ^ _01074_;
	assign _01079_ = _01078_ ^ _01068_;
	assign _01080_ = _01079_ ^ _01061_;
	assign _01081_ = _01080_ ^ _01055_;
	assign _01082_ = _01081_ ^ _06391_;
	assign _01083_ = _00752_ | _05348_;
	assign _01084_ = _05337_ & ~_00754_;
	assign _01085_ = _01083_ & ~_01084_;
	assign _01087_ = _05326_ & ~_00758_;
	assign _01088_ = _01085_ & ~_01087_;
	assign _01089_ = (_00761_ ? \mchip.wrapper.keyReg.Q [4] : _01088_);
	assign _01090_ = _00829_ | _03525_;
	assign _01091_ = _00226_ & ~_00831_;
	assign _01092_ = _01090_ & ~_01091_;
	assign _01093_ = _03503_ & ~_00835_;
	assign _01094_ = _01092_ & ~_01093_;
	assign _01095_ = (_00838_ ? _05515_ : _01094_);
	assign _01096_ = _00906_ | _05537_;
	assign _01098_ = _05371_ & ~_00909_;
	assign _01099_ = _01096_ & ~_01098_;
	assign _01100_ = _05326_ & ~_00913_;
	assign _01101_ = _01099_ & ~_01100_;
	assign _01102_ = (_00916_ ? _01110_ : _01101_);
	assign _01103_ = _00984_ | _05646_;
	assign _01104_ = _06415_ & ~_00988_;
	assign _01105_ = _01103_ & ~_01104_;
	assign _01106_ = _05482_ & ~_00991_;
	assign _01107_ = _01105_ & ~_01106_;
	assign _01109_ = (_00994_ ? _05713_ : _01107_);
	assign _01111_ = _01110_ ^ _00542_;
	assign _01112_ = _01111_ ^ _01109_;
	assign _01113_ = _01112_ ^ _01102_;
	assign _01114_ = _01113_ ^ _01095_;
	assign _01115_ = _01114_ ^ _01089_;
	assign _01116_ = _01115_ ^ _03525_;
	assign _01117_ = ~(_01116_ & _01082_);
	assign _01118_ = _01117_ | _03305_;
	assign _01120_ = _01116_ | ~_01082_;
	assign _01121_ = _04503_ & ~_01120_;
	assign _01122_ = _01118_ & ~_01121_;
	assign _01123_ = _01082_ | ~_01116_;
	assign _01124_ = _03283_ & ~_01123_;
	assign _01125_ = _01122_ & ~_01124_;
	assign _01126_ = ~(_01116_ | _01082_);
	assign _01127_ = (_01126_ ? _04471_ : _01125_);
	assign _01128_ = _00752_ | _05945_;
	assign _01129_ = _03755_ & ~_00754_;
	assign _01131_ = _01128_ & ~_01129_;
	assign _01132_ = _03744_ & ~_00758_;
	assign _01133_ = _01131_ & ~_01132_;
	assign _01134_ = (_00761_ ? _03733_ : _01133_);
	assign _01135_ = _00829_ | _05945_;
	assign _01136_ = _00271_ & ~_00831_;
	assign _01137_ = _01135_ & ~_01136_;
	assign _01138_ = _03744_ & ~_00835_;
	assign _01139_ = _01137_ & ~_01138_;
	assign _01140_ = (_00838_ ? _06099_ : _01139_);
	assign _01142_ = _00906_ | _05945_;
	assign _01143_ = _00271_ & ~_00909_;
	assign _01144_ = _01142_ & ~_01143_;
	assign _01145_ = _05911_ & ~_00913_;
	assign _01146_ = _01144_ & ~_01145_;
	assign _01147_ = (_00916_ ? _06108_ : _01146_);
	assign _01148_ = _00984_ | _06113_;
	assign _01149_ = _06111_ & ~_00988_;
	assign _01150_ = _01148_ & ~_01149_;
	assign _01151_ = _06462_ & ~_00991_;
	assign _01153_ = _01150_ & ~_01151_;
	assign _01154_ = (_00994_ ? _02616_ : _01153_);
	assign _01155_ = _00587_ ^ _06099_;
	assign _01156_ = _01155_ ^ _01154_;
	assign _01157_ = _01156_ ^ _01147_;
	assign _01158_ = _01157_ ^ _01140_;
	assign _01159_ = _01158_ ^ _01134_;
	assign _01160_ = _01159_ ^ _05945_;
	assign _01161_ = _00752_ | _06134_;
	assign _01162_ = _06131_ & ~_00754_;
	assign _01164_ = _01161_ & ~_01162_;
	assign _01165_ = _06130_ & ~_00758_;
	assign _01166_ = _01164_ & ~_01165_;
	assign _01167_ = (_00761_ ? _06129_ : _01166_);
	assign _01168_ = _00829_ | _06146_;
	assign _01169_ = _06131_ & ~_00831_;
	assign _01170_ = _01168_ & ~_01169_;
	assign _01171_ = _06130_ & ~_00835_;
	assign _01172_ = _01170_ & ~_01171_;
	assign _01173_ = (_00838_ ? _01188_ : _01172_);
	assign _01175_ = _00906_ | _06134_;
	assign _01176_ = _06131_ & ~_00909_;
	assign _01177_ = _01175_ & ~_01176_;
	assign _01178_ = _06130_ & ~_00913_;
	assign _01179_ = _01177_ & ~_01178_;
	assign _01180_ = (_00916_ ? _06160_ : _01179_);
	assign _01181_ = _00984_ | _06163_;
	assign _01182_ = _06162_ & ~_00988_;
	assign _01183_ = _01181_ & ~_01182_;
	assign _01184_ = _06139_ & ~_00991_;
	assign _01186_ = _01183_ & ~_01184_;
	assign _01187_ = (_00994_ ? _01188_ : _01186_);
	assign _01189_ = ~_01188_;
	assign _01190_ = _00621_ ^ _01189_;
	assign _01191_ = _01190_ ^ _01187_;
	assign _01192_ = _01191_ ^ _01180_;
	assign _01193_ = _01192_ ^ _01173_;
	assign _01194_ = _01193_ ^ _01167_;
	assign _01195_ = _01194_ ^ _06134_;
	assign _01197_ = _01195_ | _01160_;
	assign _01198_ = _01197_ | _03305_;
	assign _01199_ = _01159_ ^ _05934_;
	assign _01200_ = ~(_01199_ & _01195_);
	assign _01201_ = _03294_ & ~_01200_;
	assign _01202_ = _01198_ & ~_01201_;
	assign _01203_ = _01199_ | _01195_;
	assign _01204_ = _03283_ & ~_01203_;
	assign _01205_ = _01202_ & ~_01204_;
	assign _01206_ = _01195_ & ~_01199_;
	assign _01208_ = (_01206_ ? _04558_ : _01205_);
	assign _01209_ = _00752_ | _06192_;
	assign _01210_ = _00344_ & ~_00754_;
	assign _01211_ = _01209_ & ~_01210_;
	assign _01212_ = _03052_ & ~_00758_;
	assign _01213_ = _01211_ & ~_01212_;
	assign _01214_ = (_00761_ ? \mchip.wrapper.keyReg.Q [1] : _01213_);
	assign _01215_ = _00829_ | _06202_;
	assign _01216_ = _00352_ & ~_00831_;
	assign _01217_ = _01215_ & ~_01216_;
	assign _01219_ = _06200_ & ~_00835_;
	assign _01220_ = _01217_ & ~_01219_;
	assign _01221_ = (_00838_ ? _06211_ : _01220_);
	assign _01222_ = _00906_ | _03074_;
	assign _01223_ = _03063_ & ~_00909_;
	assign _01224_ = _01222_ & ~_01223_;
	assign _01225_ = _03052_ & ~_00913_;
	assign _01226_ = _01224_ & ~_01225_;
	assign _01227_ = (_00916_ ? _06220_ : _01226_);
	assign _01228_ = _00984_ | _06223_;
	assign _01230_ = _06222_ & ~_00988_;
	assign _01231_ = _01228_ & ~_01230_;
	assign _01232_ = _06206_ & ~_00991_;
	assign _01233_ = _01231_ & ~_01232_;
	assign _01234_ = (_00994_ ? _06231_ : _01233_);
	assign _01235_ = _00051_ ^ \mchip.wrapper.keyReg.Q [1];
	assign _01236_ = ~_01235_;
	assign _01237_ = _00666_ ^ _01236_;
	assign _01238_ = _01237_ ^ _01234_;
	assign _01239_ = _01238_ ^ _01227_;
	assign _01241_ = _01239_ ^ _01221_;
	assign _01242_ = _01241_ ^ _01214_;
	assign _01243_ = _01242_ ^ _00052_;
	assign _01244_ = _00752_ | _06243_;
	assign _01245_ = _06242_ & ~_00754_;
	assign _01246_ = _01244_ & ~_01245_;
	assign _01247_ = _06241_ & ~_00758_;
	assign _01248_ = _01246_ & ~_01247_;
	assign _01249_ = (_00761_ ? \mchip.wrapper.keyReg.Q [0] : _01248_);
	assign _01250_ = _00829_ | _00086_;
	assign _01252_ = _00386_ & ~_00831_;
	assign _01253_ = _01250_ & ~_01252_;
	assign _01254_ = _03952_ & ~_00835_;
	assign _01255_ = _01253_ & ~_01254_;
	assign _01256_ = (_00838_ ? _06259_ : _01255_);
	assign _01257_ = _00906_ | _02279_;
	assign _01258_ = _06263_ & ~_00909_;
	assign _01259_ = _01257_ & ~_01258_;
	assign _01260_ = _06248_ & ~_00913_;
	assign _01261_ = _01259_ & ~_01260_;
	assign _01263_ = (_00916_ ? _06273_ : _01261_);
	assign _01264_ = _00984_ | _06264_;
	assign _01265_ = _06266_ & ~_00988_;
	assign _01266_ = _01264_ & ~_01265_;
	assign _01267_ = _06248_ & ~_00991_;
	assign _01268_ = _01266_ & ~_01267_;
	assign _01269_ = (_00994_ ? _06280_ : _01268_);
	assign _01270_ = _00086_ ^ _06262_;
	assign _01271_ = ~_01270_;
	assign _01272_ = _00699_ ^ _01271_;
	assign _01274_ = _01272_ ^ _01269_;
	assign _01275_ = _01274_ ^ _01263_;
	assign _01276_ = _01275_ ^ _01256_;
	assign _01277_ = _01276_ ^ _01249_;
	assign _01278_ = _01277_ ^ _00088_;
	assign _01279_ = _01278_ | _01243_;
	assign _01280_ = _01279_ | _01835_;
	assign _01281_ = _01242_ ^ _00051_;
	assign _01282_ = ~(_01281_ & _01278_);
	assign _01283_ = _03294_ & ~_01282_;
	assign _01285_ = _01280_ & ~_01283_;
	assign _01286_ = _01281_ | _01278_;
	assign _01287_ = _03283_ & ~_01286_;
	assign _01288_ = _01285_ & ~_01287_;
	assign _01289_ = _01278_ & ~_01281_;
	assign _01290_ = (_01289_ ? _04558_ : _01288_);
	assign _01291_ = _00751_ ^ _06341_;
	assign _01292_ = _01291_ ^ _01290_;
	assign _01293_ = _01292_ ^ _01208_;
	assign _01294_ = _01293_ ^ _01127_;
	assign _01296_ = _01294_ ^ _01048_;
	assign _01297_ = _01296_ ^ _03096_;
	assign _01298_ = _01038_ | _03217_;
	assign _01299_ = _03206_ & ~_01040_;
	assign _01300_ = _01298_ & ~_01299_;
	assign _01301_ = _03162_ & ~_01044_;
	assign _01302_ = _01300_ & ~_01301_;
	assign _01303_ = (_01047_ ? _03195_ : _01302_);
	assign _01304_ = _01117_ | _03184_;
	assign _01305_ = _03173_ & ~_01120_;
	assign _01307_ = _01304_ & ~_01305_;
	assign _01308_ = _03162_ & ~_01123_;
	assign _01309_ = _01307_ & ~_01308_;
	assign _01310_ = (_01126_ ? _03667_ : _01309_);
	assign _01311_ = _01197_ | _03810_;
	assign _01312_ = _03239_ & ~_01200_;
	assign _01313_ = _01311_ & ~_01312_;
	assign _01314_ = _03228_ & ~_01203_;
	assign _01315_ = _01313_ & ~_01314_;
	assign _01316_ = (_01206_ ? _00996_ : _01315_);
	assign _01318_ = _01279_ | _03810_;
	assign _01319_ = _03832_ & ~_01282_;
	assign _01320_ = _01318_ & ~_01319_;
	assign _01321_ = _03876_ & ~_01286_;
	assign _01322_ = _01320_ & ~_01321_;
	assign _01323_ = (_01289_ ? _04241_ : _01322_);
	assign _01324_ = _00718_ ^ _03173_;
	assign _01325_ = _01324_ ^ _01323_;
	assign _01326_ = _01325_ ^ _01316_;
	assign _01327_ = _01326_ ^ _01310_;
	assign _01329_ = _01327_ ^ _01303_;
	assign _01330_ = _01329_ ^ _03162_;
	assign _01331_ = _01297_ | ~_01330_;
	assign _01332_ = _01331_ | ~_03074_;
	assign _01333_ = ~(_01330_ & _01297_);
	assign _01334_ = _00344_ & ~_01333_;
	assign _01335_ = _01332_ & ~_01334_;
	assign _01336_ = _01330_ | _01297_;
	assign _01337_ = _03052_ & ~_01336_;
	assign _01338_ = _01337_ | ~_01335_;
	assign _01340_ = _01297_ & ~_01330_;
	assign _01341_ = (_01340_ ? _03041_ : _01338_);
	assign _01342_ = _01038_ | _05348_;
	assign _01343_ = _05337_ & ~_01040_;
	assign _01344_ = _01342_ & ~_01343_;
	assign _01345_ = _05326_ & ~_01044_;
	assign _01346_ = _01344_ & ~_01345_;
	assign _01347_ = (_01047_ ? \mchip.wrapper.keyReg.Q [4] : _01346_);
	assign _01348_ = _01117_ | _03525_;
	assign _01349_ = _00226_ & ~_01120_;
	assign _01351_ = _01348_ & ~_01349_;
	assign _01352_ = _03503_ & ~_01123_;
	assign _01353_ = _01351_ & ~_01352_;
	assign _01354_ = (_01126_ ? _05515_ : _01353_);
	assign _01355_ = _01197_ | _05537_;
	assign _01356_ = _05371_ & ~_01200_;
	assign _01357_ = _01355_ & ~_01356_;
	assign _01358_ = _05326_ & ~_01203_;
	assign _01359_ = _01357_ & ~_01358_;
	assign _01360_ = (_01206_ ? _01110_ : _01359_);
	assign _01362_ = _01279_ | _05646_;
	assign _01363_ = _06415_ & ~_01282_;
	assign _01364_ = _01362_ & ~_01363_;
	assign _01365_ = _05482_ & ~_01286_;
	assign _01366_ = _01364_ & ~_01365_;
	assign _01367_ = (_01289_ ? _05713_ : _01366_);
	assign _01368_ = _00828_ ^ _03514_;
	assign _01369_ = _01368_ ^ _01367_;
	assign _01370_ = _01369_ ^ _01360_;
	assign _01371_ = _01370_ ^ _01354_;
	assign _01373_ = _01371_ ^ _01347_;
	assign _01374_ = _01373_ ^ _03503_;
	assign _01375_ = _01038_ | _03481_;
	assign _01376_ = _03470_ & ~_01040_;
	assign _01377_ = _01375_ & ~_01376_;
	assign _01378_ = _03459_ & ~_01044_;
	assign _01379_ = _01377_ & ~_01378_;
	assign _01380_ = (_01047_ ? _04833_ : _01379_);
	assign _01381_ = _01117_ | _04955_;
	assign _01382_ = _06371_ & ~_01120_;
	assign _01384_ = _01381_ & ~_01382_;
	assign _01385_ = _04933_ & ~_01123_;
	assign _01386_ = _01384_ & ~_01385_;
	assign _01387_ = (_01126_ ? _05032_ : _01386_);
	assign _01388_ = _01197_ | _02450_;
	assign _01389_ = _06371_ & ~_01200_;
	assign _01390_ = _01388_ & ~_01389_;
	assign _01391_ = _04933_ & ~_01203_;
	assign _01392_ = _01390_ & ~_01391_;
	assign _01393_ = (_01206_ ? _05129_ : _01392_);
	assign _01395_ = _01279_ | _05152_;
	assign _01396_ = _04855_ & ~_01282_;
	assign _01397_ = _01395_ & ~_01396_;
	assign _01398_ = _03459_ & ~_01286_;
	assign _01399_ = _01397_ & ~_01398_;
	assign _01400_ = (_01289_ ? _01735_ : _01399_);
	assign _01401_ = _00795_ ^ _06389_;
	assign _01402_ = _01401_ ^ _01400_;
	assign _01403_ = _01402_ ^ _01393_;
	assign _01404_ = _01403_ ^ _01387_;
	assign _01406_ = _01404_ ^ _01380_;
	assign _01407_ = _01406_ ^ _04888_;
	assign _01408_ = _01407_ | ~_01374_;
	assign _01409_ = ~(_01408_ | _06202_);
	assign _01410_ = _01407_ | _01374_;
	assign _01411_ = _00352_ & ~_01410_;
	assign _01412_ = _01411_ | _01409_;
	assign _01413_ = ~(_01407_ & _01374_);
	assign _01414_ = _06200_ & ~_01413_;
	assign _01415_ = _01414_ | _01412_;
	assign _01417_ = _01407_ & ~_01374_;
	assign _01418_ = (_01417_ ? _06210_ : _01415_);
	assign _01419_ = _01038_ | _06134_;
	assign _01420_ = _06131_ & ~_01040_;
	assign _01421_ = _01419_ & ~_01420_;
	assign _01422_ = _06130_ & ~_01044_;
	assign _01423_ = _01421_ & ~_01422_;
	assign _01424_ = (_01047_ ? _06129_ : _01423_);
	assign _01425_ = _01117_ | _06146_;
	assign _01426_ = _06131_ & ~_01120_;
	assign _01428_ = _01425_ & ~_01426_;
	assign _01429_ = _06130_ & ~_01123_;
	assign _01430_ = _01428_ & ~_01429_;
	assign _01431_ = (_01126_ ? _01188_ : _01430_);
	assign _01432_ = _01197_ | _06134_;
	assign _01433_ = _06131_ & ~_01200_;
	assign _01434_ = _01432_ & ~_01433_;
	assign _01435_ = _06130_ & ~_01203_;
	assign _01436_ = _01434_ & ~_01435_;
	assign _01437_ = (_01206_ ? _06160_ : _01436_);
	assign _01439_ = _01279_ | _06163_;
	assign _01440_ = _06162_ & ~_01282_;
	assign _01441_ = _01439_ & ~_01440_;
	assign _01442_ = _06139_ & ~_01286_;
	assign _01443_ = _01441_ & ~_01442_;
	assign _01444_ = (_01289_ ? _01188_ : _01443_);
	assign _01445_ = _00905_ ^ _06136_;
	assign _01446_ = _01445_ ^ _01444_;
	assign _01447_ = _01446_ ^ _01437_;
	assign _01448_ = _01447_ ^ _01431_;
	assign _01450_ = _01448_ ^ _01424_;
	assign _01451_ = _01450_ ^ _06139_;
	assign _01452_ = _01038_ | _05945_;
	assign _01453_ = _03755_ & ~_01040_;
	assign _01454_ = _01452_ & ~_01453_;
	assign _01455_ = _03744_ & ~_01044_;
	assign _01456_ = _01454_ & ~_01455_;
	assign _01457_ = (_01047_ ? _03733_ : _01456_);
	assign _01458_ = _01117_ | _05945_;
	assign _01459_ = _00271_ & ~_01120_;
	assign _01461_ = _01458_ & ~_01459_;
	assign _01462_ = _03744_ & ~_01123_;
	assign _01463_ = _01461_ & ~_01462_;
	assign _01464_ = (_01126_ ? _06099_ : _01463_);
	assign _01465_ = _01197_ | _05945_;
	assign _01466_ = _00271_ & ~_01200_;
	assign _01467_ = _01465_ & ~_01466_;
	assign _01468_ = _05911_ & ~_01203_;
	assign _01469_ = _01467_ & ~_01468_;
	assign _01470_ = (_01206_ ? _06108_ : _01469_);
	assign _01472_ = _01279_ | _06113_;
	assign _01473_ = _06111_ & ~_01282_;
	assign _01474_ = _01472_ & ~_01473_;
	assign _01475_ = _06462_ & ~_01286_;
	assign _01476_ = _01474_ & ~_01475_;
	assign _01477_ = (_01289_ ? _02616_ : _01476_);
	assign _01478_ = _00872_ ^ _00271_;
	assign _01479_ = _01478_ ^ _01477_;
	assign _01480_ = _01479_ ^ _01470_;
	assign _01481_ = _01480_ ^ _01464_;
	assign _01483_ = _01481_ ^ _01457_;
	assign _01484_ = _01483_ ^ _05911_;
	assign _01485_ = _01484_ | _01451_;
	assign _01486_ = _00051_ & ~_01485_;
	assign _01487_ = _01484_ | ~_01451_;
	assign _01488_ = _03063_ & ~_01487_;
	assign _01489_ = _01488_ | _01486_;
	assign _01490_ = _01451_ | ~_01484_;
	assign _01491_ = _03052_ & ~_01490_;
	assign _01492_ = _01491_ | _01489_;
	assign _01494_ = _01484_ & _01451_;
	assign _01495_ = (_01494_ ? _06219_ : _01492_);
	assign _01496_ = _01038_ | _06192_;
	assign _01497_ = _00344_ & ~_01040_;
	assign _01498_ = _01496_ & ~_01497_;
	assign _01499_ = _03052_ & ~_01044_;
	assign _01500_ = _01498_ & ~_01499_;
	assign _01501_ = (_01047_ ? \mchip.wrapper.keyReg.Q [1] : _01500_);
	assign _01502_ = _01117_ | _06202_;
	assign _01503_ = _00352_ & ~_01120_;
	assign _01505_ = _01502_ & ~_01503_;
	assign _01506_ = _06200_ & ~_01123_;
	assign _01507_ = _01505_ & ~_01506_;
	assign _01508_ = (_01126_ ? _06211_ : _01507_);
	assign _01509_ = _01197_ | _03074_;
	assign _01510_ = _03063_ & ~_01200_;
	assign _01511_ = _01509_ & ~_01510_;
	assign _01512_ = _03052_ & ~_01203_;
	assign _01513_ = _01511_ & ~_01512_;
	assign _01514_ = (_01206_ ? _06220_ : _01513_);
	assign _01516_ = _01279_ | _06223_;
	assign _01517_ = _06222_ & ~_01282_;
	assign _01518_ = _01516_ & ~_01517_;
	assign _01519_ = _06206_ & ~_01286_;
	assign _01520_ = _01518_ & ~_01519_;
	assign _01521_ = (_01289_ ? _06231_ : _01520_);
	assign _01522_ = _00950_ ^ _03063_;
	assign _01523_ = _01522_ ^ _01521_;
	assign _01524_ = _01523_ ^ _01514_;
	assign _01525_ = _01524_ ^ _01508_;
	assign _01527_ = _01525_ ^ _01501_;
	assign _01528_ = _01527_ ^ _06191_;
	assign _01529_ = _01038_ | _06243_;
	assign _01530_ = _06242_ & ~_01040_;
	assign _01531_ = _01529_ & ~_01530_;
	assign _01532_ = _06241_ & ~_01044_;
	assign _01533_ = _01531_ & ~_01532_;
	assign _01534_ = (_01047_ ? \mchip.wrapper.keyReg.Q [0] : _01533_);
	assign _01535_ = _01117_ | _00086_;
	assign _01536_ = _00386_ & ~_01120_;
	assign _01538_ = _01535_ & ~_01536_;
	assign _01539_ = _03952_ & ~_01123_;
	assign _01540_ = _01538_ & ~_01539_;
	assign _01541_ = (_01126_ ? _06259_ : _01540_);
	assign _01542_ = _01197_ | _02279_;
	assign _01543_ = _06263_ & ~_01200_;
	assign _01544_ = _01542_ & ~_01543_;
	assign _01545_ = _06248_ & ~_01203_;
	assign _01546_ = _01544_ & ~_01545_;
	assign _01547_ = (_01206_ ? _06273_ : _01546_);
	assign _01549_ = _01279_ | _06264_;
	assign _01550_ = _06266_ & ~_01282_;
	assign _01551_ = _01549_ & ~_01550_;
	assign _01552_ = _06248_ & ~_01286_;
	assign _01553_ = _01551_ & ~_01552_;
	assign _01554_ = (_01289_ ? _06280_ : _01553_);
	assign _01555_ = _00983_ ^ _00386_;
	assign _01556_ = _01555_ ^ _01554_;
	assign _01557_ = _01556_ ^ _01547_;
	assign _01558_ = _01557_ ^ _01541_;
	assign _01560_ = _01558_ ^ _01534_;
	assign _01561_ = _01560_ ^ _06240_;
	assign _01562_ = _01561_ | _01528_;
	assign _01563_ = _01562_ | _06223_;
	assign _01564_ = _01560_ ^ _03952_;
	assign _01565_ = _01564_ | _01528_;
	assign _01566_ = _06222_ & ~_01565_;
	assign _01567_ = _01563_ & ~_01566_;
	assign _01568_ = ~(_01564_ & _01528_);
	assign _01569_ = ~(_01568_ | _06200_);
	assign _01571_ = _01567_ & ~_01569_;
	assign _01572_ = _01528_ & ~_01564_;
	assign _01573_ = (_01572_ ? _06231_ : _01571_);
	assign _01574_ = _01243_ ^ _03041_;
	assign _01575_ = _01574_ ^ _01573_;
	assign _01576_ = _01575_ ^ _01495_;
	assign _01577_ = _01576_ ^ _01418_;
	assign _01578_ = ~(_01577_ ^ _01341_);
	assign _01579_ = _01331_ | ~_00089_;
	assign _01580_ = _06242_ & ~_01333_;
	assign _01582_ = _01579_ & ~_01580_;
	assign _01583_ = ~(_01336_ | _06248_);
	assign _01584_ = _01583_ | ~_01582_;
	assign _01585_ = (_01340_ ? _06262_ : _01584_);
	assign _01586_ = ~(_01408_ | _00086_);
	assign _01587_ = _00386_ & ~_01410_;
	assign _01588_ = _01587_ | _01586_;
	assign _01589_ = _03952_ & ~_01413_;
	assign _01590_ = _01589_ | _01588_;
	assign _01591_ = (_01417_ ? _06258_ : _01590_);
	assign _01593_ = _06264_ & ~_01485_;
	assign _01594_ = _06263_ & ~_01487_;
	assign _01595_ = _01594_ | _01593_;
	assign _01596_ = _06248_ & ~_01490_;
	assign _01597_ = _01596_ | _01595_;
	assign _01598_ = (_01494_ ? _06272_ : _01597_);
	assign _01599_ = _01562_ | _06264_;
	assign _01600_ = ~(_01565_ | _06263_);
	assign _01601_ = _01599_ & ~_01600_;
	assign _01602_ = _06248_ & ~_01568_;
	assign _01604_ = _01601_ & ~_01602_;
	assign _01605_ = (_01572_ ? _06280_ : _01604_);
	assign _01606_ = _01278_ ^ _06262_;
	assign _01607_ = _01606_ ^ _01605_;
	assign _01608_ = _01607_ ^ _01598_;
	assign _01609_ = _01608_ ^ _01591_;
	assign _01610_ = _01609_ ^ _01585_;
	assign _01611_ = _01578_ & ~_01610_;
	assign _01612_ = ~(_01331_ | _05945_);
	assign _01613_ = _03755_ & ~_01333_;
	assign _01615_ = _01613_ | _01612_;
	assign _01616_ = _03744_ & ~_01336_;
	assign _01617_ = _01616_ | _01615_;
	assign _01618_ = (_01340_ ? \mchip.wrapper.keyReg.Q [3] : _01617_);
	assign _01619_ = _01408_ | _05945_;
	assign _01620_ = _00271_ & ~_01410_;
	assign _01621_ = _01619_ & ~_01620_;
	assign _01622_ = _03744_ & ~_01413_;
	assign _01623_ = _01621_ & ~_01622_;
	assign _01624_ = (_01417_ ? _06099_ : _01623_);
	assign _01626_ = _01485_ | _05945_;
	assign _01627_ = _00271_ & ~_01487_;
	assign _01628_ = _01626_ & ~_01627_;
	assign _01629_ = _05911_ & ~_01490_;
	assign _01630_ = _01628_ & ~_01629_;
	assign _01631_ = (_01494_ ? _06108_ : _01630_);
	assign _01632_ = ~(_01562_ | _06113_);
	assign _01633_ = _06111_ & ~_01565_;
	assign _01634_ = _01633_ | _01632_;
	assign _01635_ = _06462_ & ~_01568_;
	assign _01637_ = _01635_ | _01634_;
	assign _01638_ = (_01572_ ? _06099_ : _01637_);
	assign _01639_ = _01160_ ^ _03733_;
	assign _01640_ = _01639_ ^ _01638_;
	assign _01641_ = _01640_ ^ _01631_;
	assign _01642_ = _01641_ ^ _01624_;
	assign _01643_ = _01642_ ^ _01618_;
	assign _01644_ = _01331_ | _06134_;
	assign _01645_ = _06131_ & ~_01333_;
	assign _01646_ = _01644_ & ~_01645_;
	assign _01648_ = _06130_ & ~_01336_;
	assign _01649_ = _01646_ & ~_01648_;
	assign _01650_ = (_01340_ ? _06129_ : _01649_);
	assign _01651_ = ~(_01408_ | _06146_);
	assign _01652_ = _06131_ & ~_01410_;
	assign _01653_ = _01652_ | _01651_;
	assign _01654_ = _06130_ & ~_01413_;
	assign _01655_ = _01654_ | _01653_;
	assign _01656_ = (_01417_ ? _01189_ : _01655_);
	assign _01658_ = _06133_ & ~_01485_;
	assign _01659_ = _06131_ & ~_01487_;
	assign _01660_ = _01659_ | _01658_;
	assign _01661_ = _06130_ & ~_01490_;
	assign _01662_ = _01661_ | _01660_;
	assign _01663_ = (_01494_ ? _06159_ : _01662_);
	assign _01664_ = _01562_ | _06163_;
	assign _01665_ = _06162_ & ~_01565_;
	assign _01666_ = _01664_ & ~_01665_;
	assign _01667_ = ~(_01568_ | _06130_);
	assign _01669_ = _01666_ & ~_01667_;
	assign _01670_ = (_01572_ ? _01188_ : _01669_);
	assign _01671_ = _01195_ ^ \mchip.wrapper.keyReg.Q [2];
	assign _01672_ = _01671_ ^ _01670_;
	assign _01673_ = _01672_ ^ _01663_;
	assign _01674_ = _01673_ ^ _01656_;
	assign _01675_ = _01674_ ^ _01650_;
	assign _01676_ = ~(_01675_ & _01643_);
	assign _01677_ = _01611_ & ~_01676_;
	assign _01678_ = ~(_01610_ & _01578_);
	assign _01680_ = ~(_01678_ | _01676_);
	assign _01681_ = _01610_ | _01578_;
	assign _01682_ = _01681_ | _01676_;
	assign _01683_ = _01643_ | ~_01675_;
	assign _01684_ = _01683_ | ~_01611_;
	assign _01685_ = ~(_01683_ | _01681_);
	assign _01686_ = _01675_ | _01643_;
	assign _01687_ = _01578_ | ~_01610_;
	assign _01688_ = ~(_01687_ | _01686_);
	assign _01689_ = ~(_01686_ | _01681_);
	assign _01691_ = _01689_ | ~_01688_;
	assign _01692_ = ~(_01686_ | _01678_);
	assign _01693_ = _01691_ & ~_01692_;
	assign _01694_ = _01611_ & ~_01686_;
	assign _01695_ = _01694_ | ~_01693_;
	assign _01696_ = ~(_01687_ | _01683_);
	assign _01697_ = _01695_ & ~_01696_;
	assign _01698_ = _01697_ | _01685_;
	assign _01699_ = _01683_ | _01678_;
	assign _01700_ = _01699_ & ~_01698_;
	assign _01702_ = _01700_ & _01684_;
	assign _01703_ = _01675_ | ~_01643_;
	assign _01704_ = ~(_01703_ | _01687_);
	assign _01705_ = _01702_ & ~_01704_;
	assign _01706_ = ~(_01703_ | _01681_);
	assign _01707_ = _01705_ & ~_01706_;
	assign _01708_ = ~(_01703_ | _01678_);
	assign _01709_ = _01707_ & ~_01708_;
	assign _01710_ = _01611_ & ~_01703_;
	assign _01711_ = _01710_ | _01709_;
	assign _01713_ = _01687_ | _01676_;
	assign _01714_ = _01713_ & _01711_;
	assign _01715_ = _01682_ & ~_01714_;
	assign _01716_ = _01715_ | _01680_;
	assign _01717_ = _01716_ | _01677_;
	assign _01718_ = _03030_ & ~_01717_;
	assign _01719_ = _04591_ & ~_03019_;
	assign _01720_ = _01331_ | ~_06355_;
	assign _01721_ = _03470_ & ~_01333_;
	assign _01722_ = _01720_ & ~_01721_;
	assign _01724_ = _03459_ & ~_01336_;
	assign _01725_ = _01724_ | ~_01722_;
	assign _01726_ = (_01340_ ? \mchip.wrapper.keyReg.Q [5] : _01725_);
	assign _01727_ = ~_05032_;
	assign _01728_ = ~(_01408_ | _04955_);
	assign _01729_ = _06371_ & ~_01410_;
	assign _01730_ = _01729_ | _01728_;
	assign _01731_ = _04933_ & ~_01413_;
	assign _01732_ = _01731_ | _01730_;
	assign _01733_ = (_01417_ ? _01727_ : _01732_);
	assign _01736_ = _04955_ & ~_01485_;
	assign _01737_ = _06371_ & ~_01487_;
	assign _01738_ = _01737_ | _01736_;
	assign _01739_ = _04933_ & ~_01490_;
	assign _01740_ = _01739_ | _01738_;
	assign _01741_ = (_01494_ ? _01735_ : _01740_);
	assign _01742_ = _01562_ | _05152_;
	assign _01743_ = ~(_01565_ | _03470_);
	assign _01744_ = _01742_ & ~_01743_;
	assign _01746_ = _03459_ & ~_01568_;
	assign _01747_ = _01744_ & ~_01746_;
	assign _01748_ = (_01572_ ? _01735_ : _01747_);
	assign _01749_ = _01082_ ^ _04833_;
	assign _01750_ = _01749_ ^ _01748_;
	assign _01751_ = _01750_ ^ _01741_;
	assign _01752_ = _01751_ ^ _01733_;
	assign _01753_ = ~(_01752_ ^ _01726_);
	assign _01754_ = _01331_ | _05348_;
	assign _01755_ = _05337_ & ~_01333_;
	assign _01757_ = _01754_ & ~_01755_;
	assign _01758_ = _05326_ & ~_01336_;
	assign _01759_ = _01758_ | ~_01757_;
	assign _01760_ = (_01340_ ? _05624_ : _01759_);
	assign _01761_ = ~(_01408_ | _03525_);
	assign _01762_ = _00226_ & ~_01410_;
	assign _01763_ = _01762_ | _01761_;
	assign _01764_ = _03503_ & ~_01413_;
	assign _01765_ = ~(_01764_ | _01763_);
	assign _01766_ = (_01417_ ? _05515_ : _01765_);
	assign _01768_ = ~(_01485_ | _05537_);
	assign _01769_ = _05371_ & ~_01487_;
	assign _01770_ = _01769_ | _01768_;
	assign _01771_ = _05326_ & ~_01490_;
	assign _01772_ = ~(_01771_ | _01770_);
	assign _01773_ = (_01494_ ? _01110_ : _01772_);
	assign _01774_ = _01562_ | _05646_;
	assign _01775_ = _06415_ & ~_01565_;
	assign _01776_ = _01774_ & ~_01775_;
	assign _01777_ = ~(_01568_ | _03503_);
	assign _01779_ = _01776_ & ~_01777_;
	assign _01780_ = (_01572_ ? _05713_ : _01779_);
	assign _01781_ = _01116_ ^ \mchip.wrapper.keyReg.Q [4];
	assign _01782_ = ~(_01781_ ^ _01780_);
	assign _01783_ = _01782_ ^ _01773_;
	assign _01784_ = ~(_01783_ ^ _01766_);
	assign _01785_ = _01784_ ^ _01760_;
	assign _01786_ = _01753_ & ~_01785_;
	assign _01787_ = _03261_ & ~_01331_;
	assign _01788_ = _03206_ & ~_01333_;
	assign _01790_ = _01788_ | _01787_;
	assign _01791_ = _03162_ & ~_01336_;
	assign _01792_ = _01791_ | _01790_;
	assign _01793_ = (_01340_ ? \mchip.wrapper.keyReg.Q [7] : _01792_);
	assign _01794_ = _01408_ | _03184_;
	assign _01795_ = _03173_ & ~_01410_;
	assign _01796_ = _01794_ & ~_01795_;
	assign _01797_ = _03162_ & ~_01413_;
	assign _01798_ = _01796_ & ~_01797_;
	assign _01799_ = (_01417_ ? _03667_ : _01798_);
	assign _01801_ = _01485_ | _03810_;
	assign _01802_ = _03239_ & ~_01487_;
	assign _01803_ = _01801_ & ~_01802_;
	assign _01804_ = _03228_ & ~_01490_;
	assign _01805_ = _01803_ & ~_01804_;
	assign _01806_ = (_01494_ ? _00996_ : _01805_);
	assign _01807_ = ~(_01562_ | _03810_);
	assign _01808_ = _03832_ & ~_01565_;
	assign _01809_ = _01808_ | _01807_;
	assign _01810_ = ~(_01568_ | _03228_);
	assign _01812_ = _01810_ | _01809_;
	assign _01813_ = (_01572_ ? _04230_ : _01812_);
	assign _01814_ = _01003_ ^ \mchip.wrapper.keyReg.Q [7];
	assign _01815_ = _01814_ ^ _01813_;
	assign _01816_ = _01815_ ^ _01806_;
	assign _01817_ = _01816_ ^ _01799_;
	assign _01818_ = _01817_ ^ _01793_;
	assign _01819_ = _01331_ | ~_06308_;
	assign _01820_ = _03129_ & ~_01333_;
	assign _01821_ = _01819_ & ~_01820_;
	assign _01823_ = _03085_ & ~_01336_;
	assign _01824_ = _01821_ & ~_01823_;
	assign _01825_ = (_01340_ ? _03107_ : _01824_);
	assign _01826_ = ~_04471_;
	assign _01827_ = ~(_01408_ | _03305_);
	assign _01828_ = ~(_01410_ | _03294_);
	assign _01829_ = _01828_ | _01827_;
	assign _01830_ = _03283_ & ~_01413_;
	assign _01831_ = _01830_ | _01829_;
	assign _01832_ = (_01417_ ? _01826_ : _01831_);
	assign _01834_ = ~_04558_;
	assign _01836_ = _01835_ & ~_01485_;
	assign _01837_ = _03294_ & ~_01487_;
	assign _01838_ = _01837_ | _01836_;
	assign _01839_ = _03283_ & ~_01490_;
	assign _01840_ = _01839_ | _01838_;
	assign _01841_ = (_01494_ ? _01834_ : _01840_);
	assign _01842_ = _01562_ | _01835_;
	assign _01843_ = _03294_ & ~_01565_;
	assign _01845_ = _01842_ & ~_01843_;
	assign _01846_ = _03283_ & ~_01568_;
	assign _01847_ = _01845_ & ~_01846_;
	assign _01848_ = (_01572_ ? _04558_ : _01847_);
	assign _01849_ = _01037_ ^ \mchip.wrapper.keyReg.Q [6];
	assign _01850_ = _01849_ ^ _01848_;
	assign _01851_ = _01850_ ^ _01841_;
	assign _01852_ = _01851_ ^ _01832_;
	assign _01853_ = _01852_ ^ _01825_;
	assign _01854_ = ~(_01853_ & _01818_);
	assign _01856_ = _01786_ & ~_01854_;
	assign _01857_ = ~(_01785_ & _01753_);
	assign _01858_ = ~(_01857_ | _01854_);
	assign _01859_ = _01785_ | _01753_;
	assign _01860_ = _01859_ | _01854_;
	assign _01861_ = _01818_ | ~_01853_;
	assign _01862_ = _01861_ | ~_01786_;
	assign _01863_ = ~(_01861_ | _01859_);
	assign _01864_ = _01853_ | _01818_;
	assign _01865_ = _01753_ | ~_01785_;
	assign _01867_ = ~(_01865_ | _01864_);
	assign _01868_ = ~(_01864_ | _01859_);
	assign _01869_ = _01868_ | ~_01867_;
	assign _01870_ = ~(_01864_ | _01857_);
	assign _01871_ = _01869_ & ~_01870_;
	assign _01872_ = _01786_ & ~_01864_;
	assign _01873_ = _01872_ | ~_01871_;
	assign _01874_ = ~(_01865_ | _01861_);
	assign _01875_ = _01873_ & ~_01874_;
	assign _01876_ = _01875_ | _01863_;
	assign _01878_ = _01861_ | _01857_;
	assign _01879_ = _01878_ & ~_01876_;
	assign _01880_ = _01879_ & _01862_;
	assign _01881_ = _01853_ | ~_01818_;
	assign _01882_ = ~(_01881_ | _01865_);
	assign _01883_ = _01880_ & ~_01882_;
	assign _01884_ = ~(_01881_ | _01859_);
	assign _01885_ = _01883_ & ~_01884_;
	assign _01886_ = ~(_01881_ | _01857_);
	assign _01887_ = _01885_ & ~_01886_;
	assign _01889_ = _01786_ & ~_01881_;
	assign _01890_ = _01889_ | _01887_;
	assign _01891_ = _01865_ | _01854_;
	assign _01892_ = _01891_ & _01890_;
	assign _01893_ = _01860_ & ~_01892_;
	assign _01894_ = _01893_ | _01858_;
	assign _01895_ = _01894_ | _01856_;
	assign _01896_ = _01719_ & ~_01895_;
	assign _01897_ = _01896_ | _01718_;
	assign _01898_ = _06444_ & ~_03019_;
	assign _01900_ = ~(_01562_ | _01485_);
	assign _01901_ = ~(_01565_ | _01485_);
	assign _01902_ = ~(_01568_ | _01485_);
	assign _01903_ = ~_01902_;
	assign _01904_ = _01565_ | _01490_;
	assign _01905_ = ~(_01568_ | _01490_);
	assign _01906_ = _01494_ & ~_01568_;
	assign _01907_ = ~(_01561_ & _01528_);
	assign _01908_ = _01494_ & ~_01907_;
	assign _01909_ = _01906_ | ~_01908_;
	assign _01911_ = _01494_ & ~_01565_;
	assign _01912_ = _01909_ & ~_01911_;
	assign _01913_ = _01494_ & ~_01562_;
	assign _01914_ = _01913_ | ~_01912_;
	assign _01915_ = ~(_01907_ | _01490_);
	assign _01916_ = _01914_ & ~_01915_;
	assign _01917_ = _01916_ | _01905_;
	assign _01918_ = _01904_ & ~_01917_;
	assign _01919_ = ~(_01562_ | _01490_);
	assign _01920_ = _01918_ & ~_01919_;
	assign _01922_ = ~(_01907_ | _01487_);
	assign _01923_ = _01920_ & ~_01922_;
	assign _01924_ = ~(_01568_ | _01487_);
	assign _01925_ = _01923_ & ~_01924_;
	assign _01926_ = ~(_01565_ | _01487_);
	assign _01927_ = _01925_ & ~_01926_;
	assign _01928_ = ~(_01562_ | _01487_);
	assign _01929_ = _01928_ | _01927_;
	assign _01930_ = ~(_01907_ | _01485_);
	assign _01931_ = ~_01930_;
	assign _01933_ = _01931_ & _01929_;
	assign _01934_ = _01903_ & ~_01933_;
	assign _01935_ = _01934_ | _01901_;
	assign _01936_ = _01935_ | _01900_;
	assign _01937_ = _01898_ & ~_01936_;
	assign _01938_ = _00492_ & ~_03019_;
	assign _01939_ = ~(_01408_ | _01331_);
	assign _01940_ = ~(_01410_ | _01331_);
	assign _01941_ = ~(_01413_ | _01331_);
	assign _01942_ = ~_01941_;
	assign _01944_ = ~(_01410_ | _01336_);
	assign _01945_ = ~_01944_;
	assign _01946_ = ~(_01413_ | _01336_);
	assign _01947_ = _01340_ & ~_01374_;
	assign _01948_ = _01340_ & ~_01408_;
	assign _01949_ = _01948_ | _01947_;
	assign _01950_ = _01417_ & ~_01336_;
	assign _01951_ = _01949_ & ~_01950_;
	assign _01952_ = _01951_ | _01946_;
	assign _01953_ = _01945_ & ~_01952_;
	assign _01955_ = ~(_01408_ | _01336_);
	assign _01956_ = _01953_ & ~_01955_;
	assign _01957_ = _01417_ & ~_01333_;
	assign _01958_ = _01956_ & ~_01957_;
	assign _01959_ = ~(_01413_ | _01333_);
	assign _01960_ = _01958_ & ~_01959_;
	assign _01961_ = ~(_01410_ | _01333_);
	assign _01962_ = _01960_ & ~_01961_;
	assign _01963_ = ~(_01408_ | _01333_);
	assign _01964_ = _01963_ | _01962_;
	assign _01966_ = _01331_ | ~_01417_;
	assign _01967_ = _01966_ & _01964_;
	assign _01968_ = _01942_ & ~_01967_;
	assign _01969_ = _01968_ | _01940_;
	assign _01970_ = _01969_ | _01939_;
	assign _01971_ = _01938_ & ~_01970_;
	assign _01972_ = _01971_ | _01937_;
	assign _01973_ = _01972_ | _01897_;
	assign _01974_ = ~(io_in[4] & io_in[5]);
	assign _01975_ = _01031_ & ~_01974_;
	assign _01977_ = ~(\mchip.wrapper.intxtReg.Q [8] & \mchip.wrapper.intxtReg.Q [9]);
	assign _01978_ = _06222_ & _00032_;
	assign _01979_ = _01977_ & ~_01978_;
	assign _01980_ = _00054_ & ~_06200_;
	assign _01981_ = _01979_ & ~_01980_;
	assign _01982_ = (_00153_ ? _06231_ : _01981_);
	assign _01983_ = _03074_ | _00010_;
	assign _01984_ = _03063_ & _00318_;
	assign _01985_ = _01983_ & ~_01984_;
	assign _01986_ = _03052_ & _00087_;
	assign _01988_ = _01985_ & ~_01986_;
	assign _01989_ = (_00131_ ? _06220_ : _01988_);
	assign _01990_ = _00547_ & ~_06201_;
	assign _01991_ = _00525_ & ~_01990_;
	assign _01992_ = _06200_ & _00569_;
	assign _01993_ = _01991_ & ~_01992_;
	assign _01994_ = (_00668_ ? _06211_ : _01993_);
	assign _01995_ = _00602_ | ~_03052_;
	assign _01996_ = _00833_ & ~_03063_;
	assign _01998_ = _00514_ | _01996_;
	assign _01999_ = _01995_ & ~_01998_;
	assign _02000_ = (_00646_ ? \mchip.wrapper.keyReg.Q [1] : _01999_);
	assign _02001_ = _02000_ ^ _01994_;
	assign _02002_ = _02001_ ^ _01989_;
	assign _02003_ = _02002_ ^ _01982_;
	assign _02004_ = _02003_ ^ \mchip.wrapper.intxtReg.Q [1];
	assign _02005_ = _02004_ ^ _03041_;
	assign _02006_ = _02005_ ^ _00052_;
	assign _02008_ = ~_06231_;
	assign _02009_ = ~_06223_;
	assign _02010_ = ~(_03052_ ^ \mchip.wrapper.intxtReg.Q [9]);
	assign _02011_ = ~_06466_;
	assign _02012_ = _06264_ | _02011_;
	assign _02013_ = _00032_ & ~_06263_;
	assign _02014_ = _02012_ & ~_02013_;
	assign _02015_ = _00054_ & ~_06241_;
	assign _02016_ = _02014_ & ~_02015_;
	assign _02017_ = (_00153_ ? _06280_ : _02016_);
	assign _02019_ = _06263_ & _00318_;
	assign _02020_ = _00010_ & ~_02019_;
	assign _02021_ = _00087_ & ~_06241_;
	assign _02022_ = _02020_ & ~_02021_;
	assign _02023_ = (_00131_ ? _06273_ : _02022_);
	assign _02024_ = _00086_ | _00525_;
	assign _02025_ = _00547_ & ~_03963_;
	assign _02026_ = _02024_ & ~_02025_;
	assign _02027_ = _03952_ & _00569_;
	assign _02029_ = _02026_ & ~_02027_;
	assign _02030_ = (_00668_ ? _06259_ : _02029_);
	assign _02031_ = _00602_ | ~_06241_;
	assign _02032_ = _06242_ & _00833_;
	assign _02033_ = _00514_ & ~_06243_;
	assign _02034_ = _02033_ | _02032_;
	assign _02035_ = _02031_ & ~_02034_;
	assign _02036_ = (_00646_ ? \mchip.wrapper.keyReg.Q [0] : _02035_);
	assign _02037_ = _02036_ ^ _02030_;
	assign _02038_ = _02037_ ^ _02023_;
	assign _02040_ = _02038_ ^ _02017_;
	assign _02041_ = _02040_ ^ \mchip.wrapper.intxtReg.Q [0];
	assign _02042_ = _02041_ ^ \mchip.wrapper.keyReg.Q [0];
	assign _02043_ = _02005_ | ~_02042_;
	assign _02044_ = _02043_ | _06223_;
	assign _02045_ = _02042_ | _02005_;
	assign _02046_ = _06222_ & ~_02045_;
	assign _02047_ = _02044_ & ~_02046_;
	assign _02048_ = ~(_02042_ & _02005_);
	assign _02049_ = _06206_ & ~_02048_;
	assign _02051_ = _02047_ & ~_02049_;
	assign _02052_ = _02005_ & ~_02042_;
	assign _02053_ = (_02052_ ? _06231_ : _02051_);
	assign _02054_ = _06111_ & _00032_;
	assign _02055_ = _01977_ & ~_02054_;
	assign _02056_ = _00054_ & ~_06110_;
	assign _02057_ = _02055_ & ~_02056_;
	assign _02058_ = (_00153_ ? _02616_ : _02057_);
	assign _02060_ = _00318_ & ~_03755_;
	assign _02061_ = _00010_ & ~_02060_;
	assign _02062_ = _00087_ & ~_03744_;
	assign _02063_ = _02061_ & ~_02062_;
	assign _02064_ = (_00131_ ? _06108_ : _02063_);
	assign _02065_ = _00547_ & ~_03755_;
	assign _02066_ = _00525_ & ~_02065_;
	assign _02067_ = _03744_ & _00569_;
	assign _02068_ = _02066_ & ~_02067_;
	assign _02070_ = (_00668_ ? _06099_ : _02068_);
	assign _02071_ = _00602_ | ~_03744_;
	assign _02072_ = _03755_ & _00833_;
	assign _02073_ = _00514_ | _02072_;
	assign _02074_ = _02071_ & ~_02073_;
	assign _02075_ = (_00646_ ? _03733_ : _02074_);
	assign _02076_ = _02075_ ^ _02070_;
	assign _02077_ = _02076_ ^ _02064_;
	assign _02078_ = _02077_ ^ _02058_;
	assign _02080_ = _02078_ ^ \mchip.wrapper.intxtReg.Q [3];
	assign _02081_ = _02080_ ^ \mchip.wrapper.keyReg.Q [3];
	assign _02082_ = _06162_ & _00032_;
	assign _02083_ = _01977_ & ~_02082_;
	assign _02084_ = _00054_ & ~_06130_;
	assign _02085_ = _02083_ & ~_02084_;
	assign _02086_ = (_00153_ ? _01188_ : _02085_);
	assign _02087_ = _00010_ | ~_06133_;
	assign _02088_ = _06131_ & _00318_;
	assign _02090_ = _02087_ & ~_02088_;
	assign _02091_ = _06130_ & _00087_;
	assign _02092_ = _02090_ & ~_02091_;
	assign _02093_ = (_00131_ ? _06160_ : _02092_);
	assign _02094_ = _06131_ & _00547_;
	assign _02095_ = _00525_ & ~_02094_;
	assign _02096_ = _06130_ & _00569_;
	assign _02097_ = _02095_ & ~_02096_;
	assign _02098_ = (_00668_ ? _01188_ : _02097_);
	assign _02100_ = _00602_ | ~_06130_;
	assign _02101_ = _06131_ & _00833_;
	assign _02102_ = _06133_ & _00514_;
	assign _02103_ = _02102_ | _02101_;
	assign _02104_ = _02100_ & ~_02103_;
	assign _02105_ = (_00646_ ? _06129_ : _02104_);
	assign _02106_ = _02105_ ^ _02098_;
	assign _02107_ = _02106_ ^ _02093_;
	assign _02108_ = _02107_ ^ _02086_;
	assign _02109_ = _02108_ ^ \mchip.wrapper.intxtReg.Q [2];
	assign _02111_ = _02109_ ^ _06129_;
	assign _02112_ = ~(_02111_ & _02081_);
	assign _02113_ = _02112_ | _03074_;
	assign _02114_ = ~_02081_;
	assign _02115_ = _02111_ | _02114_;
	assign _02116_ = _03063_ & ~_02115_;
	assign _02117_ = _02113_ & ~_02116_;
	assign _02118_ = ~(_02111_ & _02114_);
	assign _02119_ = _03052_ & ~_02118_;
	assign _02120_ = _02117_ & ~_02119_;
	assign _02122_ = _02114_ & ~_02111_;
	assign _02123_ = (_02122_ ? _06220_ : _02120_);
	assign _02124_ = _00032_ & ~_03470_;
	assign _02125_ = _01977_ & ~_02124_;
	assign _02126_ = _03459_ & _00054_;
	assign _02127_ = _02125_ & ~_02126_;
	assign _02128_ = (_00153_ ? _01735_ : _02127_);
	assign _02129_ = _00318_ & ~_04944_;
	assign _02131_ = _00010_ & ~_02129_;
	assign _02132_ = _04933_ & _00087_;
	assign _02133_ = _02131_ & ~_02132_;
	assign _02134_ = (_00131_ ? _05129_ : _02133_);
	assign _02135_ = _04955_ | _00525_;
	assign _02136_ = _00547_ & ~_04944_;
	assign _02137_ = _02135_ & ~_02136_;
	assign _02138_ = _04933_ & _00569_;
	assign _02139_ = _02137_ & ~_02138_;
	assign _02140_ = (_00668_ ? _05032_ : _02139_);
	assign _02142_ = _00602_ | ~_03459_;
	assign _02143_ = _03470_ & _00833_;
	assign _02144_ = _00514_ & ~_03481_;
	assign _02145_ = _02144_ | _02143_;
	assign _02146_ = _02142_ & ~_02145_;
	assign _02147_ = (_00646_ ? _04833_ : _02146_);
	assign _02148_ = _02147_ ^ _02140_;
	assign _02149_ = _02148_ ^ _02134_;
	assign _02150_ = _02149_ ^ _02128_;
	assign _02151_ = _02150_ ^ \mchip.wrapper.intxtReg.Q [5];
	assign _02153_ = _02151_ ^ \mchip.wrapper.keyReg.Q [5];
	assign _02154_ = _05646_ | _02011_;
	assign _02155_ = _00032_ & ~_05635_;
	assign _02156_ = _02154_ & ~_02155_;
	assign _02157_ = _00054_ & ~_03503_;
	assign _02158_ = _02156_ & ~_02157_;
	assign _02159_ = (_00153_ ? _05713_ : _02158_);
	assign _02160_ = _05537_ | _00010_;
	assign _02161_ = _00318_ & ~_05337_;
	assign _02162_ = _02160_ & ~_02161_;
	assign _02164_ = _05326_ & _00087_;
	assign _02165_ = _02162_ & ~_02164_;
	assign _02166_ = (_00131_ ? _01110_ : _02165_);
	assign _02167_ = _03525_ | _00525_;
	assign _02168_ = _00547_ & ~_03514_;
	assign _02169_ = _02167_ & ~_02168_;
	assign _02170_ = _03503_ & _00569_;
	assign _02171_ = _02169_ & ~_02170_;
	assign _02172_ = (_00668_ ? _05515_ : _02171_);
	assign _02173_ = _00602_ | ~_05326_;
	assign _02175_ = _05337_ & _00833_;
	assign _02176_ = _00514_ & ~_05348_;
	assign _02177_ = _02176_ | _02175_;
	assign _02178_ = _02173_ & ~_02177_;
	assign _02179_ = (_00646_ ? \mchip.wrapper.keyReg.Q [4] : _02178_);
	assign _02180_ = _02179_ ^ _02172_;
	assign _02181_ = _02180_ ^ _02166_;
	assign _02182_ = _02181_ ^ _02159_;
	assign _02183_ = _02182_ ^ \mchip.wrapper.intxtReg.Q [4];
	assign _02184_ = _02183_ ^ _05624_;
	assign _02186_ = _02184_ | _02153_;
	assign _02187_ = _02186_ | _06202_;
	assign _02188_ = _02183_ ^ \mchip.wrapper.keyReg.Q [4];
	assign _02189_ = _02188_ | _02153_;
	assign _02190_ = _00352_ & ~_02189_;
	assign _02191_ = _02187_ & ~_02190_;
	assign _02192_ = ~(_02188_ & _02153_);
	assign _02193_ = _06200_ & ~_02192_;
	assign _02194_ = _02191_ & ~_02193_;
	assign _02195_ = _02153_ & ~_02188_;
	assign _02197_ = (_02195_ ? _06211_ : _02194_);
	assign _02198_ = _00032_ & ~_03239_;
	assign _02199_ = _01977_ & ~_02198_;
	assign _02200_ = _00054_ & ~_03228_;
	assign _02201_ = _02199_ & ~_02200_;
	assign _02202_ = (_00153_ ? _04241_ : _02201_);
	assign _02203_ = _03239_ & _00318_;
	assign _02204_ = _00010_ & ~_02203_;
	assign _02206_ = _03228_ & _00087_;
	assign _02207_ = _02204_ & ~_02206_;
	assign _02208_ = (_00131_ ? _00996_ : _02207_);
	assign _02209_ = _03184_ | _00525_;
	assign _02210_ = _03173_ & _00547_;
	assign _02211_ = _02209_ & ~_02210_;
	assign _02212_ = _03162_ & _00569_;
	assign _02213_ = _02211_ & ~_02212_;
	assign _02214_ = (_00668_ ? _03667_ : _02213_);
	assign _02215_ = _00602_ | ~_03162_;
	assign _02217_ = _03206_ & _00833_;
	assign _02218_ = _00514_ & ~_03217_;
	assign _02219_ = _02218_ | _02217_;
	assign _02220_ = _02215_ & ~_02219_;
	assign _02221_ = (_00646_ ? _03195_ : _02220_);
	assign _02222_ = _02221_ ^ _02214_;
	assign _02223_ = _02222_ ^ _02208_;
	assign _02224_ = _02223_ ^ _02202_;
	assign _02225_ = _02224_ ^ \mchip.wrapper.intxtReg.Q [7];
	assign _02226_ = _02225_ ^ _03195_;
	assign _02228_ = ~(_03305_ & _06466_);
	assign _02229_ = _03294_ & _00032_;
	assign _02230_ = _02228_ & ~_02229_;
	assign _02231_ = _03283_ & _00054_;
	assign _02232_ = _02230_ & ~_02231_;
	assign _02233_ = (_00153_ ? _04558_ : _02232_);
	assign _02234_ = _03305_ | _00010_;
	assign _02235_ = _03294_ & _00318_;
	assign _02236_ = _02234_ & ~_02235_;
	assign _02237_ = _03283_ & _00087_;
	assign _02239_ = _02236_ & ~_02237_;
	assign _02240_ = (_00131_ ? _04558_ : _02239_);
	assign _02241_ = _03305_ | _00525_;
	assign _02242_ = _00547_ & ~_03294_;
	assign _02243_ = _02241_ & ~_02242_;
	assign _02244_ = _03283_ & _00569_;
	assign _02245_ = _02243_ & ~_02244_;
	assign _02246_ = (_00668_ ? _04471_ : _02245_);
	assign _02247_ = _00602_ | ~_03085_;
	assign _02248_ = _03129_ & _00833_;
	assign _02250_ = _00514_ & ~_03140_;
	assign _02251_ = _02250_ | _02248_;
	assign _02252_ = _02247_ & ~_02251_;
	assign _02253_ = (_00646_ ? _03107_ : _02252_);
	assign _02254_ = _02253_ ^ _02246_;
	assign _02255_ = _02254_ ^ _02240_;
	assign _02256_ = _02255_ ^ _02233_;
	assign _02257_ = _02256_ ^ \mchip.wrapper.intxtReg.Q [6];
	assign _02258_ = _02257_ ^ _03107_;
	assign _02259_ = _02258_ | _02226_;
	assign _02261_ = _03074_ & ~_02259_;
	assign _02262_ = _02257_ ^ \mchip.wrapper.keyReg.Q [6];
	assign _02263_ = _02262_ | _02226_;
	assign _02264_ = _00344_ & ~_02263_;
	assign _02265_ = _02264_ | _02261_;
	assign _02266_ = ~(_02262_ & _02226_);
	assign _02267_ = _03052_ & ~_02266_;
	assign _02268_ = _02267_ | _02265_;
	assign _02269_ = _02226_ & ~_02262_;
	assign _02270_ = (_02269_ ? _03041_ : _02268_);
	assign _02272_ = _02270_ ^ _02197_;
	assign _02273_ = _02272_ ^ _02123_;
	assign _02274_ = _02273_ ^ _02053_;
	assign _02275_ = _02274_ ^ _02010_;
	assign _02276_ = _02275_ ^ _00344_;
	assign _02277_ = _03952_ ^ \mchip.wrapper.intxtReg.Q [8];
	assign _02278_ = ~_06280_;
	assign _02280_ = _02279_ & ~_02043_;
	assign _02281_ = _06266_ & ~_02045_;
	assign _02283_ = _02281_ | _02280_;
	assign _02284_ = _06248_ & ~_02048_;
	assign _02285_ = _02284_ | _02283_;
	assign _02286_ = (_02052_ ? _02278_ : _02285_);
	assign _02287_ = _06264_ & ~_02112_;
	assign _02288_ = _06263_ & ~_02115_;
	assign _02289_ = _02288_ | _02287_;
	assign _02290_ = _06248_ & ~_02118_;
	assign _02291_ = _02290_ | _02289_;
	assign _02292_ = (_02122_ ? _06272_ : _02291_);
	assign _02294_ = _04122_ & ~_02186_;
	assign _02295_ = _00386_ & ~_02189_;
	assign _02296_ = _02295_ | _02294_;
	assign _02297_ = _03952_ & ~_02192_;
	assign _02298_ = _02297_ | _02296_;
	assign _02299_ = (_02195_ ? _06258_ : _02298_);
	assign _02300_ = _02266_ | _06248_;
	assign _02301_ = _00089_ & ~_02259_;
	assign _02302_ = _06242_ & ~_02263_;
	assign _02303_ = _02302_ | _02301_;
	assign _02305_ = _02300_ & ~_02303_;
	assign _02306_ = (_02269_ ? \mchip.wrapper.keyReg.Q [0] : _02305_);
	assign _02307_ = _02306_ ^ _02299_;
	assign _02308_ = _02307_ ^ _02292_;
	assign _02309_ = _02308_ ^ _02286_;
	assign _02310_ = _02309_ ^ _02277_;
	assign _02311_ = _02310_ ^ _00386_;
	assign _02312_ = ~(_02311_ & _02276_);
	assign _02313_ = _02009_ & ~_02312_;
	assign _02314_ = _02311_ | ~_02276_;
	assign _02316_ = _06222_ & ~_02314_;
	assign _02317_ = _02316_ | _02313_;
	assign _02318_ = _02276_ | ~_02311_;
	assign _02319_ = _06206_ & ~_02318_;
	assign _02320_ = _02319_ | _02317_;
	assign _02321_ = ~(_02311_ | _02276_);
	assign _02322_ = (_02321_ ? _02008_ : _02320_);
	assign _02323_ = ~(_03744_ ^ \mchip.wrapper.intxtReg.Q [11]);
	assign _02324_ = _02043_ | _06113_;
	assign _02325_ = _06111_ & ~_02045_;
	assign _02327_ = _02324_ & ~_02325_;
	assign _02328_ = _06462_ & ~_02048_;
	assign _02329_ = _02327_ & ~_02328_;
	assign _02330_ = (_02052_ ? _02616_ : _02329_);
	assign _02331_ = _02112_ | _05945_;
	assign _02332_ = _00271_ & ~_02115_;
	assign _02333_ = _02331_ & ~_02332_;
	assign _02334_ = _05911_ & ~_02118_;
	assign _02335_ = _02333_ & ~_02334_;
	assign _02336_ = (_02122_ ? _06108_ : _02335_);
	assign _02338_ = _02186_ | _05945_;
	assign _02339_ = _00271_ & ~_02189_;
	assign _02340_ = _02338_ & ~_02339_;
	assign _02341_ = _03744_ & ~_02192_;
	assign _02342_ = _02340_ & ~_02341_;
	assign _02343_ = (_02195_ ? _06099_ : _02342_);
	assign _02344_ = _05934_ & ~_02259_;
	assign _02345_ = _03755_ & ~_02263_;
	assign _02346_ = _02345_ | _02344_;
	assign _02347_ = _03744_ & ~_02266_;
	assign _02349_ = _02347_ | _02346_;
	assign _02350_ = (_02269_ ? \mchip.wrapper.keyReg.Q [3] : _02349_);
	assign _02351_ = _02350_ ^ _02343_;
	assign _02352_ = _02351_ ^ _02336_;
	assign _02353_ = _02352_ ^ _02330_;
	assign _02354_ = _02353_ ^ _02323_;
	assign _02355_ = _02354_ ^ _03755_;
	assign _02356_ = ~(_06130_ ^ \mchip.wrapper.intxtReg.Q [10]);
	assign _02357_ = _02043_ | _06163_;
	assign _02358_ = _06162_ & ~_02045_;
	assign _02360_ = _02357_ & ~_02358_;
	assign _02361_ = _06139_ & ~_02048_;
	assign _02362_ = _02360_ & ~_02361_;
	assign _02363_ = (_02052_ ? _01188_ : _02362_);
	assign _02364_ = _02112_ | _06134_;
	assign _02365_ = _06131_ & ~_02115_;
	assign _02366_ = _02364_ & ~_02365_;
	assign _02367_ = _06130_ & ~_02118_;
	assign _02368_ = _02366_ & ~_02367_;
	assign _02369_ = (_02122_ ? _06160_ : _02368_);
	assign _02371_ = _02186_ | _06146_;
	assign _02372_ = _06131_ & ~_02189_;
	assign _02373_ = _02371_ & ~_02372_;
	assign _02374_ = _06130_ & ~_02192_;
	assign _02375_ = _02373_ & ~_02374_;
	assign _02376_ = (_02195_ ? _01188_ : _02375_);
	assign _02377_ = _06133_ & ~_02259_;
	assign _02378_ = _06131_ & ~_02263_;
	assign _02379_ = _02378_ | _02377_;
	assign _02380_ = _06130_ & ~_02266_;
	assign _02382_ = _02380_ | _02379_;
	assign _02383_ = (_02269_ ? \mchip.wrapper.keyReg.Q [2] : _02382_);
	assign _02384_ = _02383_ ^ _02376_;
	assign _02385_ = _02384_ ^ _02369_;
	assign _02386_ = _02385_ ^ _02363_;
	assign _02387_ = _02386_ ^ _02356_;
	assign _02388_ = _02387_ ^ _06131_;
	assign _02389_ = ~(_02388_ & _02355_);
	assign _02390_ = _00051_ & ~_02389_;
	assign _02391_ = _02388_ | ~_02355_;
	assign _02393_ = _03063_ & ~_02391_;
	assign _02394_ = _02393_ | _02390_;
	assign _02395_ = _02355_ | ~_02388_;
	assign _02396_ = _03052_ & ~_02395_;
	assign _02397_ = _02396_ | _02394_;
	assign _02398_ = ~(_02388_ | _02355_);
	assign _02399_ = (_02398_ ? _06219_ : _02397_);
	assign _02400_ = ~_06202_;
	assign _02401_ = ~(_03503_ ^ \mchip.wrapper.intxtReg.Q [12]);
	assign _02402_ = _02043_ | _05646_;
	assign _02404_ = _06415_ & ~_02045_;
	assign _02405_ = _02402_ & ~_02404_;
	assign _02406_ = _05482_ & ~_02048_;
	assign _02407_ = _02405_ & ~_02406_;
	assign _02408_ = (_02052_ ? _05713_ : _02407_);
	assign _02409_ = _02112_ | _05537_;
	assign _02410_ = _05371_ & ~_02115_;
	assign _02411_ = _02409_ & ~_02410_;
	assign _02412_ = _05326_ & ~_02118_;
	assign _02413_ = _02411_ & ~_02412_;
	assign _02415_ = (_02122_ ? _01110_ : _02413_);
	assign _02416_ = _02186_ | _03525_;
	assign _02417_ = _00226_ & ~_02189_;
	assign _02418_ = _02416_ & ~_02417_;
	assign _02419_ = _03503_ & ~_02192_;
	assign _02420_ = _02418_ & ~_02419_;
	assign _02421_ = (_02195_ ? _05515_ : _02420_);
	assign _02422_ = _06393_ & ~_02259_;
	assign _02423_ = _05337_ & ~_02263_;
	assign _02424_ = _02423_ | _02422_;
	assign _02426_ = _05326_ & ~_02266_;
	assign _02427_ = _02426_ | _02424_;
	assign _02428_ = (_02269_ ? _05624_ : _02427_);
	assign _02429_ = _02428_ ^ _02421_;
	assign _02430_ = _02429_ ^ _02415_;
	assign _02431_ = _02430_ ^ _02408_;
	assign _02432_ = _02431_ ^ _02401_;
	assign _02433_ = _02432_ ^ _00226_;
	assign _02434_ = _03459_ ^ \mchip.wrapper.intxtReg.Q [13];
	assign _02435_ = ~_05152_;
	assign _02437_ = _02435_ & ~_02043_;
	assign _02438_ = _04855_ & ~_02045_;
	assign _02439_ = _02438_ | _02437_;
	assign _02440_ = _03459_ & ~_02048_;
	assign _02441_ = _02440_ | _02439_;
	assign _02442_ = (_02052_ ? _05129_ : _02441_);
	assign _02443_ = _04955_ & ~_02112_;
	assign _02444_ = _06371_ & ~_02115_;
	assign _02445_ = _02444_ | _02443_;
	assign _02446_ = _04933_ & ~_02118_;
	assign _02448_ = _02446_ | _02445_;
	assign _02449_ = (_02122_ ? _01735_ : _02448_);
	assign _02451_ = _02450_ & ~_02186_;
	assign _02452_ = _06371_ & ~_02189_;
	assign _02453_ = _02452_ | _02451_;
	assign _02454_ = _04933_ & ~_02192_;
	assign _02455_ = _02454_ | _02453_;
	assign _02456_ = (_02195_ ? _01727_ : _02455_);
	assign _02457_ = _02266_ | _04888_;
	assign _02459_ = _06355_ & ~_02259_;
	assign _02460_ = _03470_ & ~_02263_;
	assign _02461_ = _02460_ | _02459_;
	assign _02462_ = _02457_ & ~_02461_;
	assign _02463_ = (_02269_ ? _04833_ : _02462_);
	assign _02464_ = _02463_ ^ _02456_;
	assign _02465_ = _02464_ ^ _02449_;
	assign _02466_ = _02465_ ^ _02442_;
	assign _02467_ = _02466_ ^ _02434_;
	assign _02468_ = _02467_ ^ _06389_;
	assign _02470_ = _02468_ | _02433_;
	assign _02471_ = _02400_ & ~_02470_;
	assign _02472_ = _02432_ ^ _03514_;
	assign _02473_ = _02468_ | _02472_;
	assign _02474_ = _00352_ & ~_02473_;
	assign _02475_ = _02474_ | _02471_;
	assign _02476_ = ~(_02468_ & _02472_);
	assign _02477_ = _06200_ & ~_02476_;
	assign _02478_ = _02477_ | _02475_;
	assign _02479_ = _02468_ & ~_02472_;
	assign _02481_ = (_02479_ ? _06210_ : _02478_);
	assign _02482_ = _03162_ ^ \mchip.wrapper.intxtReg.Q [15];
	assign _02483_ = _03799_ & ~_02043_;
	assign _02484_ = _03832_ & ~_02045_;
	assign _02485_ = _02484_ | _02483_;
	assign _02486_ = _03876_ & ~_02048_;
	assign _02487_ = _02486_ | _02485_;
	assign _02488_ = (_02052_ ? _04230_ : _02487_);
	assign _02489_ = ~_00996_;
	assign _02490_ = _03799_ & ~_02112_;
	assign _02492_ = _03239_ & ~_02115_;
	assign _02493_ = _02492_ | _02490_;
	assign _02494_ = _03228_ & ~_02118_;
	assign _02495_ = _02494_ | _02493_;
	assign _02496_ = (_02122_ ? _02489_ : _02495_);
	assign _02497_ = ~_03667_;
	assign _02498_ = ~_03184_;
	assign _02499_ = _02498_ & ~_02186_;
	assign _02500_ = _03173_ & ~_02189_;
	assign _02501_ = _02500_ | _02499_;
	assign _02503_ = _03162_ & ~_02192_;
	assign _02504_ = _02503_ | _02501_;
	assign _02505_ = (_02195_ ? _02497_ : _02504_);
	assign _02506_ = _02266_ | _03382_;
	assign _02507_ = _03261_ & ~_02259_;
	assign _02508_ = _03206_ & ~_02263_;
	assign _02509_ = _02508_ | _02507_;
	assign _02510_ = _02506_ & ~_02509_;
	assign _02511_ = (_02269_ ? _03195_ : _02510_);
	assign _02512_ = _02511_ ^ _02505_;
	assign _02514_ = _02512_ ^ _02496_;
	assign _02515_ = _02514_ ^ _02488_;
	assign _02516_ = _02515_ ^ _02482_;
	assign _02517_ = _02516_ ^ _03173_;
	assign _02518_ = ~(_03085_ ^ \mchip.wrapper.intxtReg.Q [14]);
	assign _02519_ = _02043_ | _01835_;
	assign _02520_ = _03294_ & ~_02045_;
	assign _02521_ = _02519_ & ~_02520_;
	assign _02522_ = _03283_ & ~_02048_;
	assign _02523_ = _02521_ & ~_02522_;
	assign _02525_ = (_02052_ ? _04558_ : _02523_);
	assign _02526_ = _02112_ | _03305_;
	assign _02527_ = _03294_ & ~_02115_;
	assign _02528_ = _02526_ & ~_02527_;
	assign _02529_ = _03283_ & ~_02118_;
	assign _02530_ = _02528_ & ~_02529_;
	assign _02531_ = (_02122_ ? _04558_ : _02530_);
	assign _02532_ = _02186_ | _03305_;
	assign _02533_ = _04503_ & ~_02189_;
	assign _02534_ = _02532_ & ~_02533_;
	assign _02536_ = _03283_ & ~_02192_;
	assign _02537_ = _02534_ & ~_02536_;
	assign _02538_ = (_02195_ ? _04471_ : _02537_);
	assign _02539_ = _06308_ & ~_02259_;
	assign _02540_ = _03129_ & ~_02263_;
	assign _02541_ = _02540_ | _02539_;
	assign _02542_ = _03085_ & ~_02266_;
	assign _02543_ = _02542_ | _02541_;
	assign _02544_ = (_02269_ ? \mchip.wrapper.keyReg.Q [6] : _02543_);
	assign _02545_ = _02544_ ^ _02538_;
	assign _02547_ = _02545_ ^ _02531_;
	assign _02548_ = _02547_ ^ _02525_;
	assign _02549_ = _02548_ ^ _02518_;
	assign _02550_ = _02549_ ^ _06341_;
	assign _02551_ = ~(_02550_ & _02517_);
	assign _02552_ = _02551_ | _06191_;
	assign _02553_ = ~_06341_;
	assign _02554_ = _02549_ ^ _02553_;
	assign _02555_ = _02554_ | _02517_;
	assign _02556_ = _03074_ & ~_02555_;
	assign _02558_ = _02550_ | _02517_;
	assign _02559_ = _00344_ & ~_02558_;
	assign _02560_ = _02559_ | _02556_;
	assign _02561_ = _02552_ & ~_02560_;
	assign _02562_ = _02517_ & ~_02550_;
	assign _02563_ = (_02562_ ? \mchip.wrapper.keyReg.Q [1] : _02561_);
	assign _02564_ = _02563_ ^ _02481_;
	assign _02565_ = _02564_ ^ _02399_;
	assign _02566_ = _02565_ ^ _02322_;
	assign _02567_ = _02566_ ^ _02006_;
	assign _02569_ = _02567_ ^ _01236_;
	assign _02570_ = _02569_ ^ _03074_;
	assign _02571_ = _02276_ ^ _03052_;
	assign _02572_ = _02042_ ^ _00086_;
	assign _02573_ = _02279_ & ~_02312_;
	assign _02574_ = _06266_ & ~_02314_;
	assign _02575_ = _02574_ | _02573_;
	assign _02576_ = _06248_ & ~_02318_;
	assign _02577_ = _02576_ | _02575_;
	assign _02578_ = (_02321_ ? _02278_ : _02577_);
	assign _02580_ = _06264_ & ~_02389_;
	assign _02581_ = _06263_ & ~_02391_;
	assign _02582_ = _02581_ | _02580_;
	assign _02583_ = _06248_ & ~_02395_;
	assign _02584_ = _02583_ | _02582_;
	assign _02585_ = (_02398_ ? _06272_ : _02584_);
	assign _02586_ = _04122_ & ~_02470_;
	assign _02587_ = _00386_ & ~_02473_;
	assign _02588_ = _02587_ | _02586_;
	assign _02589_ = _03952_ & ~_02476_;
	assign _02591_ = _02589_ | _02588_;
	assign _02592_ = (_02479_ ? _06258_ : _02591_);
	assign _02593_ = _02551_ | _06248_;
	assign _02594_ = _00089_ & ~_02555_;
	assign _02595_ = _06242_ & ~_02558_;
	assign _02596_ = _02595_ | _02594_;
	assign _02597_ = _02593_ & ~_02596_;
	assign _02598_ = (_02562_ ? \mchip.wrapper.keyReg.Q [0] : _02597_);
	assign _02599_ = _02598_ ^ _02592_;
	assign _02600_ = _02599_ ^ _02585_;
	assign _02602_ = _02600_ ^ _02578_;
	assign _02603_ = _02602_ ^ _02572_;
	assign _02604_ = _02603_ ^ _01271_;
	assign _02605_ = ~(_02604_ & _02569_);
	assign _02606_ = _02009_ & ~_02605_;
	assign _02607_ = _02604_ | ~_02569_;
	assign _02608_ = _06222_ & ~_02607_;
	assign _02609_ = _02608_ | _02606_;
	assign _02610_ = _02569_ | ~_02604_;
	assign _02611_ = _06206_ & ~_02610_;
	assign _02613_ = _02611_ | _02609_;
	assign _02614_ = ~(_02604_ | _02569_);
	assign _02615_ = (_02614_ ? _02008_ : _02613_);
	assign _02617_ = _02081_ ^ _05945_;
	assign _02618_ = _02312_ | _06113_;
	assign _02619_ = _06111_ & ~_02314_;
	assign _02620_ = _02618_ & ~_02619_;
	assign _02621_ = _06462_ & ~_02318_;
	assign _02622_ = _02620_ & ~_02621_;
	assign _02624_ = (_02321_ ? _02616_ : _02622_);
	assign _02625_ = _02389_ | _05945_;
	assign _02626_ = _00271_ & ~_02391_;
	assign _02627_ = _02625_ & ~_02626_;
	assign _02628_ = _05911_ & ~_02395_;
	assign _02629_ = _02627_ & ~_02628_;
	assign _02630_ = (_02398_ ? _06108_ : _02629_);
	assign _02631_ = _02470_ | _05945_;
	assign _02632_ = _00271_ & ~_02473_;
	assign _02633_ = _02631_ & ~_02632_;
	assign _02635_ = _03744_ & ~_02476_;
	assign _02636_ = _02633_ & ~_02635_;
	assign _02637_ = (_02479_ ? _06099_ : _02636_);
	assign _02638_ = _05934_ & ~_02555_;
	assign _02639_ = _03755_ & ~_02558_;
	assign _02640_ = _02639_ | _02638_;
	assign _02641_ = _03744_ & ~_02551_;
	assign _02642_ = _02641_ | _02640_;
	assign _02643_ = (_02562_ ? \mchip.wrapper.keyReg.Q [3] : _02642_);
	assign _02644_ = _02643_ ^ _02637_;
	assign _02646_ = _02644_ ^ _02630_;
	assign _02647_ = _02646_ ^ _02624_;
	assign _02648_ = _02647_ ^ _02617_;
	assign _02649_ = _02648_ ^ _02616_;
	assign _02650_ = _02111_ ^ _06133_;
	assign _02651_ = ~_06163_;
	assign _02652_ = _02651_ & ~_02312_;
	assign _02653_ = _06162_ & ~_02314_;
	assign _02654_ = _02653_ | _02652_;
	assign _02655_ = _06139_ & ~_02318_;
	assign _02657_ = _02655_ | _02654_;
	assign _02658_ = (_02321_ ? _01189_ : _02657_);
	assign _02659_ = _06133_ & ~_02389_;
	assign _02660_ = _06131_ & ~_02391_;
	assign _02661_ = _02660_ | _02659_;
	assign _02662_ = _06130_ & ~_02395_;
	assign _02663_ = _02662_ | _02661_;
	assign _02664_ = (_02398_ ? _06159_ : _02663_);
	assign _02665_ = _06145_ & ~_02470_;
	assign _02666_ = _06131_ & ~_02473_;
	assign _02668_ = _02666_ | _02665_;
	assign _02669_ = _06130_ & ~_02476_;
	assign _02670_ = _02669_ | _02668_;
	assign _02671_ = (_02479_ ? _01189_ : _02670_);
	assign _02672_ = _02551_ | _06139_;
	assign _02673_ = _06133_ & ~_02555_;
	assign _02674_ = _06131_ & ~_02558_;
	assign _02675_ = _02674_ | _02673_;
	assign _02676_ = _02672_ & ~_02675_;
	assign _02677_ = (_02562_ ? _06129_ : _02676_);
	assign _02679_ = _02677_ ^ _02671_;
	assign _02680_ = _02679_ ^ _02664_;
	assign _02681_ = _02680_ ^ _02658_;
	assign _02682_ = _02681_ ^ _02650_;
	assign _02683_ = _02682_ ^ _01189_;
	assign _02684_ = ~(_02683_ & _02649_);
	assign _02685_ = _00051_ & ~_02684_;
	assign _02686_ = _02683_ | ~_02649_;
	assign _02687_ = _03063_ & ~_02686_;
	assign _02688_ = _02687_ | _02685_;
	assign _02690_ = _02649_ | ~_02683_;
	assign _02691_ = _03052_ & ~_02690_;
	assign _02692_ = _02691_ | _02688_;
	assign _02693_ = ~(_02683_ | _02649_);
	assign _02694_ = (_02693_ ? _06219_ : _02692_);
	assign _02695_ = ~(_02153_ ^ _06391_);
	assign _02696_ = _02435_ & ~_02312_;
	assign _02697_ = _04855_ & ~_02314_;
	assign _02698_ = _02697_ | _02696_;
	assign _02699_ = _03459_ & ~_02318_;
	assign _02701_ = _02699_ | _02698_;
	assign _02702_ = (_02321_ ? _05129_ : _02701_);
	assign _02703_ = _04955_ & ~_02389_;
	assign _02704_ = _06371_ & ~_02391_;
	assign _02705_ = _02704_ | _02703_;
	assign _02706_ = _04933_ & ~_02395_;
	assign _02707_ = _02706_ | _02705_;
	assign _02708_ = (_02398_ ? _01735_ : _02707_);
	assign _02709_ = _02450_ & ~_02470_;
	assign _02710_ = _06371_ & ~_02473_;
	assign _02712_ = _02710_ | _02709_;
	assign _02713_ = _04933_ & ~_02476_;
	assign _02714_ = _02713_ | _02712_;
	assign _02715_ = (_02479_ ? _01727_ : _02714_);
	assign _02716_ = _02551_ | _04888_;
	assign _02717_ = _06355_ & ~_02555_;
	assign _02718_ = _03470_ & ~_02558_;
	assign _02719_ = _02718_ | _02717_;
	assign _02720_ = _02716_ & ~_02719_;
	assign _02721_ = (_02562_ ? _04833_ : _02720_);
	assign _02723_ = _02721_ ^ _02715_;
	assign _02724_ = _02723_ ^ _02708_;
	assign _02725_ = _02724_ ^ _02702_;
	assign _02726_ = _02725_ ^ _02695_;
	assign _02727_ = _02726_ ^ _01076_;
	assign _02728_ = ~_01110_;
	assign _02729_ = _02184_ ^ _03525_;
	assign _02730_ = _02312_ | _05646_;
	assign _02731_ = _06415_ & ~_02314_;
	assign _02732_ = _02730_ & ~_02731_;
	assign _02734_ = _05482_ & ~_02318_;
	assign _02735_ = _02732_ & ~_02734_;
	assign _02736_ = (_02321_ ? _05713_ : _02735_);
	assign _02737_ = _02389_ | _05537_;
	assign _02738_ = _05371_ & ~_02391_;
	assign _02739_ = _02737_ & ~_02738_;
	assign _02740_ = _05326_ & ~_02395_;
	assign _02741_ = _02739_ & ~_02740_;
	assign _02742_ = (_02398_ ? _01110_ : _02741_);
	assign _02743_ = _02470_ | _03525_;
	assign _02745_ = _00226_ & ~_02473_;
	assign _02746_ = _02743_ & ~_02745_;
	assign _02747_ = _03503_ & ~_02476_;
	assign _02748_ = _02746_ & ~_02747_;
	assign _02749_ = (_02479_ ? _05515_ : _02748_);
	assign _02750_ = _06393_ & ~_02555_;
	assign _02751_ = _05337_ & ~_02558_;
	assign _02752_ = _02751_ | _02750_;
	assign _02753_ = _05326_ & ~_02551_;
	assign _02754_ = _02753_ | _02752_;
	assign _02756_ = (_02562_ ? _05624_ : _02754_);
	assign _02757_ = _02756_ ^ _02749_;
	assign _02758_ = _02757_ ^ _02742_;
	assign _02759_ = _02758_ ^ _02736_;
	assign _02760_ = _02759_ ^ _02729_;
	assign _02761_ = _02760_ ^ _02728_;
	assign _02762_ = _02761_ | _02727_;
	assign _02763_ = _02400_ & ~_02762_;
	assign _02764_ = _02760_ ^ _01110_;
	assign _02765_ = _02764_ | _02727_;
	assign _02767_ = _00352_ & ~_02765_;
	assign _02768_ = _02767_ | _02763_;
	assign _02769_ = ~(_02764_ & _02727_);
	assign _02770_ = _06200_ & ~_02769_;
	assign _02771_ = _02770_ | _02768_;
	assign _02772_ = _02727_ & ~_02764_;
	assign _02773_ = (_02772_ ? _06210_ : _02771_);
	assign _02774_ = ~(_02226_ ^ _03184_);
	assign _02775_ = _03799_ & ~_02312_;
	assign _02776_ = _03832_ & ~_02314_;
	assign _02778_ = _02776_ | _02775_;
	assign _02779_ = _03876_ & ~_02318_;
	assign _02780_ = _02779_ | _02778_;
	assign _02781_ = (_02321_ ? _04230_ : _02780_);
	assign _02782_ = _03799_ & ~_02389_;
	assign _02783_ = _03239_ & ~_02391_;
	assign _02784_ = _02783_ | _02782_;
	assign _02785_ = _03228_ & ~_02395_;
	assign _02786_ = _02785_ | _02784_;
	assign _02787_ = (_02398_ ? _02489_ : _02786_);
	assign _02789_ = _02498_ & ~_02470_;
	assign _02790_ = _03173_ & ~_02473_;
	assign _02791_ = _02790_ | _02789_;
	assign _02792_ = _03162_ & ~_02476_;
	assign _02793_ = _02792_ | _02791_;
	assign _02794_ = (_02479_ ? _02497_ : _02793_);
	assign _02795_ = _02551_ | _03382_;
	assign _02796_ = _03261_ & ~_02555_;
	assign _02797_ = _03206_ & ~_02558_;
	assign _02798_ = _02797_ | _02796_;
	assign _02800_ = _02795_ & ~_02798_;
	assign _02801_ = (_02562_ ? _03195_ : _02800_);
	assign _02802_ = _02801_ ^ _02794_;
	assign _02803_ = _02802_ ^ _02787_;
	assign _02804_ = _02803_ ^ _02781_;
	assign _02805_ = _02804_ ^ _02774_;
	assign _02806_ = _02805_ ^ _00996_;
	assign _02807_ = _02258_ ^ _06342_;
	assign _02808_ = _02312_ | _01835_;
	assign _02809_ = _03294_ & ~_02314_;
	assign _02811_ = _02808_ & ~_02809_;
	assign _02812_ = _03283_ & ~_02318_;
	assign _02813_ = _02811_ & ~_02812_;
	assign _02814_ = (_02321_ ? _04558_ : _02813_);
	assign _02815_ = _02389_ | _03305_;
	assign _02816_ = _03294_ & ~_02391_;
	assign _02817_ = _02815_ & ~_02816_;
	assign _02818_ = _03283_ & ~_02395_;
	assign _02819_ = _02817_ & ~_02818_;
	assign _02820_ = (_02398_ ? _04558_ : _02819_);
	assign _02822_ = _02470_ | _03305_;
	assign _02823_ = _04503_ & ~_02473_;
	assign _02824_ = _02822_ & ~_02823_;
	assign _02825_ = _03283_ & ~_02476_;
	assign _02826_ = _02824_ & ~_02825_;
	assign _02827_ = (_02479_ ? _04471_ : _02826_);
	assign _02828_ = _06308_ & ~_02555_;
	assign _02829_ = _03129_ & ~_02558_;
	assign _02830_ = _02829_ | _02828_;
	assign _02831_ = _03085_ & ~_02551_;
	assign _02833_ = _02831_ | _02830_;
	assign _02834_ = (_02562_ ? \mchip.wrapper.keyReg.Q [6] : _02833_);
	assign _02835_ = _02834_ ^ _02827_;
	assign _02836_ = _02835_ ^ _02820_;
	assign _02837_ = _02836_ ^ _02814_;
	assign _02838_ = _02837_ ^ _02807_;
	assign _02839_ = _02838_ ^ _01030_;
	assign _02840_ = ~(_02839_ & _02806_);
	assign _02841_ = _02840_ | _06191_;
	assign _02842_ = ~_01030_;
	assign _02844_ = _02838_ ^ _02842_;
	assign _02845_ = _02844_ | _02806_;
	assign _02846_ = _03074_ & ~_02845_;
	assign _02847_ = _02839_ | _02806_;
	assign _02848_ = _00344_ & ~_02847_;
	assign _02849_ = _02848_ | _02846_;
	assign _02850_ = _02841_ & ~_02849_;
	assign _02851_ = _02806_ & ~_02839_;
	assign _02852_ = (_02851_ ? \mchip.wrapper.keyReg.Q [1] : _02850_);
	assign _02853_ = _02852_ ^ _02773_;
	assign _02855_ = _02853_ ^ _02694_;
	assign _02856_ = _02855_ ^ _02615_;
	assign _02857_ = _02856_ ^ _02571_;
	assign _02858_ = _02857_ ^ _00344_;
	assign _02859_ = _02311_ ^ _03952_;
	assign _02860_ = _02279_ & ~_02605_;
	assign _02861_ = _06266_ & ~_02607_;
	assign _02862_ = _02861_ | _02860_;
	assign _02863_ = _06248_ & ~_02610_;
	assign _02864_ = _02863_ | _02862_;
	assign _02866_ = (_02614_ ? _02278_ : _02864_);
	assign _02867_ = _06264_ & ~_02684_;
	assign _02868_ = _06263_ & ~_02686_;
	assign _02869_ = _02868_ | _02867_;
	assign _02870_ = _06248_ & ~_02690_;
	assign _02871_ = _02870_ | _02869_;
	assign _02872_ = (_02693_ ? _06272_ : _02871_);
	assign _02873_ = _04122_ & ~_02762_;
	assign _02874_ = _00386_ & ~_02765_;
	assign _02875_ = _02874_ | _02873_;
	assign _02877_ = _03952_ & ~_02769_;
	assign _02878_ = _02877_ | _02875_;
	assign _02879_ = (_02772_ ? _06258_ : _02878_);
	assign _02880_ = _02840_ | _06248_;
	assign _02881_ = _00089_ & ~_02845_;
	assign _02882_ = _06242_ & ~_02847_;
	assign _02883_ = _02882_ | _02881_;
	assign _02884_ = _02880_ & ~_02883_;
	assign _02885_ = (_02851_ ? \mchip.wrapper.keyReg.Q [0] : _02884_);
	assign _02886_ = _02885_ ^ _02879_;
	assign _02888_ = _02886_ ^ _02872_;
	assign _02889_ = _02888_ ^ _02866_;
	assign _02890_ = _02889_ ^ _02859_;
	assign _02891_ = _02890_ ^ _00386_;
	assign _02892_ = ~(_02891_ & _02858_);
	assign _02893_ = _02892_ | _06223_;
	assign _02894_ = _02891_ | ~_02858_;
	assign _02895_ = _06222_ & ~_02894_;
	assign _02896_ = _02893_ & ~_02895_;
	assign _02897_ = _02858_ | ~_02891_;
	assign _02899_ = _06206_ & ~_02897_;
	assign _02900_ = _02896_ & ~_02899_;
	assign _02901_ = ~(_02891_ | _02858_);
	assign _02902_ = (_02901_ ? _06231_ : _02900_);
	assign _02903_ = _02355_ ^ _03744_;
	assign _02904_ = ~(_02605_ | _06113_);
	assign _02905_ = _06111_ & ~_02607_;
	assign _02906_ = _02905_ | _02904_;
	assign _02907_ = _06462_ & ~_02610_;
	assign _02908_ = _02907_ | _02906_;
	assign _02910_ = (_02614_ ? _06099_ : _02908_);
	assign _02911_ = _05934_ & ~_02684_;
	assign _02912_ = _00271_ & ~_02686_;
	assign _02913_ = _02912_ | _02911_;
	assign _02914_ = _05911_ & ~_02690_;
	assign _02915_ = _02914_ | _02913_;
	assign _02916_ = (_02693_ ? _06107_ : _02915_);
	assign _02917_ = _05934_ & ~_02762_;
	assign _02918_ = _00271_ & ~_02765_;
	assign _02919_ = _02918_ | _02917_;
	assign _02921_ = _03744_ & ~_02769_;
	assign _02922_ = _02921_ | _02919_;
	assign _02923_ = (_02772_ ? _02616_ : _02922_);
	assign _02924_ = _02840_ | _05911_;
	assign _02925_ = _05934_ & ~_02845_;
	assign _02926_ = _03755_ & ~_02847_;
	assign _02927_ = _02926_ | _02925_;
	assign _02928_ = _02924_ & ~_02927_;
	assign _02929_ = (_02851_ ? _03733_ : _02928_);
	assign _02930_ = _02929_ ^ _02923_;
	assign _02932_ = _02930_ ^ _02916_;
	assign _02933_ = _02932_ ^ _02910_;
	assign _02934_ = _02933_ ^ _02903_;
	assign _02935_ = _02934_ ^ _00271_;
	assign _02936_ = _02388_ ^ _03689_;
	assign _02937_ = _02651_ & ~_02605_;
	assign _02938_ = _06162_ & ~_02607_;
	assign _02939_ = _02938_ | _02937_;
	assign _02940_ = _06139_ & ~_02610_;
	assign _02941_ = _02940_ | _02939_;
	assign _02943_ = (_02614_ ? _01189_ : _02941_);
	assign _02944_ = _06133_ & ~_02684_;
	assign _02945_ = _06131_ & ~_02686_;
	assign _02946_ = _02945_ | _02944_;
	assign _02947_ = _06130_ & ~_02690_;
	assign _02948_ = _02947_ | _02946_;
	assign _02949_ = (_02693_ ? _06159_ : _02948_);
	assign _02950_ = _06145_ & ~_02762_;
	assign _02951_ = _06131_ & ~_02765_;
	assign _02952_ = _02951_ | _02950_;
	assign _02954_ = _06130_ & ~_02769_;
	assign _02955_ = _02954_ | _02952_;
	assign _02956_ = (_02772_ ? _01189_ : _02955_);
	assign _02957_ = _02840_ | _06139_;
	assign _02958_ = _06133_ & ~_02845_;
	assign _02959_ = _06131_ & ~_02847_;
	assign _02960_ = _02959_ | _02958_;
	assign _02961_ = _02957_ & ~_02960_;
	assign _02962_ = (_02851_ ? _06129_ : _02961_);
	assign _02963_ = _02962_ ^ _02956_;
	assign _02965_ = _02963_ ^ _02949_;
	assign _02966_ = _02965_ ^ _02943_;
	assign _02967_ = _02966_ ^ _02936_;
	assign _02968_ = ~(_02967_ ^ _03700_);
	assign _02969_ = ~(_02968_ & _02935_);
	assign _02970_ = _02969_ | _03074_;
	assign _02971_ = _02968_ | ~_02935_;
	assign _02972_ = _03063_ & ~_02971_;
	assign _02973_ = _02970_ & ~_02972_;
	assign _02974_ = _02935_ | ~_02968_;
	assign _02976_ = _03052_ & ~_02974_;
	assign _02977_ = _02973_ & ~_02976_;
	assign _02978_ = ~(_02968_ | _02935_);
	assign _02979_ = (_02978_ ? _06220_ : _02977_);
	assign _02980_ = _02468_ ^ _04888_;
	assign _02981_ = _02435_ & ~_02605_;
	assign _02982_ = _04855_ & ~_02607_;
	assign _02983_ = _02982_ | _02981_;
	assign _02984_ = _03459_ & ~_02610_;
	assign _02985_ = _02984_ | _02983_;
	assign _02987_ = (_02614_ ? _05129_ : _02985_);
	assign _02988_ = _04955_ & ~_02684_;
	assign _02989_ = _06371_ & ~_02686_;
	assign _02990_ = _02989_ | _02988_;
	assign _02991_ = _04933_ & ~_02690_;
	assign _02992_ = _02991_ | _02990_;
	assign _02993_ = (_02693_ ? _01735_ : _02992_);
	assign _02994_ = _02450_ & ~_02762_;
	assign _02995_ = _06371_ & ~_02765_;
	assign _02996_ = _02995_ | _02994_;
	assign _02998_ = _04933_ & ~_02769_;
	assign _02999_ = _02998_ | _02996_;
	assign _03000_ = (_02772_ ? _01727_ : _02999_);
	assign _03001_ = _02840_ | _04888_;
	assign _03002_ = _06355_ & ~_02845_;
	assign _03003_ = _03470_ & ~_02847_;
	assign _03004_ = _03003_ | _03002_;
	assign _03005_ = _03001_ & ~_03004_;
	assign _03006_ = (_02851_ ? _04833_ : _03005_);
	assign _03007_ = _03006_ ^ _03000_;
	assign _03009_ = _03007_ ^ _02993_;
	assign _03010_ = _03009_ ^ _02987_;
	assign _03011_ = _03010_ ^ _02980_;
	assign _03012_ = _03011_ ^ _03470_;
	assign _03013_ = _02472_ ^ _05482_;
	assign _03014_ = _02605_ | _05646_;
	assign _03015_ = _06415_ & ~_02607_;
	assign _03016_ = _03014_ & ~_03015_;
	assign _03017_ = _05482_ & ~_02610_;
	assign _03018_ = _03016_ & ~_03017_;
	assign _03020_ = (_02614_ ? _05713_ : _03018_);
	assign _03021_ = _02684_ | _05537_;
	assign _03022_ = _05371_ & ~_02686_;
	assign _03023_ = _03021_ & ~_03022_;
	assign _03024_ = _05326_ & ~_02690_;
	assign _03025_ = _03023_ & ~_03024_;
	assign _03026_ = (_02693_ ? _01110_ : _03025_);
	assign _03027_ = _02762_ | _03525_;
	assign _03028_ = _00226_ & ~_02765_;
	assign _03029_ = _03027_ & ~_03028_;
	assign _03031_ = _03503_ & ~_02769_;
	assign _03032_ = _03029_ & ~_03031_;
	assign _03033_ = (_02772_ ? _05515_ : _03032_);
	assign _03034_ = _06393_ & ~_02845_;
	assign _03035_ = _05337_ & ~_02847_;
	assign _03036_ = _03035_ | _03034_;
	assign _03037_ = _05326_ & ~_02840_;
	assign _03038_ = _03037_ | _03036_;
	assign _03039_ = (_02851_ ? _05624_ : _03038_);
	assign _03040_ = _03039_ ^ _03033_;
	assign _03042_ = _03040_ ^ _03026_;
	assign _03043_ = _03042_ ^ _03020_;
	assign _03044_ = _03043_ ^ _03013_;
	assign _03045_ = _03044_ ^ _00226_;
	assign _03046_ = _03045_ | _03012_;
	assign _03047_ = _03046_ | _06202_;
	assign _03048_ = _03011_ ^ _04855_;
	assign _03049_ = ~(_03048_ & _03045_);
	assign _03050_ = _00352_ & ~_03049_;
	assign _03051_ = _03047_ & ~_03050_;
	assign _03053_ = _03048_ | _03045_;
	assign _03054_ = _06200_ & ~_03053_;
	assign _03055_ = _03051_ & ~_03054_;
	assign _03056_ = _03045_ & ~_03048_;
	assign _03057_ = (_03056_ ? _06211_ : _03055_);
	assign _03058_ = _02517_ ^ _03876_;
	assign _03059_ = _03799_ & ~_02605_;
	assign _03060_ = _03832_ & ~_02607_;
	assign _03061_ = _03060_ | _03059_;
	assign _03062_ = _03876_ & ~_02610_;
	assign _03064_ = _03062_ | _03061_;
	assign _03065_ = (_02614_ ? _04230_ : _03064_);
	assign _03066_ = _03799_ & ~_02684_;
	assign _03067_ = _03239_ & ~_02686_;
	assign _03068_ = _03067_ | _03066_;
	assign _03069_ = _03228_ & ~_02690_;
	assign _03070_ = _03069_ | _03068_;
	assign _03071_ = (_02693_ ? _02489_ : _03070_);
	assign _03072_ = _02498_ & ~_02762_;
	assign _03073_ = _03173_ & ~_02765_;
	assign _03075_ = _03073_ | _03072_;
	assign _03076_ = _03162_ & ~_02769_;
	assign _03077_ = _03076_ | _03075_;
	assign _03078_ = (_02772_ ? _02497_ : _03077_);
	assign _03079_ = _02840_ | _03382_;
	assign _03080_ = _03261_ & ~_02845_;
	assign _03081_ = _03206_ & ~_02847_;
	assign _03082_ = _03081_ | _03080_;
	assign _03083_ = _03079_ & ~_03082_;
	assign _03084_ = (_02851_ ? _03195_ : _03083_);
	assign _03086_ = _03084_ ^ _03078_;
	assign _03087_ = _03086_ ^ _03071_;
	assign _03088_ = _03087_ ^ _03065_;
	assign _03089_ = _03088_ ^ _03058_;
	assign _03090_ = _03089_ ^ _03239_;
	assign _03091_ = _02550_ ^ _03283_;
	assign _03092_ = _03305_ & ~_02605_;
	assign _03093_ = _03294_ & ~_02607_;
	assign _03094_ = _03093_ | _03092_;
	assign _03095_ = _03283_ & ~_02610_;
	assign _03097_ = _03095_ | _03094_;
	assign _03098_ = (_02614_ ? _01834_ : _03097_);
	assign _03099_ = _01835_ & ~_02684_;
	assign _03100_ = _03294_ & ~_02686_;
	assign _03101_ = _03100_ | _03099_;
	assign _03102_ = _03283_ & ~_02690_;
	assign _03103_ = _03102_ | _03101_;
	assign _03104_ = (_02693_ ? _01834_ : _03103_);
	assign _03105_ = _01835_ & ~_02762_;
	assign _03106_ = _04503_ & ~_02765_;
	assign _03108_ = _03106_ | _03105_;
	assign _03109_ = _03283_ & ~_02769_;
	assign _03110_ = _03109_ | _03108_;
	assign _03111_ = (_02772_ ? _01826_ : _03110_);
	assign _03112_ = _02840_ | _03096_;
	assign _03113_ = _06308_ & ~_02845_;
	assign _03114_ = _03129_ & ~_02847_;
	assign _03115_ = _03114_ | _03113_;
	assign _03116_ = _03112_ & ~_03115_;
	assign _03117_ = (_02851_ ? _03107_ : _03116_);
	assign _03119_ = _03117_ ^ _03111_;
	assign _03120_ = _03119_ ^ _03104_;
	assign _03121_ = _03120_ ^ _03098_;
	assign _03122_ = _03121_ ^ _03091_;
	assign _03123_ = _03122_ ^ _03294_;
	assign _03124_ = _03123_ | _03090_;
	assign _03125_ = _03074_ & ~_03124_;
	assign _03126_ = _03089_ ^ _03832_;
	assign _03127_ = ~(_03126_ & _03123_);
	assign _03128_ = _00344_ & ~_03127_;
	assign _03130_ = _03128_ | _03125_;
	assign _03131_ = _03126_ | _03123_;
	assign _03132_ = _03052_ & ~_03131_;
	assign _03133_ = _03132_ | _03130_;
	assign _03134_ = _03123_ & ~_03126_;
	assign _03135_ = (_03134_ ? _03041_ : _03133_);
	assign _03136_ = _03135_ ^ _03057_;
	assign _03137_ = _03136_ ^ _02979_;
	assign _03138_ = _03137_ ^ _02902_;
	assign _03139_ = _03138_ ^ _02570_;
	assign _03141_ = _03139_ ^ \mchip.wrapper.keyReg.Q [1];
	assign _03142_ = _03141_ ^ _00052_;
	assign _03143_ = _02858_ ^ _06191_;
	assign _03144_ = _02604_ ^ _00086_;
	assign _03145_ = _02892_ | _06264_;
	assign _03146_ = _06266_ & ~_02894_;
	assign _03147_ = _03145_ & ~_03146_;
	assign _03148_ = _06248_ & ~_02897_;
	assign _03149_ = _03147_ & ~_03148_;
	assign _03150_ = (_02901_ ? _06280_ : _03149_);
	assign _03152_ = _02969_ | _02279_;
	assign _03153_ = _06263_ & ~_02971_;
	assign _03154_ = _03152_ & ~_03153_;
	assign _03155_ = _06248_ & ~_02974_;
	assign _03156_ = _03154_ & ~_03155_;
	assign _03157_ = (_02978_ ? _06273_ : _03156_);
	assign _03158_ = _03046_ | _00086_;
	assign _03159_ = _00386_ & ~_03049_;
	assign _03160_ = _03158_ & ~_03159_;
	assign _03161_ = _03952_ & ~_03053_;
	assign _03163_ = _03160_ & ~_03161_;
	assign _03164_ = (_03056_ ? _06259_ : _03163_);
	assign _03165_ = _00089_ & ~_03124_;
	assign _03166_ = _06242_ & ~_03127_;
	assign _03167_ = _03166_ | _03165_;
	assign _03168_ = _06241_ & ~_03131_;
	assign _03169_ = _03168_ | _03167_;
	assign _03170_ = (_03134_ ? _06262_ : _03169_);
	assign _03171_ = _03170_ ^ _03164_;
	assign _03172_ = _03171_ ^ _03157_;
	assign _03174_ = _03172_ ^ _03150_;
	assign _03175_ = _03174_ ^ _03144_;
	assign _03176_ = _03175_ ^ \mchip.wrapper.keyReg.Q [0];
	assign _03177_ = ~(_03176_ & _03141_);
	assign _03178_ = _03177_ | _06223_;
	assign _03179_ = _03176_ | ~_03141_;
	assign _03180_ = _06222_ & ~_03179_;
	assign _03181_ = _03178_ & ~_03180_;
	assign _03182_ = _03141_ | ~_03176_;
	assign _03183_ = _06206_ & ~_03182_;
	assign _03185_ = _03181_ & ~_03183_;
	assign _03186_ = ~(_03176_ | _03141_);
	assign _03187_ = (_03186_ ? _06231_ : _03185_);
	assign _03188_ = _02649_ ^ _00554_;
	assign _03189_ = _02892_ | _06113_;
	assign _03190_ = _06111_ & ~_02894_;
	assign _03191_ = _03189_ & ~_03190_;
	assign _03192_ = _06462_ & ~_02897_;
	assign _03193_ = _03191_ & ~_03192_;
	assign _03194_ = (_02901_ ? _02616_ : _03193_);
	assign _03196_ = _02969_ | _05945_;
	assign _03197_ = _00271_ & ~_02971_;
	assign _03198_ = _03196_ & ~_03197_;
	assign _03199_ = _05911_ & ~_02974_;
	assign _03200_ = _03198_ & ~_03199_;
	assign _03201_ = (_02978_ ? _06108_ : _03200_);
	assign _03202_ = _03046_ | _05945_;
	assign _03203_ = _00271_ & ~_03049_;
	assign _03204_ = _03202_ & ~_03203_;
	assign _03205_ = _03744_ & ~_03053_;
	assign _03207_ = _03204_ & ~_03205_;
	assign _03208_ = (_03056_ ? _06099_ : _03207_);
	assign _03209_ = _05934_ & ~_03124_;
	assign _03210_ = _03755_ & ~_03127_;
	assign _03211_ = _03210_ | _03209_;
	assign _03212_ = _03744_ & ~_03131_;
	assign _03213_ = _03212_ | _03211_;
	assign _03214_ = (_03134_ ? \mchip.wrapper.keyReg.Q [3] : _03213_);
	assign _03215_ = _03214_ ^ _03208_;
	assign _03216_ = _03215_ ^ _03201_;
	assign _03218_ = _03216_ ^ _03194_;
	assign _03219_ = _03218_ ^ _03188_;
	assign _03220_ = _03219_ ^ \mchip.wrapper.keyReg.Q [3];
	assign _03221_ = _02683_ ^ _00588_;
	assign _03222_ = _02892_ | _06163_;
	assign _03223_ = _06162_ & ~_02894_;
	assign _03224_ = _03222_ & ~_03223_;
	assign _03225_ = _06139_ & ~_02897_;
	assign _03226_ = _03224_ & ~_03225_;
	assign _03227_ = (_02901_ ? _01188_ : _03226_);
	assign _03229_ = _02969_ | _06134_;
	assign _03230_ = _06131_ & ~_02971_;
	assign _03231_ = _03229_ & ~_03230_;
	assign _03232_ = _06130_ & ~_02974_;
	assign _03233_ = _03231_ & ~_03232_;
	assign _03234_ = (_02978_ ? _06160_ : _03233_);
	assign _03235_ = _03046_ | _06146_;
	assign _03236_ = _06131_ & ~_03049_;
	assign _03237_ = _03235_ & ~_03236_;
	assign _03238_ = _06130_ & ~_03053_;
	assign _03240_ = _03237_ & ~_03238_;
	assign _03241_ = (_03056_ ? _01188_ : _03240_);
	assign _03242_ = _06133_ & ~_03124_;
	assign _03243_ = _06131_ & ~_03127_;
	assign _03244_ = _03243_ | _03242_;
	assign _03245_ = _06130_ & ~_03131_;
	assign _03246_ = _03245_ | _03244_;
	assign _03247_ = (_03134_ ? \mchip.wrapper.keyReg.Q [2] : _03246_);
	assign _03248_ = _03247_ ^ _03241_;
	assign _03249_ = _03248_ ^ _03234_;
	assign _03251_ = _03249_ ^ _03227_;
	assign _03252_ = _03251_ ^ _03221_;
	assign _03253_ = _03252_ ^ _06129_;
	assign _03254_ = ~(_03253_ & _03220_);
	assign _03255_ = _03254_ | _03074_;
	assign _03256_ = _03253_ | ~_03220_;
	assign _03257_ = _03063_ & ~_03256_;
	assign _03258_ = _03255_ & ~_03257_;
	assign _03259_ = _03220_ | ~_03253_;
	assign _03260_ = _03052_ & ~_03259_;
	assign _03262_ = _03258_ & ~_03260_;
	assign _03263_ = ~(_03253_ | _03220_);
	assign _03264_ = (_03263_ ? _06220_ : _03262_);
	assign _03265_ = _02727_ ^ _06355_;
	assign _03266_ = _02892_ | _05152_;
	assign _03267_ = _04855_ & ~_02894_;
	assign _03268_ = _03266_ & ~_03267_;
	assign _03269_ = _03459_ & ~_02897_;
	assign _03270_ = _03268_ & ~_03269_;
	assign _03271_ = (_02901_ ? _01735_ : _03270_);
	assign _03273_ = _02969_ | _02450_;
	assign _03274_ = _06371_ & ~_02971_;
	assign _03275_ = _03273_ & ~_03274_;
	assign _03276_ = _04933_ & ~_02974_;
	assign _03277_ = _03275_ & ~_03276_;
	assign _03278_ = (_02978_ ? _05129_ : _03277_);
	assign _03279_ = _03046_ | _04955_;
	assign _03280_ = _06371_ & ~_03049_;
	assign _03281_ = _03279_ & ~_03280_;
	assign _03282_ = _04933_ & ~_03053_;
	assign _03284_ = _03281_ & ~_03282_;
	assign _03285_ = (_03056_ ? _05032_ : _03284_);
	assign _03286_ = _06355_ & ~_03124_;
	assign _03287_ = _03470_ & ~_03127_;
	assign _03288_ = _03287_ | _03286_;
	assign _03289_ = _03459_ & ~_03131_;
	assign _03290_ = _03289_ | _03288_;
	assign _03291_ = (_03134_ ? \mchip.wrapper.keyReg.Q [5] : _03290_);
	assign _03292_ = _03291_ ^ _03285_;
	assign _03293_ = _03292_ ^ _03278_;
	assign _03295_ = _03293_ ^ _03271_;
	assign _03296_ = _03295_ ^ _03265_;
	assign _03297_ = _03296_ ^ \mchip.wrapper.keyReg.Q [5];
	assign _03298_ = _02764_ ^ _03525_;
	assign _03299_ = _02892_ | _05646_;
	assign _03300_ = _06415_ & ~_02894_;
	assign _03301_ = _03299_ & ~_03300_;
	assign _03302_ = _05482_ & ~_02897_;
	assign _03303_ = _03301_ & ~_03302_;
	assign _03304_ = (_02901_ ? _05713_ : _03303_);
	assign _03306_ = _02969_ | _05537_;
	assign _03307_ = _05371_ & ~_02971_;
	assign _03308_ = _03306_ & ~_03307_;
	assign _03309_ = _05326_ & ~_02974_;
	assign _03310_ = _03308_ & ~_03309_;
	assign _03311_ = (_02978_ ? _01110_ : _03310_);
	assign _03312_ = _03046_ | _03525_;
	assign _03313_ = _00226_ & ~_03049_;
	assign _03314_ = _03312_ & ~_03313_;
	assign _03315_ = _03503_ & ~_03053_;
	assign _03317_ = _03314_ & ~_03315_;
	assign _03318_ = (_03056_ ? _05515_ : _03317_);
	assign _03319_ = _06393_ & ~_03124_;
	assign _03320_ = _05337_ & ~_03127_;
	assign _03321_ = _03320_ | _03319_;
	assign _03322_ = _05326_ & ~_03131_;
	assign _03323_ = _03322_ | _03321_;
	assign _03324_ = (_03134_ ? _05624_ : _03323_);
	assign _03325_ = _03324_ ^ _03318_;
	assign _03326_ = _03325_ ^ _03311_;
	assign _03328_ = _03326_ ^ _03304_;
	assign _03329_ = _03328_ ^ _03298_;
	assign _03330_ = _03329_ ^ _05624_;
	assign _03331_ = _03330_ | _03297_;
	assign _03332_ = _03331_ | _06202_;
	assign _03333_ = _03296_ ^ _04833_;
	assign _03334_ = ~(_03333_ & _03330_);
	assign _03335_ = _00352_ & ~_03334_;
	assign _03336_ = _03332_ & ~_03335_;
	assign _03337_ = _03333_ | _03330_;
	assign _03339_ = _06200_ & ~_03337_;
	assign _03340_ = _03336_ & ~_03339_;
	assign _03341_ = _03330_ & ~_03333_;
	assign _03342_ = (_03341_ ? _06211_ : _03340_);
	assign _03343_ = _02806_ ^ _03250_;
	assign _03344_ = _02892_ | _03810_;
	assign _03345_ = _03832_ & ~_02894_;
	assign _03346_ = _03344_ & ~_03345_;
	assign _03347_ = _03876_ & ~_02897_;
	assign _03348_ = _03346_ & ~_03347_;
	assign _03350_ = (_02901_ ? _04241_ : _03348_);
	assign _03351_ = _02969_ | _03810_;
	assign _03352_ = _03239_ & ~_02971_;
	assign _03353_ = _03351_ & ~_03352_;
	assign _03354_ = _03228_ & ~_02974_;
	assign _03355_ = _03353_ & ~_03354_;
	assign _03356_ = (_02978_ ? _00996_ : _03355_);
	assign _03357_ = _03046_ | _03184_;
	assign _03358_ = _03173_ & ~_03049_;
	assign _03359_ = _03357_ & ~_03358_;
	assign _03361_ = _03162_ & ~_03053_;
	assign _03362_ = _03359_ & ~_03361_;
	assign _03363_ = (_03056_ ? _03667_ : _03362_);
	assign _03364_ = _03261_ & ~_03124_;
	assign _03365_ = _03206_ & ~_03127_;
	assign _03366_ = _03365_ | _03364_;
	assign _03367_ = _03162_ & ~_03131_;
	assign _03368_ = _03367_ | _03366_;
	assign _03369_ = (_03134_ ? \mchip.wrapper.keyReg.Q [7] : _03368_);
	assign _03370_ = _03369_ ^ _03363_;
	assign _03372_ = _03370_ ^ _03356_;
	assign _03373_ = _03372_ ^ _03350_;
	assign _03374_ = _03373_ ^ _03343_;
	assign _03375_ = _03374_ ^ _03195_;
	assign _03376_ = _02839_ ^ _01835_;
	assign _03377_ = _02892_ | _01835_;
	assign _03378_ = _03294_ & ~_02894_;
	assign _03379_ = _03377_ & ~_03378_;
	assign _03380_ = _03283_ & ~_02897_;
	assign _03381_ = _03379_ & ~_03380_;
	assign _03383_ = (_02901_ ? _04558_ : _03381_);
	assign _03384_ = _02969_ | _03305_;
	assign _03385_ = _03294_ & ~_02971_;
	assign _03386_ = _03384_ & ~_03385_;
	assign _03387_ = _03283_ & ~_02974_;
	assign _03388_ = _03386_ & ~_03387_;
	assign _03389_ = (_02978_ ? _04558_ : _03388_);
	assign _03390_ = _03046_ | _03305_;
	assign _03391_ = _04503_ & ~_03049_;
	assign _03392_ = _03390_ & ~_03391_;
	assign _03394_ = _03283_ & ~_03053_;
	assign _03395_ = _03392_ & ~_03394_;
	assign _03396_ = (_03056_ ? _04471_ : _03395_);
	assign _03397_ = _06308_ & ~_03124_;
	assign _03398_ = _03129_ & ~_03127_;
	assign _03399_ = _03398_ | _03397_;
	assign _03400_ = _03085_ & ~_03131_;
	assign _03401_ = _03400_ | _03399_;
	assign _03402_ = (_03134_ ? \mchip.wrapper.keyReg.Q [6] : _03401_);
	assign _03403_ = _03402_ ^ _03396_;
	assign _03405_ = _03403_ ^ _03389_;
	assign _03406_ = _03405_ ^ _03383_;
	assign _03407_ = _03406_ ^ _03376_;
	assign _03408_ = _03407_ ^ _03107_;
	assign _03409_ = _03408_ | _03375_;
	assign _03410_ = _03074_ & ~_03409_;
	assign _03411_ = _03374_ ^ \mchip.wrapper.keyReg.Q [7];
	assign _03412_ = ~(_03411_ & _03408_);
	assign _03413_ = _00344_ & ~_03412_;
	assign _03414_ = _03413_ | _03410_;
	assign _03416_ = _03411_ | _03408_;
	assign _03417_ = _03052_ & ~_03416_;
	assign _03418_ = _03417_ | _03414_;
	assign _03419_ = _03408_ & ~_03411_;
	assign _03420_ = (_03419_ ? _03041_ : _03418_);
	assign _03421_ = _03420_ ^ _03342_;
	assign _03422_ = _03421_ ^ _03264_;
	assign _03423_ = _03422_ ^ _03187_;
	assign _03424_ = _03423_ ^ _03143_;
	assign _03425_ = _03424_ ^ _00344_;
	assign _03427_ = _02891_ ^ _06240_;
	assign _03428_ = _03177_ | _06264_;
	assign _03429_ = _06266_ & ~_03179_;
	assign _03430_ = _03428_ & ~_03429_;
	assign _03431_ = _06248_ & ~_03182_;
	assign _03432_ = _03430_ & ~_03431_;
	assign _03433_ = (_03186_ ? _06280_ : _03432_);
	assign _03434_ = _03254_ | _02279_;
	assign _03435_ = _06263_ & ~_03256_;
	assign _03436_ = _03434_ & ~_03435_;
	assign _03438_ = _06248_ & ~_03259_;
	assign _03439_ = _03436_ & ~_03438_;
	assign _03440_ = (_03263_ ? _06273_ : _03439_);
	assign _03441_ = _03331_ | _00086_;
	assign _03442_ = _00386_ & ~_03334_;
	assign _03443_ = _03441_ & ~_03442_;
	assign _03444_ = _03952_ & ~_03337_;
	assign _03445_ = _03443_ & ~_03444_;
	assign _03446_ = (_03341_ ? _06259_ : _03445_);
	assign _03447_ = _00089_ & ~_03409_;
	assign _03449_ = _06242_ & ~_03412_;
	assign _03450_ = _03449_ | _03447_;
	assign _03451_ = _06241_ & ~_03416_;
	assign _03452_ = _03451_ | _03450_;
	assign _03453_ = (_03419_ ? _06262_ : _03452_);
	assign _03454_ = _03453_ ^ _03446_;
	assign _03455_ = _03454_ ^ _03440_;
	assign _03456_ = _03455_ ^ _03433_;
	assign _03457_ = _03456_ ^ _03427_;
	assign _03458_ = _03457_ ^ _03963_;
	assign _03460_ = ~(_03458_ & _03425_);
	assign _03461_ = _03460_ | _06223_;
	assign _03462_ = _03458_ | ~_03425_;
	assign _03463_ = _06222_ & ~_03462_;
	assign _03464_ = _03461_ & ~_03463_;
	assign _03465_ = _03425_ | ~_03458_;
	assign _03466_ = _06206_ & ~_03465_;
	assign _03467_ = _03464_ & ~_03466_;
	assign _03468_ = ~(_03458_ | _03425_);
	assign _03469_ = (_03468_ ? _06231_ : _03467_);
	assign _03471_ = _02935_ ^ _05911_;
	assign _03472_ = _03177_ | _06113_;
	assign _03473_ = _06111_ & ~_03179_;
	assign _03474_ = _03472_ & ~_03473_;
	assign _03475_ = _06462_ & ~_03182_;
	assign _03476_ = _03474_ & ~_03475_;
	assign _03477_ = (_03186_ ? _02616_ : _03476_);
	assign _03478_ = _03254_ | _05945_;
	assign _03479_ = _00271_ & ~_03256_;
	assign _03480_ = _03478_ & ~_03479_;
	assign _03482_ = _05911_ & ~_03259_;
	assign _03483_ = _03480_ & ~_03482_;
	assign _03484_ = (_03263_ ? _06108_ : _03483_);
	assign _03485_ = _03331_ | _05945_;
	assign _03486_ = _00271_ & ~_03334_;
	assign _03487_ = _03485_ & ~_03486_;
	assign _03488_ = _03744_ & ~_03337_;
	assign _03489_ = _03487_ & ~_03488_;
	assign _03490_ = (_03341_ ? _06099_ : _03489_);
	assign _03491_ = _05934_ & ~_03409_;
	assign _03493_ = _03755_ & ~_03412_;
	assign _03494_ = _03493_ | _03491_;
	assign _03495_ = _03744_ & ~_03416_;
	assign _03496_ = _03495_ | _03494_;
	assign _03497_ = (_03419_ ? \mchip.wrapper.keyReg.Q [3] : _03496_);
	assign _03498_ = _03497_ ^ _03490_;
	assign _03499_ = _03498_ ^ _03484_;
	assign _03500_ = _03499_ ^ _03477_;
	assign _03501_ = _03500_ ^ _03471_;
	assign _03502_ = _03501_ ^ _03755_;
	assign _03504_ = _02968_ ^ _06139_;
	assign _03505_ = _03177_ | _06163_;
	assign _03506_ = _06162_ & ~_03179_;
	assign _03507_ = _03505_ & ~_03506_;
	assign _03508_ = _06139_ & ~_03182_;
	assign _03509_ = _03507_ & ~_03508_;
	assign _03510_ = (_03186_ ? _01188_ : _03509_);
	assign _03511_ = _03254_ | _06134_;
	assign _03512_ = _06131_ & ~_03256_;
	assign _03513_ = _03511_ & ~_03512_;
	assign _03515_ = _06130_ & ~_03259_;
	assign _03516_ = _03513_ & ~_03515_;
	assign _03517_ = (_03263_ ? _06160_ : _03516_);
	assign _03518_ = _03331_ | _06146_;
	assign _03519_ = _06131_ & ~_03334_;
	assign _03520_ = _03518_ & ~_03519_;
	assign _03521_ = _06130_ & ~_03337_;
	assign _03522_ = _03520_ & ~_03521_;
	assign _03523_ = (_03341_ ? _01188_ : _03522_);
	assign _03524_ = _06133_ & ~_03409_;
	assign _03526_ = _06131_ & ~_03412_;
	assign _03527_ = _03526_ | _03524_;
	assign _03528_ = _06130_ & ~_03416_;
	assign _03529_ = _03528_ | _03527_;
	assign _03530_ = (_03419_ ? \mchip.wrapper.keyReg.Q [2] : _03529_);
	assign _03531_ = _03530_ ^ _03523_;
	assign _03532_ = _03531_ ^ _03517_;
	assign _03533_ = _03532_ ^ _03510_;
	assign _03534_ = _03533_ ^ _03504_;
	assign _03535_ = _03534_ ^ _06131_;
	assign _03537_ = ~(_03535_ & _03502_);
	assign _03538_ = _03537_ | _03074_;
	assign _03539_ = _03535_ | ~_03502_;
	assign _03540_ = _03063_ & ~_03539_;
	assign _03541_ = _03538_ & ~_03540_;
	assign _03542_ = _03502_ | ~_03535_;
	assign _03543_ = _03052_ & ~_03542_;
	assign _03544_ = _03541_ & ~_03543_;
	assign _03545_ = ~(_03535_ | _03502_);
	assign _03546_ = (_03545_ ? _06220_ : _03544_);
	assign _03548_ = _03012_ ^ _03459_;
	assign _03549_ = _03177_ | _05152_;
	assign _03550_ = _04855_ & ~_03179_;
	assign _03551_ = _03549_ & ~_03550_;
	assign _03552_ = _03459_ & ~_03182_;
	assign _03553_ = _03551_ & ~_03552_;
	assign _03554_ = (_03186_ ? _01735_ : _03553_);
	assign _03555_ = _03254_ | _02450_;
	assign _03556_ = _06371_ & ~_03256_;
	assign _03557_ = _03555_ & ~_03556_;
	assign _03558_ = _04933_ & ~_03259_;
	assign _03559_ = _03557_ & ~_03558_;
	assign _03560_ = (_03263_ ? _05129_ : _03559_);
	assign _03561_ = _03331_ | _04955_;
	assign _03562_ = _06371_ & ~_03334_;
	assign _03563_ = _03561_ & ~_03562_;
	assign _03564_ = _04933_ & ~_03337_;
	assign _03565_ = _03563_ & ~_03564_;
	assign _03566_ = (_03341_ ? _05032_ : _03565_);
	assign _03567_ = _06355_ & ~_03409_;
	assign _03569_ = _03470_ & ~_03412_;
	assign _03570_ = _03569_ | _03567_;
	assign _03571_ = _03459_ & ~_03416_;
	assign _03572_ = _03571_ | _03570_;
	assign _03573_ = (_03419_ ? \mchip.wrapper.keyReg.Q [5] : _03572_);
	assign _03574_ = _03573_ ^ _03566_;
	assign _03575_ = _03574_ ^ _03560_;
	assign _03576_ = _03575_ ^ _03554_;
	assign _03577_ = _03576_ ^ _03548_;
	assign _03578_ = ~(_03577_ ^ _06389_);
	assign _03580_ = _03045_ ^ _03503_;
	assign _03581_ = _03177_ | _05646_;
	assign _03582_ = _06415_ & ~_03179_;
	assign _03583_ = _03581_ & ~_03582_;
	assign _03584_ = _05482_ & ~_03182_;
	assign _03585_ = _03583_ & ~_03584_;
	assign _03586_ = (_03186_ ? _05713_ : _03585_);
	assign _03587_ = _03254_ | _05537_;
	assign _03588_ = _05371_ & ~_03256_;
	assign _03589_ = _03587_ & ~_03588_;
	assign _03591_ = _05326_ & ~_03259_;
	assign _03592_ = _03589_ & ~_03591_;
	assign _03593_ = (_03263_ ? _01110_ : _03592_);
	assign _03594_ = _03331_ | _03525_;
	assign _03595_ = _00226_ & ~_03334_;
	assign _03596_ = _03594_ & ~_03595_;
	assign _03597_ = _03503_ & ~_03337_;
	assign _03598_ = _03596_ & ~_03597_;
	assign _03599_ = (_03341_ ? _05515_ : _03598_);
	assign _03600_ = _06393_ & ~_03409_;
	assign _03602_ = _05337_ & ~_03412_;
	assign _03603_ = _03602_ | _03600_;
	assign _03604_ = _05326_ & ~_03416_;
	assign _03605_ = _03604_ | _03603_;
	assign _03606_ = (_03419_ ? _05624_ : _03605_);
	assign _03607_ = _03606_ ^ _03599_;
	assign _03608_ = _03607_ ^ _03593_;
	assign _03609_ = _03608_ ^ _03586_;
	assign _03610_ = _03609_ ^ _03580_;
	assign _03611_ = _03610_ ^ _00226_;
	assign _03613_ = _03611_ | _03578_;
	assign _03614_ = _03613_ | _06202_;
	assign _03615_ = _03577_ ^ _06389_;
	assign _03616_ = ~(_03615_ & _03611_);
	assign _03617_ = _00352_ & ~_03616_;
	assign _03618_ = _03614_ & ~_03617_;
	assign _03619_ = _03615_ | _03611_;
	assign _03620_ = _06200_ & ~_03619_;
	assign _03621_ = _03618_ & ~_03620_;
	assign _03622_ = _03611_ & ~_03615_;
	assign _03624_ = (_03622_ ? _06211_ : _03621_);
	assign _03625_ = _03090_ ^ _03162_;
	assign _03626_ = _03177_ | _03810_;
	assign _03627_ = _03832_ & ~_03179_;
	assign _03628_ = _03626_ & ~_03627_;
	assign _03629_ = _03876_ & ~_03182_;
	assign _03630_ = _03628_ & ~_03629_;
	assign _03631_ = (_03186_ ? _04241_ : _03630_);
	assign _03632_ = _03254_ | _03810_;
	assign _03633_ = _03239_ & ~_03256_;
	assign _03635_ = _03632_ & ~_03633_;
	assign _03636_ = _03228_ & ~_03259_;
	assign _03637_ = _03635_ & ~_03636_;
	assign _03638_ = (_03263_ ? _00996_ : _03637_);
	assign _03639_ = _03331_ | _03184_;
	assign _03640_ = _03173_ & ~_03334_;
	assign _03641_ = _03639_ & ~_03640_;
	assign _03642_ = _03162_ & ~_03337_;
	assign _03643_ = _03641_ & ~_03642_;
	assign _03644_ = (_03341_ ? _03667_ : _03643_);
	assign _03646_ = _03261_ & ~_03409_;
	assign _03647_ = _03206_ & ~_03412_;
	assign _03648_ = _03647_ | _03646_;
	assign _03649_ = _03162_ & ~_03416_;
	assign _03650_ = _03649_ | _03648_;
	assign _03651_ = (_03419_ ? \mchip.wrapper.keyReg.Q [7] : _03650_);
	assign _03652_ = _03651_ ^ _03644_;
	assign _03653_ = _03652_ ^ _03638_;
	assign _03654_ = _03653_ ^ _03631_;
	assign _03655_ = _03654_ ^ _03625_;
	assign _03657_ = _03655_ ^ _03579_;
	assign _03658_ = _03123_ ^ _03085_;
	assign _03659_ = _03177_ | _01835_;
	assign _03660_ = _03294_ & ~_03179_;
	assign _03661_ = _03659_ & ~_03660_;
	assign _03662_ = _03283_ & ~_03182_;
	assign _03663_ = _03661_ & ~_03662_;
	assign _03664_ = (_03186_ ? _04558_ : _03663_);
	assign _03665_ = _03254_ | _03305_;
	assign _03666_ = _03294_ & ~_03256_;
	assign _03668_ = _03665_ & ~_03666_;
	assign _03669_ = _03283_ & ~_03259_;
	assign _03670_ = _03668_ & ~_03669_;
	assign _03671_ = (_03263_ ? _04558_ : _03670_);
	assign _03672_ = _03331_ | _03305_;
	assign _03673_ = _04503_ & ~_03334_;
	assign _03674_ = _03672_ & ~_03673_;
	assign _03675_ = _03283_ & ~_03337_;
	assign _03676_ = _03674_ & ~_03675_;
	assign _03677_ = (_03341_ ? _04471_ : _03676_);
	assign _03679_ = _06308_ & ~_03409_;
	assign _03680_ = _03129_ & ~_03412_;
	assign _03681_ = _03680_ | _03679_;
	assign _03682_ = _03085_ & ~_03416_;
	assign _03683_ = _03682_ | _03681_;
	assign _03684_ = (_03419_ ? \mchip.wrapper.keyReg.Q [6] : _03683_);
	assign _03685_ = _03684_ ^ _03677_;
	assign _03686_ = _03685_ ^ _03671_;
	assign _03687_ = _03686_ ^ _03664_;
	assign _03688_ = _03687_ ^ _03658_;
	assign _03690_ = _03688_ ^ _02553_;
	assign _03691_ = _03690_ | _03657_;
	assign _03692_ = _03074_ & ~_03691_;
	assign _03693_ = _03655_ ^ _03173_;
	assign _03694_ = ~(_03693_ & _03690_);
	assign _03695_ = _00344_ & ~_03694_;
	assign _03696_ = _03695_ | _03692_;
	assign _03697_ = _03693_ | _03690_;
	assign _03698_ = _03052_ & ~_03697_;
	assign _03699_ = _03698_ | _03696_;
	assign _03701_ = _03690_ & ~_03693_;
	assign _03702_ = (_03701_ ? _03041_ : _03699_);
	assign _03703_ = _03702_ ^ _03624_;
	assign _03704_ = _03703_ ^ _03546_;
	assign _03705_ = _03704_ ^ _03469_;
	assign _03706_ = _03705_ ^ _03142_;
	assign _03707_ = _03706_ ^ _01235_;
	assign _03708_ = _03707_ ^ _00051_;
	assign _03709_ = _03176_ ^ _00088_;
	assign _03710_ = _03460_ | _06264_;
	assign _03712_ = _06266_ & ~_03462_;
	assign _03713_ = _03710_ & ~_03712_;
	assign _03714_ = _06248_ & ~_03465_;
	assign _03715_ = _03713_ & ~_03714_;
	assign _03716_ = (_03468_ ? _06280_ : _03715_);
	assign _03717_ = _03537_ | _02279_;
	assign _03718_ = _06263_ & ~_03539_;
	assign _03719_ = _03717_ & ~_03718_;
	assign _03720_ = _06248_ & ~_03542_;
	assign _03721_ = _03719_ & ~_03720_;
	assign _03723_ = (_03545_ ? _06273_ : _03721_);
	assign _03724_ = _03613_ | _00086_;
	assign _03725_ = _00386_ & ~_03616_;
	assign _03726_ = _03724_ & ~_03725_;
	assign _03727_ = _03952_ & ~_03619_;
	assign _03728_ = _03726_ & ~_03727_;
	assign _03729_ = (_03622_ ? _06259_ : _03728_);
	assign _03730_ = _00089_ & ~_03691_;
	assign _03731_ = _06242_ & ~_03694_;
	assign _03732_ = _03731_ | _03730_;
	assign _03734_ = _06241_ & ~_03697_;
	assign _03735_ = _03734_ | _03732_;
	assign _03736_ = (_03701_ ? _06262_ : _03735_);
	assign _03737_ = _03736_ ^ _03729_;
	assign _03738_ = _03737_ ^ _03723_;
	assign _03739_ = _03738_ ^ _03716_;
	assign _03740_ = _03739_ ^ _03709_;
	assign _03741_ = _03740_ ^ _01270_;
	assign _03742_ = _03741_ ^ _04122_;
	assign _03743_ = _03742_ & _03708_;
	assign _03745_ = _03220_ ^ _05945_;
	assign _03746_ = _03460_ | _06113_;
	assign _03747_ = _06111_ & ~_03462_;
	assign _03748_ = _03746_ & ~_03747_;
	assign _03749_ = _06462_ & ~_03465_;
	assign _03750_ = _03748_ & ~_03749_;
	assign _03751_ = (_03468_ ? _02616_ : _03750_);
	assign _03752_ = _03537_ | _05945_;
	assign _03753_ = _00271_ & ~_03539_;
	assign _03754_ = _03752_ & ~_03753_;
	assign _03756_ = _05911_ & ~_03542_;
	assign _03757_ = _03754_ & ~_03756_;
	assign _03758_ = (_03545_ ? _06108_ : _03757_);
	assign _03759_ = _03613_ | _05945_;
	assign _03760_ = _00271_ & ~_03616_;
	assign _03761_ = _03759_ & ~_03760_;
	assign _03762_ = _03744_ & ~_03619_;
	assign _03763_ = _03761_ & ~_03762_;
	assign _03764_ = (_03622_ ? _06099_ : _03763_);
	assign _03765_ = _05934_ & ~_03691_;
	assign _03767_ = _03755_ & ~_03694_;
	assign _03768_ = _03767_ | _03765_;
	assign _03769_ = _03744_ & ~_03697_;
	assign _03770_ = _03769_ | _03768_;
	assign _03771_ = (_03701_ ? \mchip.wrapper.keyReg.Q [3] : _03770_);
	assign _03772_ = _03771_ ^ _03764_;
	assign _03773_ = _03772_ ^ _03758_;
	assign _03774_ = _03773_ ^ _03751_;
	assign _03775_ = _03774_ ^ _03745_;
	assign _03776_ = _03775_ ^ _02616_;
	assign _03778_ = _03776_ ^ _03766_;
	assign _03779_ = _03253_ ^ _06134_;
	assign _03780_ = _03460_ | _06163_;
	assign _03781_ = _06162_ & ~_03462_;
	assign _03782_ = _03780_ & ~_03781_;
	assign _03783_ = _06139_ & ~_03465_;
	assign _03784_ = _03782_ & ~_03783_;
	assign _03785_ = (_03468_ ? _01188_ : _03784_);
	assign _03786_ = _03537_ | _06134_;
	assign _03787_ = _06131_ & ~_03539_;
	assign _03789_ = _03786_ & ~_03787_;
	assign _03790_ = _06130_ & ~_03542_;
	assign _03791_ = _03789_ & ~_03790_;
	assign _03792_ = (_03545_ ? _06160_ : _03791_);
	assign _03793_ = _03613_ | _06146_;
	assign _03794_ = _06131_ & ~_03616_;
	assign _03795_ = _03793_ & ~_03794_;
	assign _03796_ = _06130_ & ~_03619_;
	assign _03797_ = _03795_ & ~_03796_;
	assign _03798_ = (_03622_ ? _01188_ : _03797_);
	assign _03800_ = _06133_ & ~_03691_;
	assign _03801_ = _06131_ & ~_03694_;
	assign _03802_ = _03801_ | _03800_;
	assign _03803_ = _06130_ & ~_03697_;
	assign _03804_ = _03803_ | _03802_;
	assign _03805_ = (_03701_ ? \mchip.wrapper.keyReg.Q [2] : _03804_);
	assign _03806_ = _03805_ ^ _03798_;
	assign _03807_ = _03806_ ^ _03792_;
	assign _03808_ = _03807_ ^ _03785_;
	assign _03809_ = _03808_ ^ _03779_;
	assign _03811_ = _03809_ ^ _01188_;
	assign _03812_ = _03811_ ^ _03711_;
	assign _03813_ = ~(_03812_ & _03778_);
	assign _03814_ = _03743_ & ~_03813_;
	assign _03815_ = _03742_ | ~_03708_;
	assign _03816_ = ~(_03815_ | _03813_);
	assign _03817_ = _03708_ | ~_03742_;
	assign _03818_ = ~(_03817_ | _03813_);
	assign _03819_ = ~_03818_;
	assign _03820_ = _03778_ | ~_03812_;
	assign _03822_ = _03820_ | _03815_;
	assign _03823_ = ~(_03820_ | _03817_);
	assign _03824_ = _03812_ | _03778_;
	assign _03825_ = ~(_03824_ | _03817_);
	assign _03826_ = _03742_ | _03708_;
	assign _03827_ = ~(_03826_ | _03824_);
	assign _03828_ = _03825_ | ~_03827_;
	assign _03829_ = ~(_03824_ | _03815_);
	assign _03830_ = _03828_ & ~_03829_;
	assign _03831_ = _03743_ & ~_03824_;
	assign _03833_ = _03831_ | ~_03830_;
	assign _03834_ = ~(_03826_ | _03820_);
	assign _03835_ = _03833_ & ~_03834_;
	assign _03836_ = _03835_ | _03823_;
	assign _03837_ = _03822_ & ~_03836_;
	assign _03838_ = _03743_ & ~_03820_;
	assign _03839_ = _03837_ & ~_03838_;
	assign _03840_ = _03812_ | ~_03778_;
	assign _03841_ = ~(_03840_ | _03826_);
	assign _03842_ = _03839_ & ~_03841_;
	assign _03844_ = ~(_03840_ | _03817_);
	assign _03845_ = _03842_ & ~_03844_;
	assign _03846_ = ~(_03840_ | _03815_);
	assign _03847_ = _03845_ & ~_03846_;
	assign _03848_ = _03743_ & ~_03840_;
	assign _03849_ = _03848_ | _03847_;
	assign _03850_ = ~(_03826_ | _03813_);
	assign _03851_ = ~_03850_;
	assign _03852_ = _03851_ & _03849_;
	assign _03853_ = _03819_ & ~_03852_;
	assign _03855_ = _03853_ | _03816_;
	assign _03856_ = _03855_ | _03814_;
	assign _03857_ = _01975_ & ~_03856_;
	assign _03858_ = _04591_ & ~_01974_;
	assign _03859_ = _03297_ ^ _06391_;
	assign _03860_ = _03460_ | _05152_;
	assign _03861_ = _04855_ & ~_03462_;
	assign _03862_ = _03860_ & ~_03861_;
	assign _03863_ = _03459_ & ~_03465_;
	assign _03864_ = _03862_ & ~_03863_;
	assign _03866_ = (_03468_ ? _01735_ : _03864_);
	assign _03867_ = _03537_ | _02450_;
	assign _03868_ = _06371_ & ~_03539_;
	assign _03869_ = _03867_ & ~_03868_;
	assign _03870_ = _04933_ & ~_03542_;
	assign _03871_ = _03869_ & ~_03870_;
	assign _03872_ = (_03545_ ? _05129_ : _03871_);
	assign _03873_ = _03613_ | _04955_;
	assign _03874_ = _06371_ & ~_03616_;
	assign _03875_ = _03873_ & ~_03874_;
	assign _03877_ = _04933_ & ~_03619_;
	assign _03878_ = _03875_ & ~_03877_;
	assign _03879_ = (_03622_ ? _05032_ : _03878_);
	assign _03880_ = _06355_ & ~_03691_;
	assign _03881_ = _03470_ & ~_03694_;
	assign _03882_ = _03881_ | _03880_;
	assign _03883_ = _03459_ & ~_03697_;
	assign _03884_ = _03883_ | _03882_;
	assign _03885_ = (_03701_ ? \mchip.wrapper.keyReg.Q [5] : _03884_);
	assign _03886_ = _03885_ ^ _03879_;
	assign _03888_ = _03886_ ^ _03872_;
	assign _03889_ = _03888_ ^ _03866_;
	assign _03890_ = _03889_ ^ _03859_;
	assign _03891_ = ~(_03890_ ^ _01076_);
	assign _03892_ = _03891_ ^ _03481_;
	assign _03893_ = _03330_ ^ _03525_;
	assign _03894_ = _03460_ | _05646_;
	assign _03895_ = _06415_ & ~_03462_;
	assign _03896_ = _03894_ & ~_03895_;
	assign _03897_ = _05482_ & ~_03465_;
	assign _03899_ = _03896_ & ~_03897_;
	assign _03900_ = (_03468_ ? _05713_ : _03899_);
	assign _03901_ = _03537_ | _05537_;
	assign _03902_ = _05371_ & ~_03539_;
	assign _03903_ = _03901_ & ~_03902_;
	assign _03904_ = _05326_ & ~_03542_;
	assign _03905_ = _03903_ & ~_03904_;
	assign _03906_ = (_03545_ ? _01110_ : _03905_);
	assign _03907_ = _03613_ | _03525_;
	assign _03908_ = _00226_ & ~_03616_;
	assign _03910_ = _03907_ & ~_03908_;
	assign _03911_ = _03503_ & ~_03619_;
	assign _03912_ = _03910_ & ~_03911_;
	assign _03913_ = (_03622_ ? _05515_ : _03912_);
	assign _03914_ = _06393_ & ~_03691_;
	assign _03915_ = _05337_ & ~_03694_;
	assign _03916_ = _03915_ | _03914_;
	assign _03917_ = _05326_ & ~_03697_;
	assign _03918_ = _03917_ | _03916_;
	assign _03919_ = (_03701_ ? _05624_ : _03918_);
	assign _03921_ = _03919_ ^ _03913_;
	assign _03922_ = _03921_ ^ _03906_;
	assign _03923_ = _03922_ ^ _03900_;
	assign _03924_ = _03923_ ^ _03893_;
	assign _03925_ = _03924_ ^ _02728_;
	assign _03926_ = _03925_ ^ _03525_;
	assign _03927_ = _03926_ & _03892_;
	assign _03928_ = _03375_ ^ _03184_;
	assign _03929_ = _03460_ | _03810_;
	assign _03930_ = _03832_ & ~_03462_;
	assign _03931_ = _03929_ & ~_03930_;
	assign _03932_ = _03876_ & ~_03465_;
	assign _03933_ = _03931_ & ~_03932_;
	assign _03934_ = (_03468_ ? _04241_ : _03933_);
	assign _03935_ = _03537_ | _03810_;
	assign _03936_ = _03239_ & ~_03539_;
	assign _03937_ = _03935_ & ~_03936_;
	assign _03938_ = _03228_ & ~_03542_;
	assign _03939_ = _03937_ & ~_03938_;
	assign _03940_ = (_03545_ ? _00996_ : _03939_);
	assign _03942_ = _03613_ | _03184_;
	assign _03943_ = _03173_ & ~_03616_;
	assign _03944_ = _03942_ & ~_03943_;
	assign _03945_ = _03162_ & ~_03619_;
	assign _03946_ = _03944_ & ~_03945_;
	assign _03947_ = (_03622_ ? _03667_ : _03946_);
	assign _03948_ = _03261_ & ~_03691_;
	assign _03949_ = _03206_ & ~_03694_;
	assign _03950_ = _03949_ | _03948_;
	assign _03951_ = _03162_ & ~_03697_;
	assign _03953_ = _03951_ | _03950_;
	assign _03954_ = (_03701_ ? \mchip.wrapper.keyReg.Q [7] : _03953_);
	assign _03955_ = _03954_ ^ _03947_;
	assign _03956_ = _03955_ ^ _03940_;
	assign _03957_ = _03956_ ^ _03934_;
	assign _03958_ = _03957_ ^ _03928_;
	assign _03959_ = ~(_03958_ ^ _00996_);
	assign _03960_ = ~(_03959_ ^ _03250_);
	assign _03961_ = _03408_ ^ _06342_;
	assign _03962_ = _03460_ | _01835_;
	assign _03964_ = _03294_ & ~_03462_;
	assign _03965_ = _03962_ & ~_03964_;
	assign _03966_ = _03283_ & ~_03465_;
	assign _03967_ = _03965_ & ~_03966_;
	assign _03968_ = (_03468_ ? _04558_ : _03967_);
	assign _03969_ = _03537_ | _03305_;
	assign _03970_ = _03294_ & ~_03539_;
	assign _03971_ = _03969_ & ~_03970_;
	assign _03972_ = _03283_ & ~_03542_;
	assign _03973_ = _03971_ & ~_03972_;
	assign _03974_ = (_03545_ ? _04558_ : _03973_);
	assign _03975_ = _03613_ | _03305_;
	assign _03976_ = _04503_ & ~_03616_;
	assign _03977_ = _03975_ & ~_03976_;
	assign _03978_ = _03283_ & ~_03619_;
	assign _03979_ = _03977_ & ~_03978_;
	assign _03980_ = (_03622_ ? _04471_ : _03979_);
	assign _03981_ = _06308_ & ~_03691_;
	assign _03982_ = _03129_ & ~_03694_;
	assign _03983_ = _03982_ | _03981_;
	assign _03985_ = _03085_ & ~_03697_;
	assign _03986_ = _03985_ | _03983_;
	assign _03987_ = (_03701_ ? \mchip.wrapper.keyReg.Q [6] : _03986_);
	assign _03988_ = _03987_ ^ _03980_;
	assign _03989_ = _03988_ ^ _03974_;
	assign _03990_ = _03989_ ^ _03968_;
	assign _03991_ = _03990_ ^ _03961_;
	assign _03992_ = _03991_ ^ _02842_;
	assign _03993_ = _03992_ ^ _01835_;
	assign _03994_ = ~(_03993_ & _03960_);
	assign _03995_ = _03927_ & ~_03994_;
	assign _03996_ = _03926_ | ~_03892_;
	assign _03997_ = ~(_03996_ | _03994_);
	assign _03998_ = _03892_ | ~_03926_;
	assign _03999_ = ~(_03998_ | _03994_);
	assign _04000_ = ~_03999_;
	assign _04001_ = _03960_ | ~_03993_;
	assign _04002_ = _04001_ | _03996_;
	assign _04003_ = ~(_04001_ | _03998_);
	assign _04004_ = _03993_ | _03960_;
	assign _04005_ = ~(_04004_ | _03998_);
	assign _04006_ = _03926_ | _03892_;
	assign _04007_ = ~(_04006_ | _04004_);
	assign _04008_ = _04005_ | ~_04007_;
	assign _04009_ = ~(_04004_ | _03996_);
	assign _04010_ = _04008_ & ~_04009_;
	assign _04011_ = _03927_ & ~_04004_;
	assign _04012_ = _04011_ | ~_04010_;
	assign _04013_ = ~(_04006_ | _04001_);
	assign _04014_ = _04012_ & ~_04013_;
	assign _04016_ = _04014_ | _04003_;
	assign _04017_ = _04002_ & ~_04016_;
	assign _04018_ = _03927_ & ~_04001_;
	assign _04019_ = _04017_ & ~_04018_;
	assign _04020_ = _03993_ | ~_03960_;
	assign _04021_ = ~(_04020_ | _04006_);
	assign _04022_ = _04019_ & ~_04021_;
	assign _04023_ = ~(_04020_ | _03998_);
	assign _04024_ = _04022_ & ~_04023_;
	assign _04025_ = ~(_04020_ | _03996_);
	assign _04027_ = _04024_ & ~_04025_;
	assign _04028_ = _03927_ & ~_04020_;
	assign _04029_ = _04028_ | _04027_;
	assign _04030_ = ~(_04006_ | _03994_);
	assign _04031_ = ~_04030_;
	assign _04032_ = _04031_ & _04029_;
	assign _04033_ = _04000_ & ~_04032_;
	assign _04034_ = _04033_ | _03997_;
	assign _04035_ = _04034_ | _03995_;
	assign _04036_ = _03858_ & ~_04035_;
	assign _04037_ = _04036_ | _03857_;
	assign _04038_ = _06444_ & ~_01974_;
	assign _04039_ = _03425_ ^ _06191_;
	assign _04040_ = ~(_03741_ & _03707_);
	assign _04041_ = _04040_ | _06223_;
	assign _04042_ = _03741_ | ~_03707_;
	assign _04043_ = _06222_ & ~_04042_;
	assign _04044_ = _04041_ & ~_04043_;
	assign _04045_ = _03707_ | ~_03741_;
	assign _04046_ = _06206_ & ~_04045_;
	assign _04047_ = _04044_ & ~_04046_;
	assign _04048_ = ~(_03741_ | _03707_);
	assign _04049_ = (_04048_ ? _06231_ : _04047_);
	assign _04050_ = ~(_03811_ & _03776_);
	assign _04051_ = _04050_ | _03074_;
	assign _04052_ = _03811_ | ~_03776_;
	assign _04053_ = _03063_ & ~_04052_;
	assign _04054_ = _04051_ & ~_04053_;
	assign _04055_ = _03776_ | ~_03811_;
	assign _04056_ = _03052_ & ~_04055_;
	assign _04057_ = _04054_ & ~_04056_;
	assign _04058_ = ~(_03811_ | _03776_);
	assign _04059_ = (_04058_ ? _06220_ : _04057_);
	assign _04060_ = _03925_ | _03891_;
	assign _04061_ = _04060_ | _06202_;
	assign _04062_ = _03890_ ^ _01076_;
	assign _04063_ = ~(_04062_ & _03925_);
	assign _04064_ = _00352_ & ~_04063_;
	assign _04065_ = _04061_ & ~_04064_;
	assign _04066_ = _04062_ | _03925_;
	assign _04068_ = _06200_ & ~_04066_;
	assign _04069_ = _04065_ & ~_04068_;
	assign _04070_ = _03925_ & ~_04062_;
	assign _04071_ = (_04070_ ? _06211_ : _04069_);
	assign _04072_ = _03992_ | _03959_;
	assign _04073_ = _03074_ & ~_04072_;
	assign _04074_ = _03958_ ^ _00996_;
	assign _04075_ = ~(_04074_ & _03992_);
	assign _04076_ = _00344_ & ~_04075_;
	assign _04077_ = _04076_ | _04073_;
	assign _04079_ = _04074_ | _03992_;
	assign _04080_ = _03052_ & ~_04079_;
	assign _04081_ = _04080_ | _04077_;
	assign _04082_ = _03992_ & ~_04074_;
	assign _04083_ = (_04082_ ? _03041_ : _04081_);
	assign _04084_ = _04083_ ^ _04071_;
	assign _04085_ = _04084_ ^ _04059_;
	assign _04086_ = _04085_ ^ _04049_;
	assign _04087_ = _04086_ ^ _04039_;
	assign _04088_ = _04087_ ^ _03063_;
	assign _04090_ = _03458_ ^ _06240_;
	assign _04091_ = _04040_ | _06264_;
	assign _04092_ = _06266_ & ~_04042_;
	assign _04093_ = _04091_ & ~_04092_;
	assign _04094_ = _06248_ & ~_04045_;
	assign _04095_ = _04093_ & ~_04094_;
	assign _04096_ = (_04048_ ? _06280_ : _04095_);
	assign _04097_ = _04050_ | _02279_;
	assign _04098_ = _06263_ & ~_04052_;
	assign _04099_ = _04097_ & ~_04098_;
	assign _04101_ = _06248_ & ~_04055_;
	assign _04102_ = _04099_ & ~_04101_;
	assign _04103_ = (_04058_ ? _06273_ : _04102_);
	assign _04104_ = _04060_ | _00086_;
	assign _04105_ = _00386_ & ~_04063_;
	assign _04106_ = _04104_ & ~_04105_;
	assign _04107_ = _03952_ & ~_04066_;
	assign _04108_ = _04106_ & ~_04107_;
	assign _04109_ = (_04070_ ? _06259_ : _04108_);
	assign _04110_ = _00089_ & ~_04072_;
	assign _04112_ = _06242_ & ~_04075_;
	assign _04113_ = _04112_ | _04110_;
	assign _04114_ = _06241_ & ~_04079_;
	assign _04115_ = _04114_ | _04113_;
	assign _04116_ = (_04082_ ? _06262_ : _04115_);
	assign _04117_ = _04116_ ^ _04109_;
	assign _04118_ = _04117_ ^ _04103_;
	assign _04119_ = _04118_ ^ _04096_;
	assign _04120_ = _04119_ ^ _04090_;
	assign _04121_ = _04120_ ^ _00386_;
	assign _04123_ = _04088_ & ~_04121_;
	assign _04124_ = _03502_ ^ _05911_;
	assign _04125_ = _04040_ | _06113_;
	assign _04126_ = _06111_ & ~_04042_;
	assign _04127_ = _04125_ & ~_04126_;
	assign _04128_ = _06462_ & ~_04045_;
	assign _04129_ = _04127_ & ~_04128_;
	assign _04130_ = (_04048_ ? _02616_ : _04129_);
	assign _04131_ = _04050_ | _05945_;
	assign _04132_ = _00271_ & ~_04052_;
	assign _04134_ = _04131_ & ~_04132_;
	assign _04135_ = _05911_ & ~_04055_;
	assign _04136_ = _04134_ & ~_04135_;
	assign _04137_ = (_04058_ ? _06108_ : _04136_);
	assign _04138_ = _04060_ | _05945_;
	assign _04139_ = _00271_ & ~_04063_;
	assign _04140_ = _04138_ & ~_04139_;
	assign _04141_ = _03744_ & ~_04066_;
	assign _04142_ = _04140_ & ~_04141_;
	assign _04143_ = (_04070_ ? _06099_ : _04142_);
	assign _04145_ = _05934_ & ~_04072_;
	assign _04146_ = _03755_ & ~_04075_;
	assign _04147_ = _04146_ | _04145_;
	assign _04148_ = _03744_ & ~_04079_;
	assign _04149_ = _04148_ | _04147_;
	assign _04150_ = (_04082_ ? \mchip.wrapper.keyReg.Q [3] : _04149_);
	assign _04151_ = _04150_ ^ _04143_;
	assign _04152_ = _04151_ ^ _04137_;
	assign _04153_ = _04152_ ^ _04130_;
	assign _04154_ = _04153_ ^ _04124_;
	assign _04155_ = _04154_ ^ _03755_;
	assign _04156_ = _03535_ ^ _06128_;
	assign _04157_ = _04040_ | _06163_;
	assign _04158_ = _06162_ & ~_04042_;
	assign _04159_ = _04157_ & ~_04158_;
	assign _04160_ = _06139_ & ~_04045_;
	assign _04161_ = _04159_ & ~_04160_;
	assign _04162_ = (_04048_ ? _01188_ : _04161_);
	assign _04163_ = _04050_ | _06134_;
	assign _04164_ = _06131_ & ~_04052_;
	assign _04166_ = _04163_ & ~_04164_;
	assign _04167_ = _06130_ & ~_04055_;
	assign _04168_ = _04166_ & ~_04167_;
	assign _04169_ = (_04058_ ? _06160_ : _04168_);
	assign _04170_ = _04060_ | _06146_;
	assign _04171_ = _06131_ & ~_04063_;
	assign _04172_ = _04170_ & ~_04171_;
	assign _04173_ = _06130_ & ~_04066_;
	assign _04174_ = _04172_ & ~_04173_;
	assign _04175_ = (_04070_ ? _01188_ : _04174_);
	assign _04177_ = _06133_ & ~_04072_;
	assign _04178_ = _06131_ & ~_04075_;
	assign _04179_ = _04178_ | _04177_;
	assign _04180_ = _06130_ & ~_04079_;
	assign _04181_ = _04180_ | _04179_;
	assign _04182_ = (_04082_ ? \mchip.wrapper.keyReg.Q [2] : _04181_);
	assign _04183_ = _04182_ ^ _04175_;
	assign _04184_ = _04183_ ^ _04169_;
	assign _04185_ = _04184_ ^ _04162_;
	assign _04186_ = _04185_ ^ _04156_;
	assign _04188_ = _04186_ ^ _03700_;
	assign _04189_ = ~(_04188_ & _04155_);
	assign _04190_ = _04123_ & ~_04189_;
	assign _04191_ = ~(_04121_ & _04088_);
	assign _04192_ = ~(_04191_ | _04189_);
	assign _04193_ = _04121_ | _04088_;
	assign _04194_ = ~(_04193_ | _04189_);
	assign _04195_ = ~_04194_;
	assign _04196_ = _04155_ | ~_04188_;
	assign _04197_ = _04196_ | ~_04123_;
	assign _04199_ = ~(_04196_ | _04193_);
	assign _04200_ = _04188_ | _04155_;
	assign _04201_ = _04200_ | _04193_;
	assign _04202_ = _04088_ | ~_04121_;
	assign _04203_ = ~(_04202_ | _04200_);
	assign _04204_ = ~(_04203_ & _04201_);
	assign _04205_ = ~(_04200_ | _04191_);
	assign _04206_ = _04204_ & ~_04205_;
	assign _04207_ = _04123_ & ~_04200_;
	assign _04208_ = _04207_ | ~_04206_;
	assign _04210_ = ~(_04202_ | _04196_);
	assign _04211_ = _04208_ & ~_04210_;
	assign _04212_ = _04211_ | _04199_;
	assign _04213_ = _04196_ | _04191_;
	assign _04214_ = _04213_ & ~_04212_;
	assign _04215_ = _04214_ & _04197_;
	assign _04216_ = _04188_ | ~_04155_;
	assign _04217_ = ~(_04216_ | _04202_);
	assign _04218_ = _04215_ & ~_04217_;
	assign _04219_ = ~(_04216_ | _04193_);
	assign _04220_ = _04218_ & ~_04219_;
	assign _04221_ = ~(_04216_ | _04191_);
	assign _04222_ = _04220_ & ~_04221_;
	assign _04223_ = _04123_ & ~_04216_;
	assign _04224_ = _04223_ | _04222_;
	assign _04225_ = _04202_ | _04189_;
	assign _04226_ = _04225_ & _04224_;
	assign _04227_ = _04195_ & ~_04226_;
	assign _04228_ = _04227_ | _04192_;
	assign _04229_ = _04228_ | _04190_;
	assign _04231_ = _04038_ & ~_04229_;
	assign _04232_ = _00492_ & ~_01974_;
	assign _04233_ = _03578_ ^ _03459_;
	assign _04234_ = _04040_ | _05152_;
	assign _04235_ = _04855_ & ~_04042_;
	assign _04236_ = _04234_ & ~_04235_;
	assign _04237_ = _03459_ & ~_04045_;
	assign _04238_ = _04236_ & ~_04237_;
	assign _04239_ = (_04048_ ? _01735_ : _04238_);
	assign _04240_ = _04050_ | _02450_;
	assign _04242_ = _06371_ & ~_04052_;
	assign _04243_ = _04240_ & ~_04242_;
	assign _04244_ = _04933_ & ~_04055_;
	assign _04245_ = _04243_ & ~_04244_;
	assign _04246_ = (_04058_ ? _05129_ : _04245_);
	assign _04247_ = _04060_ | _04955_;
	assign _04248_ = _06371_ & ~_04063_;
	assign _04249_ = _04247_ & ~_04248_;
	assign _04250_ = _04933_ & ~_04066_;
	assign _04251_ = _04249_ & ~_04250_;
	assign _04253_ = (_04070_ ? _05032_ : _04251_);
	assign _04254_ = _06355_ & ~_04072_;
	assign _04255_ = _03470_ & ~_04075_;
	assign _04256_ = _04255_ | _04254_;
	assign _04257_ = _03459_ & ~_04079_;
	assign _04258_ = _04257_ | _04256_;
	assign _04259_ = (_04082_ ? \mchip.wrapper.keyReg.Q [5] : _04258_);
	assign _04260_ = _04259_ ^ _04253_;
	assign _04261_ = _04260_ ^ _04246_;
	assign _04262_ = _04261_ ^ _04239_;
	assign _04264_ = _04262_ ^ _04233_;
	assign _04265_ = _04264_ ^ _03470_;
	assign _04266_ = _03611_ ^ _03503_;
	assign _04267_ = _04040_ | _05646_;
	assign _04268_ = _06415_ & ~_04042_;
	assign _04269_ = _04267_ & ~_04268_;
	assign _04270_ = _05482_ & ~_04045_;
	assign _04271_ = _04269_ & ~_04270_;
	assign _04272_ = (_04048_ ? _05713_ : _04271_);
	assign _04273_ = _04050_ | _05537_;
	assign _04275_ = _05371_ & ~_04052_;
	assign _04276_ = _04273_ & ~_04275_;
	assign _04277_ = _05326_ & ~_04055_;
	assign _04278_ = _04276_ & ~_04277_;
	assign _04279_ = (_04058_ ? _01110_ : _04278_);
	assign _04280_ = _04060_ | _03525_;
	assign _04281_ = _00226_ & ~_04063_;
	assign _04282_ = _04280_ & ~_04281_;
	assign _04283_ = _03503_ & ~_04066_;
	assign _04284_ = _04282_ & ~_04283_;
	assign _04286_ = (_04070_ ? _05515_ : _04284_);
	assign _04287_ = _06393_ & ~_04072_;
	assign _04288_ = _05337_ & ~_04075_;
	assign _04289_ = _04288_ | _04287_;
	assign _04290_ = _05326_ & ~_04079_;
	assign _04291_ = _04290_ | _04289_;
	assign _04292_ = (_04082_ ? _05624_ : _04291_);
	assign _04293_ = _04292_ ^ _04286_;
	assign _04294_ = _04293_ ^ _04279_;
	assign _04295_ = _04294_ ^ _04272_;
	assign _04297_ = _04295_ ^ _04266_;
	assign _04298_ = _04297_ ^ _00226_;
	assign _04299_ = _04265_ & ~_04298_;
	assign _04300_ = _03657_ ^ _03228_;
	assign _04301_ = _04040_ | _03810_;
	assign _04302_ = _03832_ & ~_04042_;
	assign _04303_ = _04301_ & ~_04302_;
	assign _04304_ = _03876_ & ~_04045_;
	assign _04305_ = _04303_ & ~_04304_;
	assign _04306_ = (_04048_ ? _04241_ : _04305_);
	assign _04308_ = _04050_ | _03810_;
	assign _04309_ = _03239_ & ~_04052_;
	assign _04310_ = _04308_ & ~_04309_;
	assign _04311_ = _03228_ & ~_04055_;
	assign _04312_ = _04310_ & ~_04311_;
	assign _04313_ = (_04058_ ? _00996_ : _04312_);
	assign _04314_ = _04060_ | _03184_;
	assign _04315_ = _03173_ & ~_04063_;
	assign _04316_ = _04314_ & ~_04315_;
	assign _04317_ = _03162_ & ~_04066_;
	assign _04319_ = _04316_ & ~_04317_;
	assign _04320_ = (_04070_ ? _03667_ : _04319_);
	assign _04321_ = _03261_ & ~_04072_;
	assign _04322_ = _03206_ & ~_04075_;
	assign _04323_ = _04322_ | _04321_;
	assign _04324_ = _03162_ & ~_04079_;
	assign _04325_ = _04324_ | _04323_;
	assign _04326_ = (_04082_ ? \mchip.wrapper.keyReg.Q [7] : _04325_);
	assign _04327_ = _04326_ ^ _04320_;
	assign _04328_ = _04327_ ^ _04313_;
	assign _04330_ = _04328_ ^ _04306_;
	assign _04331_ = _04330_ ^ _04300_;
	assign _04332_ = _04331_ ^ _03239_;
	assign _04333_ = _03690_ ^ _03283_;
	assign _04334_ = _04040_ | _01835_;
	assign _04335_ = _03294_ & ~_04042_;
	assign _04336_ = _04334_ & ~_04335_;
	assign _04337_ = _03283_ & ~_04045_;
	assign _04338_ = _04336_ & ~_04337_;
	assign _04339_ = (_04048_ ? _04558_ : _04338_);
	assign _04341_ = _04050_ | _03305_;
	assign _04342_ = _03294_ & ~_04052_;
	assign _04343_ = _04341_ & ~_04342_;
	assign _04344_ = _03283_ & ~_04055_;
	assign _04345_ = _04343_ & ~_04344_;
	assign _04346_ = (_04058_ ? _04558_ : _04345_);
	assign _04347_ = _04060_ | _03305_;
	assign _04348_ = _04503_ & ~_04063_;
	assign _04349_ = _04347_ & ~_04348_;
	assign _04350_ = _03283_ & ~_04066_;
	assign _04352_ = _04349_ & ~_04350_;
	assign _04353_ = (_04070_ ? _04471_ : _04352_);
	assign _04354_ = _06308_ & ~_04072_;
	assign _04355_ = _03129_ & ~_04075_;
	assign _04356_ = _04355_ | _04354_;
	assign _04357_ = _03085_ & ~_04079_;
	assign _04358_ = _04357_ | _04356_;
	assign _04359_ = (_04082_ ? \mchip.wrapper.keyReg.Q [6] : _04358_);
	assign _04360_ = _04359_ ^ _04353_;
	assign _04361_ = _04360_ ^ _04346_;
	assign _04363_ = _04361_ ^ _04339_;
	assign _04364_ = _04363_ ^ _04333_;
	assign _04365_ = _04364_ ^ _03294_;
	assign _04366_ = ~(_04365_ & _04332_);
	assign _04367_ = _04299_ & ~_04366_;
	assign _04368_ = ~(_04298_ & _04265_);
	assign _04369_ = ~(_04368_ | _04366_);
	assign _04370_ = _04298_ | _04265_;
	assign _04371_ = ~(_04370_ | _04366_);
	assign _04372_ = ~_04371_;
	assign _04374_ = _04332_ | ~_04365_;
	assign _04375_ = _04374_ | ~_04299_;
	assign _04376_ = ~(_04374_ | _04370_);
	assign _04377_ = _04365_ | _04332_;
	assign _04378_ = _04377_ | _04370_;
	assign _04379_ = _04265_ | ~_04298_;
	assign _04380_ = ~(_04379_ | _04377_);
	assign _04381_ = ~(_04380_ & _04378_);
	assign _04382_ = ~(_04377_ | _04368_);
	assign _04383_ = _04381_ & ~_04382_;
	assign _04385_ = _04299_ & ~_04377_;
	assign _04386_ = _04385_ | ~_04383_;
	assign _04387_ = ~(_04379_ | _04374_);
	assign _04388_ = _04386_ & ~_04387_;
	assign _04389_ = _04388_ | _04376_;
	assign _04390_ = _04374_ | _04368_;
	assign _04391_ = _04390_ & ~_04389_;
	assign _04392_ = _04391_ & _04375_;
	assign _04393_ = _04365_ | ~_04332_;
	assign _04394_ = ~(_04393_ | _04379_);
	assign _04395_ = _04392_ & ~_04394_;
	assign _04396_ = ~(_04393_ | _04370_);
	assign _04397_ = _04395_ & ~_04396_;
	assign _04398_ = ~(_04393_ | _04368_);
	assign _04399_ = _04397_ & ~_04398_;
	assign _04400_ = _04299_ & ~_04393_;
	assign _04401_ = _04400_ | _04399_;
	assign _04402_ = _04379_ | _04366_;
	assign _04403_ = _04402_ & _04401_;
	assign _04404_ = _04372_ & ~_04403_;
	assign _04406_ = _04404_ | _04369_;
	assign _04407_ = _04406_ | _04367_;
	assign _04408_ = _04232_ & ~_04407_;
	assign _04409_ = _04408_ | _04231_;
	assign _04410_ = _04409_ | _04037_;
	assign _04411_ = _04410_ | _01973_;
	assign _04412_ = _04411_ | _03008_;
	assign _04413_ = _04232_ | _04038_;
	assign _04414_ = _03858_ | _01975_;
	assign _04415_ = _04414_ | _04413_;
	assign _04417_ = _01719_ | _03030_;
	assign _04418_ = _01938_ | _01898_;
	assign _04419_ = _04418_ | _04417_;
	assign _04420_ = _04419_ | _04415_;
	assign _04421_ = _00503_ | _06455_;
	assign _04422_ = _04421_ | _04811_;
	assign _04423_ = _01537_ | _01053_;
	assign _04424_ = _02502_ | _02028_;
	assign _04425_ = _04424_ | _04423_;
	assign _04426_ = _04425_ | _04422_;
	assign _04428_ = _04426_ | _04420_;
	assign _04429_ = \mchip.wrapper.intxtReg.Q [1] & ~\mchip.wrapper.intxtReg.Q [0];
	assign _04430_ = \mchip.wrapper.intxtReg.Q [3] | ~\mchip.wrapper.intxtReg.Q [2];
	assign _04431_ = _04429_ & ~_04430_;
	assign _04432_ = ~_04431_;
	assign _04433_ = \mchip.wrapper.intxtReg.Q [1] | ~\mchip.wrapper.intxtReg.Q [0];
	assign _04434_ = ~(_04433_ | _04430_);
	assign _04435_ = \mchip.wrapper.intxtReg.Q [2] | \mchip.wrapper.intxtReg.Q [3];
	assign _04436_ = ~(_04435_ | _04433_);
	assign _04437_ = \mchip.wrapper.intxtReg.Q [1] | \mchip.wrapper.intxtReg.Q [0];
	assign _04439_ = ~(_04437_ | _04435_);
	assign _04440_ = _04436_ | ~_04439_;
	assign _04441_ = _04429_ & ~_04435_;
	assign _04442_ = _04440_ & ~_04441_;
	assign _04443_ = ~(\mchip.wrapper.intxtReg.Q [1] & \mchip.wrapper.intxtReg.Q [0]);
	assign _04444_ = ~(_04443_ | _04435_);
	assign _04445_ = _04444_ | ~_04442_;
	assign _04446_ = ~(_04437_ | _04430_);
	assign _04447_ = _04445_ & ~_04446_;
	assign _04448_ = _04447_ | _04434_;
	assign _04450_ = _04432_ & ~_04448_;
	assign _04451_ = ~(_04443_ | _04430_);
	assign _04452_ = _04450_ & ~_04451_;
	assign _04453_ = \mchip.wrapper.intxtReg.Q [2] | ~\mchip.wrapper.intxtReg.Q [3];
	assign _04454_ = ~(_04453_ | _04437_);
	assign _04455_ = _04452_ & ~_04454_;
	assign _04456_ = ~(_04453_ | _04433_);
	assign _04457_ = _04455_ & ~_04456_;
	assign _04458_ = _04429_ & ~_04453_;
	assign _04459_ = _04457_ & ~_04458_;
	assign _04461_ = ~(_04453_ | _04443_);
	assign _04462_ = _04461_ | _04459_;
	assign _04463_ = ~(\mchip.wrapper.intxtReg.Q [2] & \mchip.wrapper.intxtReg.Q [3]);
	assign _04464_ = ~(_04463_ | _04437_);
	assign _04465_ = ~_04464_;
	assign _04466_ = _04465_ & _04462_;
	assign _04467_ = ~(_04463_ | _04433_);
	assign _04468_ = _04467_ | _04466_;
	assign _04469_ = _04429_ & ~_04463_;
	assign _04470_ = _04468_ & ~_04469_;
	assign _04472_ = ~(_04463_ | _04443_);
	assign _04473_ = _04470_ & ~_04472_;
	assign io_out[0] = (_04428_ ? _04412_ : _04473_);
	assign _04474_ = ~_05141_;
	assign _04475_ = ~_06302_;
	assign _04476_ = ~(\mchip.wrapper.intxtReg.Q [7] | \mchip.wrapper.intxtReg.Q [6]);
	assign _04477_ = ~(_04476_ | _06207_);
	assign _04478_ = _04477_ | _06101_;
	assign _04479_ = _06022_ & ~_04478_;
	assign _04480_ = _04479_ | _06250_;
	assign _04482_ = _04480_ | _06281_;
	assign _04483_ = _04475_ & ~_04482_;
	assign _04484_ = _04483_ & ~_06324_;
	assign _04485_ = _04484_ | _06346_;
	assign _04486_ = _06379_ & ~_04485_;
	assign _04487_ = _05691_ & ~_04486_;
	assign _04488_ = _04487_ | _05360_;
	assign _04489_ = _04474_ & ~_04488_;
	assign _04490_ = _04811_ & ~_04489_;
	assign _04491_ = ~_00021_;
	assign _04493_ = ~_00350_;
	assign _04494_ = \mchip.wrapper.intxtReg.Q [10] | \mchip.wrapper.intxtReg.Q [11];
	assign _04495_ = _04494_ & ~_00252_;
	assign _04496_ = _04495_ | _00120_;
	assign _04497_ = _00109_ & ~_04496_;
	assign _04498_ = _04497_ | _00296_;
	assign _04499_ = _04498_ | _00329_;
	assign _04500_ = _04493_ & ~_04499_;
	assign _04501_ = _04500_ & ~_00372_;
	assign _04502_ = _04501_ | _00394_;
	assign _04504_ = _00426_ & ~_04502_;
	assign _04505_ = _00076_ & ~_04504_;
	assign _04506_ = _04505_ | _00043_;
	assign _04507_ = _04491_ & ~_04506_;
	assign _04508_ = _06455_ & ~_04507_;
	assign _04509_ = ~_00536_;
	assign _04510_ = ~_00866_;
	assign _04511_ = \mchip.wrapper.intxtReg.Q [14] | \mchip.wrapper.intxtReg.Q [15];
	assign _04512_ = _04511_ & ~_00767_;
	assign _04513_ = _04512_ | _00635_;
	assign _04515_ = _00624_ & ~_04513_;
	assign _04516_ = _04515_ | _00811_;
	assign _04517_ = _04516_ | _00844_;
	assign _04518_ = _04510_ & ~_04517_;
	assign _04519_ = _04518_ & ~_00888_;
	assign _04520_ = _04519_ | _00910_;
	assign _04521_ = _00943_ & ~_04520_;
	assign _04522_ = _00591_ & ~_04521_;
	assign _04523_ = _04522_ | _00558_;
	assign _04524_ = _04509_ & ~_04523_;
	assign _04526_ = _00503_ & ~_04524_;
	assign _04527_ = _04526_ | _04508_;
	assign _04528_ = _04527_ | _04490_;
	assign _04529_ = ~_01086_;
	assign _04530_ = ~_01394_;
	assign _04531_ = ~(\mchip.wrapper.keyReg.Q [3] | \mchip.wrapper.keyReg.Q [2]);
	assign _04532_ = ~(_04531_ | _01295_);
	assign _04533_ = _04532_ | _01185_;
	assign _04534_ = _01174_ & ~_04533_;
	assign _04535_ = _04534_ | _01339_;
	assign _04537_ = _04535_ | _01372_;
	assign _04538_ = _04530_ & ~_04537_;
	assign _04539_ = _04538_ & ~_01416_;
	assign _04540_ = _04539_ | _01438_;
	assign _04541_ = _01471_ & ~_04540_;
	assign _04542_ = _01141_ & ~_04541_;
	assign _04543_ = _04542_ | _01108_;
	assign _04544_ = _04529_ & ~_04543_;
	assign _04545_ = _01053_ & ~_04544_;
	assign _04546_ = ~_01570_;
	assign _04548_ = ~_01877_;
	assign _04549_ = ~_01734_;
	assign _04550_ = ~(_01712_ | _01690_);
	assign _04551_ = ~(_04550_ & _04549_);
	assign _04552_ = _04551_ | _01756_;
	assign _04553_ = ~(_04552_ | _01778_);
	assign _04554_ = _04553_ | _01668_;
	assign _04555_ = _01657_ & ~_04554_;
	assign _04556_ = _04555_ | _01822_;
	assign _04557_ = _04556_ | _01855_;
	assign _04559_ = _04548_ & ~_04557_;
	assign _04560_ = _04559_ & ~_01899_;
	assign _04561_ = _04560_ | _01921_;
	assign _04562_ = _01954_ & ~_04561_;
	assign _04563_ = _01625_ & ~_04562_;
	assign _04564_ = _04563_ | _01592_;
	assign _04565_ = _04546_ & ~_04564_;
	assign _04566_ = _01537_ & ~_04565_;
	assign _04567_ = _04566_ | _04545_;
	assign _04568_ = ~_02059_;
	assign _04570_ = ~_02359_;
	assign _04571_ = ~(\mchip.wrapper.keyReg.Q [11] | \mchip.wrapper.keyReg.Q [10]);
	assign _04572_ = ~(_04571_ | _02260_);
	assign _04573_ = _04572_ | _02152_;
	assign _04574_ = _02141_ & ~_04573_;
	assign _04575_ = _04574_ | _02304_;
	assign _04576_ = _04575_ | _02337_;
	assign _04577_ = _04570_ & ~_04576_;
	assign _04578_ = _04577_ & ~_02381_;
	assign _04579_ = _04578_ | _02403_;
	assign _04580_ = _02436_ & ~_04579_;
	assign _04581_ = _02110_ & ~_04580_;
	assign _04582_ = _04581_ | _02079_;
	assign _04583_ = _04568_ & ~_04582_;
	assign _04584_ = _02028_ & ~_04583_;
	assign _04585_ = ~_02535_;
	assign _04586_ = ~_02843_;
	assign _04587_ = ~_02700_;
	assign _04588_ = ~(_02678_ | _02656_);
	assign _04589_ = ~(_04588_ & _04587_);
	assign _04592_ = _04589_ | _02722_;
	assign _04593_ = ~(_04592_ | _02744_);
	assign _04594_ = _04593_ | _02634_;
	assign _04595_ = _02623_ & ~_04594_;
	assign _04596_ = _04595_ | _02788_;
	assign _04597_ = _04596_ | _02821_;
	assign _04598_ = _04586_ & ~_04597_;
	assign _04599_ = _04598_ & ~_02865_;
	assign _04600_ = _04599_ | _02887_;
	assign _04601_ = _02920_ & ~_04600_;
	assign _04603_ = _02590_ & ~_04601_;
	assign _04604_ = _04603_ | _02557_;
	assign _04605_ = _04585_ & ~_04604_;
	assign _04606_ = _02502_ & ~_04605_;
	assign _04607_ = _04606_ | _04584_;
	assign _04608_ = _04607_ | _04567_;
	assign _04609_ = _04608_ | _04528_;
	assign _04610_ = _01689_ | _01688_;
	assign _04611_ = _04610_ | _01692_;
	assign _04612_ = _04611_ | _01694_;
	assign _04614_ = ~(_04612_ | _01696_);
	assign _04615_ = _04614_ | _01685_;
	assign _04616_ = _01699_ & ~_04615_;
	assign _04617_ = _04616_ | ~_01684_;
	assign _04618_ = _04617_ | _01704_;
	assign _04619_ = _04618_ | _01706_;
	assign _04620_ = ~(_04619_ | _01708_);
	assign _04621_ = _04620_ | _01710_;
	assign _04622_ = _01713_ & ~_04621_;
	assign _04623_ = _01682_ & ~_04622_;
	assign _04625_ = _04623_ | _01680_;
	assign _04626_ = ~(_04625_ | _01677_);
	assign _04627_ = _03030_ & ~_04626_;
	assign _04628_ = _01868_ | _01867_;
	assign _04629_ = _04628_ | _01870_;
	assign _04630_ = _04629_ | _01872_;
	assign _04631_ = ~(_04630_ | _01874_);
	assign _04632_ = _04631_ | _01863_;
	assign _04633_ = _01878_ & ~_04632_;
	assign _04634_ = _04633_ | ~_01862_;
	assign _04636_ = _04634_ | _01882_;
	assign _04637_ = _04636_ | _01884_;
	assign _04638_ = ~(_04637_ | _01886_);
	assign _04639_ = _04638_ | _01889_;
	assign _04640_ = _01891_ & ~_04639_;
	assign _04641_ = _01860_ & ~_04640_;
	assign _04642_ = _04641_ | _01858_;
	assign _04643_ = ~(_04642_ | _01856_);
	assign _04644_ = _01719_ & ~_04643_;
	assign _04645_ = _04644_ | _04627_;
	assign _04647_ = ~_01900_;
	assign _04648_ = ~_01911_;
	assign _04649_ = ~(_01908_ | _01906_);
	assign _04650_ = ~(_04649_ & _04648_);
	assign _04651_ = _04650_ | _01913_;
	assign _04652_ = ~(_04651_ | _01915_);
	assign _04653_ = _04652_ | _01905_;
	assign _04654_ = _01904_ & ~_04653_;
	assign _04655_ = _04654_ | _01919_;
	assign _04656_ = _04655_ | _01922_;
	assign _04658_ = ~(_04656_ | _01924_);
	assign _04659_ = _04658_ & ~_01926_;
	assign _04660_ = _04659_ | _01928_;
	assign _04661_ = _01931_ & ~_04660_;
	assign _04662_ = _01903_ & ~_04661_;
	assign _04663_ = _04662_ | _01901_;
	assign _04664_ = _04647_ & ~_04663_;
	assign _04665_ = _01898_ & ~_04664_;
	assign _04666_ = ~(_01340_ | _01950_);
	assign _04668_ = _04666_ | _01946_;
	assign _04669_ = _01945_ & ~_04668_;
	assign _04670_ = _04669_ | _01955_;
	assign _04671_ = _04670_ | _01957_;
	assign _04672_ = _04671_ | _01959_;
	assign _04673_ = ~(_04672_ | _01961_);
	assign _04674_ = _04673_ | _01963_;
	assign _04675_ = _01966_ & ~_04674_;
	assign _04676_ = _01942_ & ~_04675_;
	assign _04677_ = _04676_ | _01940_;
	assign _04679_ = ~(_04677_ | _01939_);
	assign _04680_ = _01938_ & ~_04679_;
	assign _04681_ = _04680_ | _04665_;
	assign _04682_ = _04681_ | _04645_;
	assign _04683_ = ~_03814_;
	assign _04684_ = ~_03829_;
	assign _04685_ = ~(_03827_ | _03825_);
	assign _04686_ = ~(_04685_ & _04684_);
	assign _04687_ = _04686_ | _03831_;
	assign _04688_ = ~(_04687_ | _03834_);
	assign _04690_ = _04688_ | _03823_;
	assign _04691_ = _03822_ & ~_04690_;
	assign _04692_ = _04691_ | _03838_;
	assign _04693_ = _04692_ | _03841_;
	assign _04694_ = _04693_ | _03844_;
	assign _04695_ = ~(_04694_ | _03846_);
	assign _04696_ = _04695_ | _03848_;
	assign _04697_ = _03851_ & ~_04696_;
	assign _04698_ = _03819_ & ~_04697_;
	assign _04699_ = _04698_ | _03816_;
	assign _04702_ = _04683_ & ~_04699_;
	assign _04703_ = _01975_ & ~_04702_;
	assign _04704_ = ~_03995_;
	assign _04705_ = ~_04009_;
	assign _04706_ = ~(_04007_ | _04005_);
	assign _04707_ = ~(_04706_ & _04705_);
	assign _04708_ = _04707_ | _04011_;
	assign _04709_ = ~(_04708_ | _04013_);
	assign _04710_ = _04709_ | _04003_;
	assign _04711_ = _04002_ & ~_04710_;
	assign _04713_ = _04711_ | _04018_;
	assign _04714_ = _04713_ | _04021_;
	assign _04715_ = _04714_ | _04023_;
	assign _04716_ = ~(_04715_ | _04025_);
	assign _04717_ = _04716_ | _04028_;
	assign _04718_ = _04031_ & ~_04717_;
	assign _04719_ = _04000_ & ~_04718_;
	assign _04720_ = _04719_ | _03997_;
	assign _04721_ = _04704_ & ~_04720_;
	assign _04722_ = _03858_ & ~_04721_;
	assign _04724_ = _04722_ | _04703_;
	assign _04725_ = ~_04190_;
	assign _04726_ = ~_04205_;
	assign _04727_ = _04201_ & ~_04203_;
	assign _04728_ = ~(_04727_ & _04726_);
	assign _04729_ = _04728_ | _04207_;
	assign _04730_ = ~(_04729_ | _04210_);
	assign _04731_ = _04730_ | _04199_;
	assign _04732_ = _04213_ & ~_04731_;
	assign _04733_ = _04732_ | ~_04197_;
	assign _04735_ = _04733_ | _04217_;
	assign _04736_ = _04735_ | _04219_;
	assign _04737_ = ~(_04736_ | _04221_);
	assign _04738_ = _04737_ | _04223_;
	assign _04739_ = _04225_ & ~_04738_;
	assign _04740_ = _04195_ & ~_04739_;
	assign _04741_ = _04740_ | _04192_;
	assign _04742_ = _04725_ & ~_04741_;
	assign _04743_ = _04038_ & ~_04742_;
	assign _04744_ = ~_04367_;
	assign _04746_ = ~_04382_;
	assign _04747_ = _04378_ & ~_04380_;
	assign _04748_ = ~(_04747_ & _04746_);
	assign _04749_ = _04748_ | _04385_;
	assign _04750_ = ~(_04749_ | _04387_);
	assign _04751_ = _04750_ | _04376_;
	assign _04752_ = _04390_ & ~_04751_;
	assign _04753_ = _04752_ | ~_04375_;
	assign _04754_ = _04753_ | _04394_;
	assign _04755_ = _04754_ | _04396_;
	assign _04757_ = ~(_04755_ | _04398_);
	assign _04758_ = _04757_ | _04400_;
	assign _04759_ = _04402_ & ~_04758_;
	assign _04760_ = _04372_ & ~_04759_;
	assign _04761_ = _04760_ | _04369_;
	assign _04762_ = _04744_ & ~_04761_;
	assign _04763_ = _04232_ & ~_04762_;
	assign _04764_ = _04763_ | _04743_;
	assign _04765_ = _04764_ | _04724_;
	assign _04766_ = _04765_ | _04682_;
	assign _04768_ = _04766_ | _04609_;
	assign _04769_ = ~_04467_;
	assign _04770_ = ~_04456_;
	assign _04771_ = ~_04441_;
	assign _04772_ = ~(_04439_ | _04436_);
	assign _04773_ = ~(_04772_ & _04771_);
	assign _04774_ = ~(_04773_ | _04444_);
	assign _04775_ = _04774_ & ~_04446_;
	assign _04776_ = _04775_ | _04434_;
	assign _04777_ = _04432_ & ~_04776_;
	assign _04779_ = _04777_ | _04451_;
	assign _04780_ = _04779_ | _04454_;
	assign _04781_ = _04770_ & ~_04780_;
	assign _04782_ = _04781_ & ~_04458_;
	assign _04783_ = _04782_ | _04461_;
	assign _04784_ = _04465_ & ~_04783_;
	assign _04785_ = _04769_ & ~_04784_;
	assign _04786_ = _04785_ | _04469_;
	assign _04787_ = _04786_ | _04472_;
	assign io_out[1] = (_04428_ ? _04768_ : _04787_);
	assign _04789_ = ~_06346_;
	assign _04790_ = ~(_06143_ & _06121_);
	assign _04791_ = _04790_ & ~_06164_;
	assign _04792_ = _04791_ | _06185_;
	assign _04793_ = _04792_ | _06207_;
	assign _04794_ = _04793_ | _06101_;
	assign _04795_ = _04794_ | _05912_;
	assign _04796_ = _04795_ | _06250_;
	assign _04797_ = _04796_ | _06281_;
	assign _04798_ = _04797_ | _06302_;
	assign _04800_ = _04798_ | _06324_;
	assign _04801_ = _04789_ & ~_04800_;
	assign _04802_ = _06379_ & ~_04801_;
	assign _04803_ = _05691_ & ~_04802_;
	assign _04804_ = _04803_ | _05360_;
	assign _04805_ = _04474_ & ~_04804_;
	assign _04806_ = _04811_ & ~_04805_;
	assign _04807_ = ~_00394_;
	assign _04808_ = ~(_00164_ | _00142_);
	assign _04809_ = _00197_ & ~_04808_;
	assign _04812_ = _04809_ | _00219_;
	assign _04813_ = _04812_ | _00252_;
	assign _04814_ = _04813_ | _00120_;
	assign _04815_ = _04814_ | _00098_;
	assign _04816_ = _04815_ | _00296_;
	assign _04817_ = _04816_ | _00329_;
	assign _04818_ = _04817_ | _00350_;
	assign _04819_ = _04818_ | _00372_;
	assign _04820_ = _04807_ & ~_04819_;
	assign _04821_ = _00426_ & ~_04820_;
	assign _04823_ = _00076_ & ~_04821_;
	assign _04824_ = _04823_ | _00043_;
	assign _04825_ = _04491_ & ~_04824_;
	assign _04826_ = _06455_ & ~_04825_;
	assign _04827_ = ~_00910_;
	assign _04828_ = ~(_00679_ | _00657_);
	assign _04829_ = _00712_ & ~_04828_;
	assign _04830_ = _04829_ | _00734_;
	assign _04831_ = _04830_ | _00767_;
	assign _04832_ = _04831_ | _00635_;
	assign _04834_ = _04832_ | _00613_;
	assign _04835_ = _04834_ | _00811_;
	assign _04836_ = _04835_ | _00844_;
	assign _04837_ = _04836_ | _00866_;
	assign _04838_ = _04837_ | _00888_;
	assign _04839_ = _04827_ & ~_04838_;
	assign _04840_ = _00943_ & ~_04839_;
	assign _04841_ = _00591_ & ~_04840_;
	assign _04842_ = _04841_ | _00558_;
	assign _04843_ = _04509_ & ~_04842_;
	assign _04845_ = _00503_ & ~_04843_;
	assign _04846_ = _04845_ | _04826_;
	assign _04847_ = _04846_ | _04806_;
	assign _04848_ = ~_01438_;
	assign _04849_ = ~(_01229_ & _01207_);
	assign _04850_ = _04849_ & ~_01251_;
	assign _04851_ = _04850_ | _01273_;
	assign _04852_ = _04851_ | _01295_;
	assign _04853_ = _04852_ | _01185_;
	assign _04854_ = _04853_ | _01163_;
	assign _04856_ = _04854_ | _01339_;
	assign _04857_ = _04856_ | _01372_;
	assign _04858_ = _04857_ | _01394_;
	assign _04859_ = _04858_ | _01416_;
	assign _04860_ = _04848_ & ~_04859_;
	assign _04861_ = _01471_ & ~_04860_;
	assign _04862_ = _01141_ & ~_04861_;
	assign _04863_ = _04862_ | _01108_;
	assign _04864_ = _04529_ & ~_04863_;
	assign _04865_ = _01053_ & ~_04864_;
	assign _04867_ = ~_01921_;
	assign _04868_ = _04549_ & ~_04550_;
	assign _04869_ = _04868_ | _01756_;
	assign _04870_ = _04869_ | _01778_;
	assign _04871_ = _04870_ | _01668_;
	assign _04872_ = _04871_ | _01647_;
	assign _04873_ = _04872_ | _01822_;
	assign _04874_ = _04873_ | _01855_;
	assign _04875_ = _04874_ | _01877_;
	assign _04876_ = _04875_ | _01899_;
	assign _04878_ = _04867_ & ~_04876_;
	assign _04879_ = _01954_ & ~_04878_;
	assign _04880_ = _01625_ & ~_04879_;
	assign _04881_ = _04880_ | _01592_;
	assign _04882_ = _04546_ & ~_04881_;
	assign _04883_ = _01537_ & ~_04882_;
	assign _04884_ = _04883_ | _04865_;
	assign _04885_ = ~_02403_;
	assign _04886_ = ~(_02196_ & _02174_);
	assign _04887_ = _04886_ & ~_02216_;
	assign _04889_ = _04887_ | _02238_;
	assign _04890_ = _04889_ | _02260_;
	assign _04891_ = _04890_ | _02152_;
	assign _04892_ = _04891_ | _02130_;
	assign _04893_ = _04892_ | _02304_;
	assign _04894_ = _04893_ | _02337_;
	assign _04895_ = _04894_ | _02359_;
	assign _04896_ = _04895_ | _02381_;
	assign _04897_ = _04885_ & ~_04896_;
	assign _04898_ = _02436_ & ~_04897_;
	assign _04900_ = _02110_ & ~_04898_;
	assign _04901_ = _04900_ | _02079_;
	assign _04902_ = _04568_ & ~_04901_;
	assign _04903_ = _02028_ & ~_04902_;
	assign _04904_ = ~_02887_;
	assign _04905_ = _04587_ & ~_04588_;
	assign _04906_ = _04905_ | _02722_;
	assign _04907_ = _04906_ | _02744_;
	assign _04908_ = _04907_ | _02634_;
	assign _04909_ = _04908_ | _02612_;
	assign _04911_ = _04909_ | _02788_;
	assign _04912_ = _04911_ | _02821_;
	assign _04913_ = _04912_ | _02843_;
	assign _04914_ = _04913_ | _02865_;
	assign _04915_ = _04904_ & ~_04914_;
	assign _04916_ = _02920_ & ~_04915_;
	assign _04917_ = _02590_ & ~_04916_;
	assign _04918_ = _04917_ | _02557_;
	assign _04919_ = _04585_ & ~_04918_;
	assign _04920_ = _02502_ & ~_04919_;
	assign _04923_ = _04920_ | _04903_;
	assign _04924_ = _04923_ | _04884_;
	assign _04925_ = _04924_ | _04847_;
	assign _04926_ = _04610_ & ~_01692_;
	assign _04927_ = _04926_ | _01694_;
	assign _04928_ = _04927_ | _01696_;
	assign _04929_ = _04928_ | _01685_;
	assign _04930_ = _04929_ | ~_01699_;
	assign _04931_ = _04930_ | ~_01684_;
	assign _04932_ = _04931_ | _01704_;
	assign _04934_ = _04932_ | _01706_;
	assign _04935_ = _04934_ | _01708_;
	assign _04936_ = ~(_04935_ | _01710_);
	assign _04937_ = _01713_ & ~_04936_;
	assign _04938_ = _01682_ & ~_04937_;
	assign _04939_ = _04938_ | _01680_;
	assign _04940_ = ~(_04939_ | _01677_);
	assign _04941_ = _03030_ & ~_04940_;
	assign _04942_ = _04628_ & ~_01870_;
	assign _04943_ = _04942_ | _01872_;
	assign _04945_ = _04943_ | _01874_;
	assign _04946_ = _04945_ | _01863_;
	assign _04947_ = _04946_ | ~_01878_;
	assign _04948_ = _04947_ | ~_01862_;
	assign _04949_ = _04948_ | _01882_;
	assign _04950_ = _04949_ | _01884_;
	assign _04951_ = _04950_ | _01886_;
	assign _04952_ = ~(_04951_ | _01889_);
	assign _04953_ = _01891_ & ~_04952_;
	assign _04954_ = _01860_ & ~_04953_;
	assign _04956_ = _04954_ | _01858_;
	assign _04957_ = ~(_04956_ | _01856_);
	assign _04958_ = _01719_ & ~_04957_;
	assign _04959_ = _04958_ | _04941_;
	assign _04960_ = ~_01928_;
	assign _04961_ = _04648_ & ~_04649_;
	assign _04962_ = _04961_ | _01913_;
	assign _04963_ = _04962_ | _01915_;
	assign _04964_ = _04963_ | _01905_;
	assign _04965_ = _04964_ | ~_01904_;
	assign _04967_ = _04965_ | _01919_;
	assign _04968_ = _04967_ | _01922_;
	assign _04969_ = _04968_ | _01924_;
	assign _04970_ = _04969_ | _01926_;
	assign _04971_ = _04960_ & ~_04970_;
	assign _04972_ = _01931_ & ~_04971_;
	assign _04973_ = _01903_ & ~_04972_;
	assign _04974_ = _04973_ | _01901_;
	assign _04975_ = _04647_ & ~_04974_;
	assign _04976_ = _01898_ & ~_04975_;
	assign _04978_ = ~_01963_;
	assign _04979_ = _01340_ & ~_01410_;
	assign _04980_ = _01340_ & ~_01413_;
	assign _04981_ = _01417_ & _01340_;
	assign _04982_ = ~(_04981_ | _04980_);
	assign _04983_ = ~(_04982_ | _04979_);
	assign _04984_ = _04983_ | _01948_;
	assign _04985_ = _04984_ | _01950_;
	assign _04986_ = _04985_ | _01946_;
	assign _04987_ = _04986_ | _01944_;
	assign _04989_ = _04987_ | _01955_;
	assign _04990_ = _04989_ | _01957_;
	assign _04991_ = _04990_ | _01959_;
	assign _04992_ = _04991_ | _01961_;
	assign _04993_ = _04978_ & ~_04992_;
	assign _04994_ = _01966_ & ~_04993_;
	assign _04995_ = _01942_ & ~_04994_;
	assign _04996_ = ~(_04995_ | _01940_);
	assign _04997_ = _04996_ & ~_01939_;
	assign _04998_ = _01938_ & ~_04997_;
	assign _05000_ = _04998_ | _04976_;
	assign _05001_ = _05000_ | _04959_;
	assign _05002_ = _04684_ & ~_04685_;
	assign _05003_ = _05002_ | _03831_;
	assign _05004_ = _05003_ | _03834_;
	assign _05005_ = _05004_ | _03823_;
	assign _05006_ = _05005_ | ~_03822_;
	assign _05007_ = _05006_ | _03838_;
	assign _05008_ = _05007_ | _03841_;
	assign _05009_ = _05008_ | _03844_;
	assign _05011_ = _05009_ | _03846_;
	assign _05012_ = ~(_05011_ | _03848_);
	assign _05013_ = _03851_ & ~_05012_;
	assign _05014_ = _03819_ & ~_05013_;
	assign _05015_ = _05014_ | _03816_;
	assign _05016_ = _04683_ & ~_05015_;
	assign _05017_ = _01975_ & ~_05016_;
	assign _05018_ = _04705_ & ~_04706_;
	assign _05019_ = _05018_ | _04011_;
	assign _05020_ = _05019_ | _04013_;
	assign _05022_ = _05020_ | _04003_;
	assign _05023_ = _05022_ | ~_04002_;
	assign _05024_ = _05023_ | _04018_;
	assign _05025_ = _05024_ | _04021_;
	assign _05026_ = _05025_ | _04023_;
	assign _05027_ = _05026_ | _04025_;
	assign _05028_ = ~(_05027_ | _04028_);
	assign _05029_ = _04031_ & ~_05028_;
	assign _05030_ = _04000_ & ~_05029_;
	assign _05031_ = _05030_ | _03997_;
	assign _05034_ = _04704_ & ~_05031_;
	assign _05035_ = _03858_ & ~_05034_;
	assign _05036_ = _05035_ | _05017_;
	assign _05037_ = _04726_ & ~_04727_;
	assign _05038_ = _05037_ | _04207_;
	assign _05039_ = _05038_ | _04210_;
	assign _05040_ = _05039_ | _04199_;
	assign _05041_ = _05040_ | ~_04213_;
	assign _05042_ = _05041_ | ~_04197_;
	assign _05043_ = _05042_ | _04217_;
	assign _05045_ = _05043_ | _04219_;
	assign _05046_ = _05045_ | _04221_;
	assign _05047_ = ~(_05046_ | _04223_);
	assign _05048_ = _04225_ & ~_05047_;
	assign _05049_ = _04195_ & ~_05048_;
	assign _05050_ = _05049_ | _04192_;
	assign _05051_ = _04725_ & ~_05050_;
	assign _05052_ = _04038_ & ~_05051_;
	assign _05053_ = _04746_ & ~_04747_;
	assign _05054_ = _05053_ | _04385_;
	assign _05055_ = _05054_ | _04387_;
	assign _05056_ = _05055_ | _04376_;
	assign _05057_ = _05056_ | ~_04390_;
	assign _05058_ = _05057_ | ~_04375_;
	assign _05059_ = _05058_ | _04394_;
	assign _05060_ = _05059_ | _04396_;
	assign _05061_ = _05060_ | _04398_;
	assign _05062_ = ~(_05061_ | _04400_);
	assign _05063_ = _04402_ & ~_05062_;
	assign _05064_ = _04372_ & ~_05063_;
	assign _05065_ = _05064_ | _04369_;
	assign _05066_ = _04744_ & ~_05065_;
	assign _05067_ = _04232_ & ~_05066_;
	assign _05068_ = _05067_ | _05052_;
	assign _05069_ = _05068_ | _05036_;
	assign _05070_ = _05069_ | _05001_;
	assign _05071_ = _05070_ | _04925_;
	assign _05072_ = ~_04461_;
	assign _05073_ = _04771_ & ~_04772_;
	assign _05074_ = _05073_ | _04444_;
	assign _05076_ = _05074_ | _04446_;
	assign _05077_ = _05076_ | _04434_;
	assign _05078_ = _05077_ | _04431_;
	assign _05079_ = _05078_ | _04451_;
	assign _05080_ = _05079_ | _04454_;
	assign _05081_ = _05080_ | _04456_;
	assign _05082_ = _05081_ | _04458_;
	assign _05083_ = _05072_ & ~_05082_;
	assign _05084_ = _04465_ & ~_05083_;
	assign _05085_ = _04769_ & ~_05084_;
	assign _05087_ = _05085_ | _04469_;
	assign _05088_ = _05087_ | _04472_;
	assign io_out[2] = (_04428_ ? _05071_ : _05088_);
	assign _05089_ = ~_06250_;
	assign _05090_ = _05089_ & ~_06239_;
	assign _05091_ = _05090_ | _06281_;
	assign _05092_ = ~(_05091_ | _06302_);
	assign _05093_ = ~(_05092_ | _06324_);
	assign _05094_ = _05093_ | _06346_;
	assign _05095_ = _05094_ | ~_06379_;
	assign _05097_ = _05095_ | ~_05691_;
	assign _05098_ = ~(_05097_ | _05360_);
	assign _05099_ = ~(_05098_ | _05141_);
	assign _05100_ = _04811_ & ~_05099_;
	assign _05101_ = ~_00296_;
	assign _05102_ = _05101_ & ~_00285_;
	assign _05103_ = _05102_ | _00329_;
	assign _05104_ = ~(_05103_ | _00350_);
	assign _05105_ = ~(_05104_ | _00372_);
	assign _05106_ = _05105_ | _00394_;
	assign _05108_ = _05106_ | ~_00426_;
	assign _05109_ = _05108_ | ~_00076_;
	assign _05110_ = ~(_05109_ | _00043_);
	assign _05111_ = _04491_ & ~_05110_;
	assign _05112_ = _06455_ & ~_05111_;
	assign _05113_ = ~_00811_;
	assign _05114_ = _05113_ & ~_00800_;
	assign _05115_ = _05114_ | _00844_;
	assign _05116_ = ~(_05115_ | _00866_);
	assign _05117_ = ~(_05116_ | _00888_);
	assign _05119_ = _05117_ | _00910_;
	assign _05120_ = _05119_ | ~_00943_;
	assign _05121_ = _05120_ | ~_00591_;
	assign _05122_ = ~(_05121_ | _00558_);
	assign _05123_ = _04509_ & ~_05122_;
	assign _05124_ = _00503_ & ~_05123_;
	assign _05125_ = _05124_ | _05112_;
	assign _05126_ = _05125_ | _05100_;
	assign _05127_ = ~_01339_;
	assign _05128_ = _05127_ & ~_01328_;
	assign _05130_ = _05128_ | _01372_;
	assign _05131_ = ~(_05130_ | _01394_);
	assign _05132_ = ~(_05131_ | _01416_);
	assign _05133_ = _05132_ | _01438_;
	assign _05134_ = _05133_ | ~_01471_;
	assign _05135_ = _05134_ | ~_01141_;
	assign _05136_ = ~(_05135_ | _01108_);
	assign _05137_ = ~(_05136_ | _01086_);
	assign _05138_ = _01053_ & ~_05137_;
	assign _05139_ = ~_01822_;
	assign _05142_ = _05139_ & ~_01811_;
	assign _05143_ = _05142_ | _01855_;
	assign _05144_ = ~(_05143_ | _01877_);
	assign _05145_ = ~(_05144_ | _01899_);
	assign _05146_ = _05145_ | _01921_;
	assign _05147_ = _05146_ | ~_01954_;
	assign _05148_ = _05147_ | ~_01625_;
	assign _05149_ = ~(_05148_ | _01592_);
	assign _05150_ = ~(_05149_ | _01570_);
	assign _05151_ = _01537_ & ~_05150_;
	assign _05153_ = _05151_ | _05138_;
	assign _05154_ = ~_02304_;
	assign _05155_ = _05154_ & ~_02293_;
	assign _05156_ = _05155_ | _02337_;
	assign _05157_ = ~(_05156_ | _02359_);
	assign _05158_ = ~(_05157_ | _02381_);
	assign _05159_ = _05158_ | _02403_;
	assign _05160_ = _05159_ | ~_02436_;
	assign _05161_ = _05160_ | ~_02110_;
	assign _05162_ = ~(_05161_ | _02079_);
	assign _05164_ = ~(_05162_ | _02059_);
	assign _05165_ = _02028_ & ~_05164_;
	assign _05166_ = ~_02788_;
	assign _05167_ = _05166_ & ~_02777_;
	assign _05168_ = _05167_ | _02821_;
	assign _05169_ = ~(_05168_ | _02843_);
	assign _05170_ = ~(_05169_ | _02865_);
	assign _05171_ = _05170_ | _02887_;
	assign _05172_ = _05171_ | ~_02920_;
	assign _05173_ = _05172_ | ~_02590_;
	assign _05175_ = ~(_05173_ | _02557_);
	assign _05176_ = ~(_05175_ | _02535_);
	assign _05177_ = _02502_ & ~_05176_;
	assign _05178_ = _05177_ | _05165_;
	assign _05179_ = _05178_ | _05153_;
	assign _05180_ = _05179_ | _05126_;
	assign _05181_ = _01684_ & ~_01700_;
	assign _05182_ = _05181_ | _01704_;
	assign _05183_ = ~(_05182_ | _01706_);
	assign _05184_ = ~(_05183_ | _01708_);
	assign _05186_ = _05184_ | _01710_;
	assign _05187_ = _05186_ | ~_01713_;
	assign _05188_ = _05187_ | ~_01682_;
	assign _05189_ = _05188_ | _01680_;
	assign _05190_ = _05189_ & ~_01677_;
	assign _05191_ = _03030_ & ~_05190_;
	assign _05192_ = _01862_ & ~_01879_;
	assign _05193_ = _05192_ | _01882_;
	assign _05194_ = ~(_05193_ | _01884_);
	assign _05195_ = ~(_05194_ | _01886_);
	assign _05197_ = _05195_ | _01889_;
	assign _05198_ = _05197_ | ~_01891_;
	assign _05199_ = _05198_ | ~_01860_;
	assign _05200_ = _05199_ | _01858_;
	assign _05201_ = _05200_ & ~_01856_;
	assign _05202_ = _01719_ & ~_05201_;
	assign _05203_ = _05202_ | _05191_;
	assign _05204_ = ~_01919_;
	assign _05205_ = _05204_ & ~_01918_;
	assign _05206_ = _05205_ | _01922_;
	assign _05208_ = ~(_05206_ | _01924_);
	assign _05209_ = ~(_05208_ | _01926_);
	assign _05210_ = _05209_ | _01928_;
	assign _05211_ = _05210_ | ~_01931_;
	assign _05212_ = _05211_ | ~_01903_;
	assign _05213_ = ~(_05212_ | _01901_);
	assign _05214_ = ~(_05213_ | _01900_);
	assign _05215_ = _01898_ & ~_05214_;
	assign _05216_ = ~_01955_;
	assign _05217_ = _05216_ & ~_01953_;
	assign _05218_ = _05217_ | _01957_;
	assign _05219_ = ~(_05218_ | _01959_);
	assign _05220_ = ~(_05219_ | _01961_);
	assign _05221_ = _05220_ | _01963_;
	assign _05222_ = _05221_ | ~_01966_;
	assign _05223_ = _05222_ | ~_01942_;
	assign _05224_ = ~(_05223_ | _01940_);
	assign _05225_ = ~(_05224_ | _01939_);
	assign _05226_ = _01938_ & ~_05225_;
	assign _05227_ = _05226_ | _05215_;
	assign _05228_ = _05227_ | _05203_;
	assign _05229_ = ~(_03838_ | _03837_);
	assign _05230_ = _05229_ | _03841_;
	assign _05231_ = ~(_05230_ | _03844_);
	assign _05232_ = ~(_05231_ | _03846_);
	assign _05233_ = _05232_ | _03848_;
	assign _05234_ = _05233_ | ~_03851_;
	assign _05235_ = _05234_ | ~_03819_;
	assign _05236_ = ~(_05235_ | _03816_);
	assign _05237_ = ~(_05236_ | _03814_);
	assign _05239_ = _01975_ & ~_05237_;
	assign _05240_ = ~(_04018_ | _04017_);
	assign _05241_ = _05240_ | _04021_;
	assign _05242_ = ~(_05241_ | _04023_);
	assign _05243_ = ~(_05242_ | _04025_);
	assign _05244_ = _05243_ | _04028_;
	assign _05245_ = _05244_ | ~_04031_;
	assign _05246_ = _05245_ | ~_04000_;
	assign _05247_ = ~(_05246_ | _03997_);
	assign _05248_ = ~(_05247_ | _03995_);
	assign _05251_ = _03858_ & ~_05248_;
	assign _05252_ = _05251_ | _05239_;
	assign _05253_ = _04197_ & ~_04214_;
	assign _05254_ = _05253_ | _04217_;
	assign _05255_ = ~(_05254_ | _04219_);
	assign _05256_ = ~(_05255_ | _04221_);
	assign _05257_ = _05256_ | _04223_;
	assign _05258_ = _05257_ | ~_04225_;
	assign _05259_ = _05258_ | _04194_;
	assign _05260_ = ~(_05259_ | _04192_);
	assign _05262_ = _04725_ & ~_05260_;
	assign _05263_ = _04038_ & ~_05262_;
	assign _05264_ = _04375_ & ~_04391_;
	assign _05265_ = _05264_ | _04394_;
	assign _05266_ = ~(_05265_ | _04396_);
	assign _05267_ = ~(_05266_ | _04398_);
	assign _05268_ = _05267_ | _04400_;
	assign _05269_ = _05268_ | ~_04402_;
	assign _05270_ = _05269_ | _04371_;
	assign _05271_ = ~(_05270_ | _04369_);
	assign _05273_ = _04744_ & ~_05271_;
	assign _05274_ = _04232_ & ~_05273_;
	assign _05275_ = _05274_ | _05263_;
	assign _05276_ = _05275_ | _05252_;
	assign _05277_ = _05276_ | _05228_;
	assign _05278_ = _05277_ | _05180_;
	assign _05279_ = ~_04451_;
	assign _05280_ = _05279_ & ~_04450_;
	assign _05281_ = _05280_ | _04454_;
	assign _05282_ = ~(_05281_ | _04456_);
	assign _05284_ = ~(_05282_ | _04458_);
	assign _05285_ = _05284_ | _04461_;
	assign _05286_ = _05285_ | ~_04465_;
	assign _05287_ = _05286_ | _04467_;
	assign _05288_ = ~(_05287_ | _04469_);
	assign _05289_ = _05288_ | _04472_;
	assign io_out[3] = (_04428_ ? _05278_ : _05289_);
	assign _05290_ = _06185_ | _06175_;
	assign _05291_ = _05290_ | _06207_;
	assign _05292_ = ~(_05291_ | _06101_);
	assign _05294_ = _06022_ & ~_05292_;
	assign _05295_ = _05089_ & ~_05294_;
	assign _05296_ = ~(_05295_ | _06281_);
	assign _05297_ = _04475_ & ~_05296_;
	assign _05298_ = _05297_ | _06324_;
	assign _05299_ = _05298_ | _06346_;
	assign _05300_ = _05299_ | _06368_;
	assign _05301_ = _05300_ | _05581_;
	assign _05302_ = _05301_ | _05360_;
	assign _05303_ = _05302_ | _05141_;
	assign _05305_ = _04811_ & ~_05303_;
	assign _05306_ = _00219_ | _00208_;
	assign _05307_ = ~(_05306_ | _00252_);
	assign _05308_ = _05307_ & ~_00120_;
	assign _05309_ = _00109_ & ~_05308_;
	assign _05310_ = _05309_ | _00296_;
	assign _05311_ = _05310_ & ~_00329_;
	assign _05312_ = _04493_ & ~_05311_;
	assign _05313_ = _05312_ | _00372_;
	assign _05314_ = _05313_ | _00394_;
	assign _05316_ = _05314_ | _00415_;
	assign _05317_ = _05316_ | _00065_;
	assign _05318_ = _05317_ | _00043_;
	assign _05319_ = _05318_ | _00021_;
	assign _05320_ = _06455_ & ~_05319_;
	assign _05321_ = _00734_ | _00723_;
	assign _05322_ = ~(_05321_ | _00767_);
	assign _05323_ = _05322_ & ~_00635_;
	assign _05324_ = _00624_ & ~_05323_;
	assign _05325_ = _05324_ | _00811_;
	assign _05327_ = _05325_ & ~_00844_;
	assign _05328_ = _04510_ & ~_05327_;
	assign _05329_ = _05328_ | _00888_;
	assign _05330_ = _05329_ | _00910_;
	assign _05331_ = _05330_ | _00932_;
	assign _05332_ = _05331_ | _00580_;
	assign _05333_ = _05332_ | _00558_;
	assign _05334_ = _05333_ | _00536_;
	assign _05335_ = _00503_ & ~_05334_;
	assign _05336_ = _05335_ | _05320_;
	assign _05338_ = _05336_ | _05305_;
	assign _05339_ = _01273_ | _01262_;
	assign _05340_ = _05339_ | _01295_;
	assign _05341_ = ~(_05340_ | _01185_);
	assign _05342_ = _01174_ & ~_05341_;
	assign _05343_ = _05127_ & ~_05342_;
	assign _05344_ = ~(_05343_ | _01372_);
	assign _05345_ = _04530_ & ~_05344_;
	assign _05346_ = _05345_ | _01416_;
	assign _05347_ = _05346_ | _01438_;
	assign _05349_ = _05347_ | _01460_;
	assign _05350_ = _05349_ | _01130_;
	assign _05351_ = _05350_ | _01108_;
	assign _05352_ = _05351_ | _01086_;
	assign _05353_ = _01053_ & ~_05352_;
	assign _05354_ = _01756_ | _01745_;
	assign _05355_ = _05354_ | _01778_;
	assign _05356_ = ~(_05355_ | _01668_);
	assign _05357_ = _01657_ & ~_05356_;
	assign _05358_ = _05139_ & ~_05357_;
	assign _05361_ = ~(_05358_ | _01855_);
	assign _05362_ = _04548_ & ~_05361_;
	assign _05363_ = _05362_ | _01899_;
	assign _05364_ = _05363_ | _01921_;
	assign _05365_ = _05364_ | _01943_;
	assign _05366_ = _05365_ | _01614_;
	assign _05367_ = _05366_ | _01592_;
	assign _05368_ = _05367_ | _01570_;
	assign _05369_ = _01537_ & ~_05368_;
	assign _05370_ = _05369_ | _05353_;
	assign _05372_ = _02238_ | _02227_;
	assign _05373_ = _05372_ | _02260_;
	assign _05374_ = ~(_05373_ | _02152_);
	assign _05375_ = _02141_ & ~_05374_;
	assign _05376_ = _05154_ & ~_05375_;
	assign _05377_ = ~(_05376_ | _02337_);
	assign _05378_ = _04570_ & ~_05377_;
	assign _05379_ = _05378_ | _02381_;
	assign _05380_ = _05379_ | _02403_;
	assign _05381_ = _05380_ | _02425_;
	assign _05383_ = _05381_ | _02099_;
	assign _05384_ = _05383_ | _02079_;
	assign _05385_ = _05384_ | _02059_;
	assign _05386_ = _02028_ & ~_05385_;
	assign _05387_ = _02722_ | _02711_;
	assign _05388_ = _05387_ | _02744_;
	assign _05389_ = ~(_05388_ | _02634_);
	assign _05390_ = _02623_ & ~_05389_;
	assign _05391_ = _05166_ & ~_05390_;
	assign _05392_ = ~(_05391_ | _02821_);
	assign _05394_ = _04586_ & ~_05392_;
	assign _05395_ = _05394_ | _02865_;
	assign _05396_ = _05395_ | _02887_;
	assign _05397_ = _05396_ | _02909_;
	assign _05398_ = _05397_ | _02579_;
	assign _05399_ = _05398_ | _02557_;
	assign _05400_ = _05399_ | _02535_;
	assign _05401_ = _02502_ & ~_05400_;
	assign _05402_ = _05401_ | _05386_;
	assign _05403_ = _05402_ | _05370_;
	assign _05405_ = _05403_ | _05338_;
	assign _05406_ = _01694_ | _01693_;
	assign _05407_ = _05406_ | _01696_;
	assign _05408_ = ~(_05407_ | _01685_);
	assign _05409_ = _01699_ & ~_05408_;
	assign _05410_ = _01684_ & ~_05409_;
	assign _05411_ = ~(_05410_ | _01704_);
	assign _05412_ = ~(_05411_ | _01706_);
	assign _05413_ = _05412_ | _01708_;
	assign _05414_ = _05413_ | _01710_;
	assign _05416_ = _05414_ | ~_01713_;
	assign _05417_ = _05416_ | ~_01682_;
	assign _05418_ = _05417_ | _01680_;
	assign _05419_ = _05418_ | _01677_;
	assign _05420_ = _03030_ & ~_05419_;
	assign _05421_ = _01872_ | _01871_;
	assign _05422_ = _05421_ | _01874_;
	assign _05423_ = ~(_05422_ | _01863_);
	assign _05424_ = _01878_ & ~_05423_;
	assign _05425_ = _01862_ & ~_05424_;
	assign _05427_ = ~(_05425_ | _01882_);
	assign _05428_ = ~(_05427_ | _01884_);
	assign _05429_ = _05428_ | _01886_;
	assign _05430_ = _05429_ | _01889_;
	assign _05431_ = _05430_ | ~_01891_;
	assign _05432_ = _05431_ | ~_01860_;
	assign _05433_ = _05432_ | _01858_;
	assign _05434_ = _05433_ | _01856_;
	assign _05435_ = _01719_ & ~_05434_;
	assign _05436_ = _05435_ | _05420_;
	assign _05438_ = _01913_ | _01912_;
	assign _05439_ = _05438_ | _01915_;
	assign _05440_ = ~(_05439_ | _01905_);
	assign _05441_ = _01904_ & ~_05440_;
	assign _05442_ = _05204_ & ~_05441_;
	assign _05443_ = ~(_05442_ | _01922_);
	assign _05444_ = ~(_05443_ | _01924_);
	assign _05445_ = _05444_ | _01926_;
	assign _05446_ = _05445_ | _01928_;
	assign _05447_ = _05446_ | _01930_;
	assign _05449_ = _05447_ | _01902_;
	assign _05450_ = _05449_ | _01901_;
	assign _05451_ = _05450_ | _01900_;
	assign _05452_ = _01898_ & ~_05451_;
	assign _05453_ = _01374_ | ~_01340_;
	assign _05454_ = _05453_ | _01950_;
	assign _05455_ = ~(_05454_ | _01946_);
	assign _05456_ = _01945_ & ~_05455_;
	assign _05457_ = ~(_05456_ | _01955_);
	assign _05458_ = ~(_05457_ | _01957_);
	assign _05460_ = ~(_05458_ | _01959_);
	assign _05461_ = _05460_ | _01961_;
	assign _05462_ = _05461_ | _01963_;
	assign _05463_ = _05462_ | ~_01966_;
	assign _05464_ = _05463_ | ~_01942_;
	assign _05465_ = _05464_ | _01940_;
	assign _05466_ = _05465_ | _01939_;
	assign _05467_ = _01938_ & ~_05466_;
	assign _05468_ = _05467_ | _05452_;
	assign _05469_ = _05468_ | _05436_;
	assign _05472_ = _03831_ | _03830_;
	assign _05473_ = _05472_ | _03834_;
	assign _05474_ = ~(_05473_ | _03823_);
	assign _05475_ = _03822_ & ~_05474_;
	assign _05476_ = ~(_05475_ | _03838_);
	assign _05477_ = ~(_05476_ | _03841_);
	assign _05478_ = ~(_05477_ | _03844_);
	assign _05479_ = _05478_ | _03846_;
	assign _05480_ = _05479_ | _03848_;
	assign _05481_ = _05480_ | _03850_;
	assign _05483_ = _05481_ | _03818_;
	assign _05484_ = _05483_ | _03816_;
	assign _05485_ = _05484_ | _03814_;
	assign _05486_ = _01975_ & ~_05485_;
	assign _05487_ = _04011_ | _04010_;
	assign _05488_ = _05487_ | _04013_;
	assign _05489_ = ~(_05488_ | _04003_);
	assign _05490_ = _04002_ & ~_05489_;
	assign _05491_ = ~(_05490_ | _04018_);
	assign _05492_ = ~(_05491_ | _04021_);
	assign _05494_ = ~(_05492_ | _04023_);
	assign _05495_ = _05494_ | _04025_;
	assign _05496_ = _05495_ | _04028_;
	assign _05497_ = _05496_ | _04030_;
	assign _05498_ = _05497_ | _03999_;
	assign _05499_ = _05498_ | _03997_;
	assign _05500_ = _05499_ | _03995_;
	assign _05501_ = _03858_ & ~_05500_;
	assign _05502_ = _05501_ | _05486_;
	assign _05503_ = _04207_ | _04206_;
	assign _05505_ = _05503_ | _04210_;
	assign _05506_ = ~(_05505_ | _04199_);
	assign _05507_ = _04213_ & ~_05506_;
	assign _05508_ = _04197_ & ~_05507_;
	assign _05509_ = ~(_05508_ | _04217_);
	assign _05510_ = ~(_05509_ | _04219_);
	assign _05511_ = _05510_ | _04221_;
	assign _05512_ = _05511_ | _04223_;
	assign _05513_ = _05512_ | ~_04225_;
	assign _05514_ = _05513_ | ~_04195_;
	assign _05516_ = _05514_ | _04192_;
	assign _05517_ = _05516_ | _04190_;
	assign _05518_ = _04038_ & ~_05517_;
	assign _05519_ = _04385_ | _04383_;
	assign _05520_ = _05519_ | _04387_;
	assign _05521_ = ~(_05520_ | _04376_);
	assign _05522_ = _04390_ & ~_05521_;
	assign _05523_ = _04375_ & ~_05522_;
	assign _05524_ = ~(_05523_ | _04394_);
	assign _05525_ = ~(_05524_ | _04396_);
	assign _05527_ = _05525_ | _04398_;
	assign _05528_ = _05527_ | _04400_;
	assign _05529_ = _05528_ | ~_04402_;
	assign _05530_ = _05529_ | ~_04372_;
	assign _05531_ = _05530_ | _04369_;
	assign _05532_ = _05531_ | _04367_;
	assign _05533_ = _04232_ & ~_05532_;
	assign _05534_ = _05533_ | _05518_;
	assign _05535_ = _05534_ | _05502_;
	assign _05536_ = _05535_ | _05469_;
	assign _05538_ = _05536_ | _05405_;
	assign _05539_ = ~_04472_;
	assign _05540_ = _04444_ | _04442_;
	assign _05541_ = ~(_05540_ | _04446_);
	assign _05542_ = _05541_ & ~_04434_;
	assign _05543_ = _04432_ & ~_05542_;
	assign _05544_ = _05279_ & ~_05543_;
	assign _05545_ = ~(_05544_ | _04454_);
	assign _05546_ = _04770_ & ~_05545_;
	assign _05547_ = _05546_ | _04458_;
	assign _05549_ = _05547_ | _04461_;
	assign _05550_ = _05549_ | _04464_;
	assign _05551_ = _05550_ | _04467_;
	assign _05552_ = _05551_ | _04469_;
	assign _05553_ = _05539_ & ~_05552_;
	assign io_out[4] = (_04428_ ? _05538_ : _05553_);
	assign _05554_ = _06164_ | _06153_;
	assign _05555_ = ~(_05554_ | _06185_);
	assign _05556_ = _05555_ | _06207_;
	assign _05557_ = _05556_ | _06101_;
	assign _05559_ = _06022_ & ~_05557_;
	assign _05560_ = _05089_ & ~_05559_;
	assign _05561_ = _05560_ | _06281_;
	assign _05562_ = _05561_ | _06302_;
	assign _05563_ = _05562_ | _06324_;
	assign _05564_ = _05563_ | _06346_;
	assign _05565_ = _06379_ & ~_05564_;
	assign _05566_ = _05691_ & ~_05565_;
	assign _05567_ = _05566_ | _05360_;
	assign _05568_ = _05567_ | _05141_;
	assign _05570_ = _04811_ & ~_05568_;
	assign _05571_ = ~(_00197_ & _00175_);
	assign _05572_ = _00230_ & ~_05571_;
	assign _05573_ = _05572_ | _00252_;
	assign _05574_ = _05573_ | _00120_;
	assign _05575_ = _00109_ & ~_05574_;
	assign _05576_ = _05101_ & ~_05575_;
	assign _05577_ = _05576_ | _00329_;
	assign _05578_ = _05577_ | _00350_;
	assign _05579_ = _05578_ | _00372_;
	assign _05582_ = _05579_ | _00394_;
	assign _05583_ = _00426_ & ~_05582_;
	assign _05584_ = _00076_ & ~_05583_;
	assign _05585_ = _05584_ | _00043_;
	assign _05586_ = _05585_ | _00021_;
	assign _05587_ = _06455_ & ~_05586_;
	assign _05588_ = ~(_00712_ & _00690_);
	assign _05589_ = _00745_ & ~_05588_;
	assign _05590_ = _05589_ | _00767_;
	assign _05591_ = _05590_ | _00635_;
	assign _05593_ = _00624_ & ~_05591_;
	assign _05594_ = _05113_ & ~_05593_;
	assign _05595_ = _05594_ | _00844_;
	assign _05596_ = _05595_ | _00866_;
	assign _05597_ = _05596_ | _00888_;
	assign _05598_ = _05597_ | _00910_;
	assign _05599_ = _00943_ & ~_05598_;
	assign _05600_ = _00591_ & ~_05599_;
	assign _05601_ = _05600_ | _00558_;
	assign _05602_ = _05601_ | _00536_;
	assign _05603_ = _00503_ & ~_05602_;
	assign _05604_ = _05603_ | _05587_;
	assign _05605_ = _05604_ | _05570_;
	assign _05606_ = _01251_ | _01240_;
	assign _05607_ = ~(_05606_ | _01273_);
	assign _05608_ = _05607_ | _01295_;
	assign _05609_ = _05608_ | _01185_;
	assign _05610_ = _01174_ & ~_05609_;
	assign _05611_ = _05127_ & ~_05610_;
	assign _05612_ = _05611_ | _01372_;
	assign _05614_ = _05612_ | _01394_;
	assign _05615_ = _05614_ | _01416_;
	assign _05616_ = _05615_ | _01438_;
	assign _05617_ = _01471_ & ~_05616_;
	assign _05618_ = _01141_ & ~_05617_;
	assign _05619_ = _05618_ | _01108_;
	assign _05620_ = _05619_ | _01086_;
	assign _05621_ = _01053_ & ~_05620_;
	assign _05622_ = _01734_ | _01723_;
	assign _05623_ = ~(_05622_ | _01756_);
	assign _05625_ = _05623_ | _01778_;
	assign _05626_ = _05625_ | _01668_;
	assign _05627_ = _01657_ & ~_05626_;
	assign _05628_ = ~(_05627_ | _01822_);
	assign _05629_ = _05628_ | _01855_;
	assign _05630_ = _05629_ | _01877_;
	assign _05631_ = _05630_ | _01899_;
	assign _05632_ = _05631_ | _01921_;
	assign _05633_ = _01954_ & ~_05632_;
	assign _05634_ = _01625_ & ~_05633_;
	assign _05636_ = _05634_ | _01592_;
	assign _05637_ = _05636_ | _01570_;
	assign _05638_ = _01537_ & ~_05637_;
	assign _05639_ = _05638_ | _05621_;
	assign _05640_ = _02216_ | _02205_;
	assign _05641_ = ~(_05640_ | _02238_);
	assign _05642_ = _05641_ | _02260_;
	assign _05643_ = _05642_ | _02152_;
	assign _05644_ = _02141_ & ~_05643_;
	assign _05645_ = _05154_ & ~_05644_;
	assign _05647_ = _05645_ | _02337_;
	assign _05648_ = _05647_ | _02359_;
	assign _05649_ = _05648_ | _02381_;
	assign _05650_ = _05649_ | _02403_;
	assign _05651_ = _02436_ & ~_05650_;
	assign _05652_ = _02110_ & ~_05651_;
	assign _05653_ = _05652_ | _02079_;
	assign _05654_ = _05653_ | _02059_;
	assign _05655_ = _02028_ & ~_05654_;
	assign _05656_ = _02700_ | _02689_;
	assign _05658_ = ~(_05656_ | _02722_);
	assign _05659_ = _05658_ | _02744_;
	assign _05660_ = _05659_ | _02634_;
	assign _05661_ = _02623_ & ~_05660_;
	assign _05662_ = ~(_05661_ | _02788_);
	assign _05663_ = _05662_ | _02821_;
	assign _05664_ = _05663_ | _02843_;
	assign _05665_ = _05664_ | _02865_;
	assign _05666_ = _05665_ | _02887_;
	assign _05667_ = _02920_ & ~_05666_;
	assign _05669_ = _02590_ & ~_05667_;
	assign _05670_ = _05669_ | _02557_;
	assign _05671_ = _05670_ | _02535_;
	assign _05672_ = _02502_ & ~_05671_;
	assign _05673_ = _05672_ | _05655_;
	assign _05674_ = _05673_ | _05639_;
	assign _05675_ = _05674_ | _05605_;
	assign _05676_ = _01692_ | _01691_;
	assign _05677_ = ~(_05676_ | _01694_);
	assign _05678_ = _05677_ | _01696_;
	assign _05680_ = _05678_ | _01685_;
	assign _05681_ = _01699_ & ~_05680_;
	assign _05682_ = _01684_ & ~_05681_;
	assign _05683_ = _05682_ | _01704_;
	assign _05684_ = _05683_ | _01706_;
	assign _05685_ = _05684_ | _01708_;
	assign _05686_ = _05685_ | _01710_;
	assign _05687_ = _01713_ & ~_05686_;
	assign _05688_ = _01682_ & ~_05687_;
	assign _05689_ = _05688_ | _01680_;
	assign _05692_ = _05689_ | _01677_;
	assign _05693_ = _03030_ & ~_05692_;
	assign _05694_ = _01870_ | _01869_;
	assign _05695_ = ~(_05694_ | _01872_);
	assign _05696_ = _05695_ | _01874_;
	assign _05697_ = _05696_ | _01863_;
	assign _05698_ = _01878_ & ~_05697_;
	assign _05699_ = _01862_ & ~_05698_;
	assign _05700_ = _05699_ | _01882_;
	assign _05701_ = _05700_ | _01884_;
	assign _05703_ = _05701_ | _01886_;
	assign _05704_ = _05703_ | _01889_;
	assign _05705_ = _01891_ & ~_05704_;
	assign _05706_ = _01860_ & ~_05705_;
	assign _05707_ = _05706_ | _01858_;
	assign _05708_ = _05707_ | _01856_;
	assign _05709_ = _01719_ & ~_05708_;
	assign _05710_ = _05709_ | _05693_;
	assign _05711_ = _01911_ | _01909_;
	assign _05712_ = ~(_05711_ | _01913_);
	assign _05714_ = _05712_ | _01915_;
	assign _05715_ = _05714_ | _01905_;
	assign _05716_ = _01904_ & ~_05715_;
	assign _05717_ = ~(_05716_ | _01919_);
	assign _05718_ = _05717_ | _01922_;
	assign _05719_ = _05718_ | _01924_;
	assign _05720_ = _05719_ | _01926_;
	assign _05721_ = _05720_ | _01928_;
	assign _05722_ = _01931_ & ~_05721_;
	assign _05723_ = _01903_ & ~_05722_;
	assign _05725_ = _05723_ | _01901_;
	assign _05726_ = _05725_ | _01900_;
	assign _05727_ = _01898_ & ~_05726_;
	assign _05728_ = _04981_ & ~_04980_;
	assign _05729_ = _05728_ & ~_04979_;
	assign _05730_ = _05729_ & ~_01948_;
	assign _05731_ = _05730_ | _01950_;
	assign _05732_ = _05731_ | _01946_;
	assign _05733_ = _01945_ & ~_05732_;
	assign _05734_ = _05216_ & ~_05733_;
	assign _05736_ = _05734_ | _01957_;
	assign _05737_ = _05736_ | _01959_;
	assign _05738_ = _05737_ | _01961_;
	assign _05739_ = _05738_ | _01963_;
	assign _05740_ = _01966_ & ~_05739_;
	assign _05741_ = _01942_ & ~_05740_;
	assign _05742_ = _05741_ | _01940_;
	assign _05743_ = _05742_ | _01939_;
	assign _05744_ = _01938_ & ~_05743_;
	assign _05745_ = _05744_ | _05727_;
	assign _05747_ = _05745_ | _05710_;
	assign _05748_ = _03829_ | _03828_;
	assign _05749_ = ~(_05748_ | _03831_);
	assign _05750_ = _05749_ | _03834_;
	assign _05751_ = _05750_ | _03823_;
	assign _05752_ = _03822_ & ~_05751_;
	assign _05753_ = ~(_05752_ | _03838_);
	assign _05754_ = _05753_ | _03841_;
	assign _05755_ = _05754_ | _03844_;
	assign _05756_ = _05755_ | _03846_;
	assign _05758_ = _05756_ | _03848_;
	assign _05759_ = _03851_ & ~_05758_;
	assign _05760_ = _03819_ & ~_05759_;
	assign _05761_ = _05760_ | _03816_;
	assign _05762_ = _05761_ | _03814_;
	assign _05763_ = _01975_ & ~_05762_;
	assign _05764_ = _04009_ | _04008_;
	assign _05765_ = ~(_05764_ | _04011_);
	assign _05766_ = _05765_ | _04013_;
	assign _05767_ = _05766_ | _04003_;
	assign _05769_ = _04002_ & ~_05767_;
	assign _05770_ = ~(_05769_ | _04018_);
	assign _05771_ = _05770_ | _04021_;
	assign _05772_ = _05771_ | _04023_;
	assign _05773_ = _05772_ | _04025_;
	assign _05774_ = _05773_ | _04028_;
	assign _05775_ = _04031_ & ~_05774_;
	assign _05776_ = _04000_ & ~_05775_;
	assign _05777_ = _05776_ | _03997_;
	assign _05778_ = _05777_ | _03995_;
	assign _05780_ = _03858_ & ~_05778_;
	assign _05781_ = _05780_ | _05763_;
	assign _05782_ = _04205_ | _04204_;
	assign _05783_ = ~(_05782_ | _04207_);
	assign _05784_ = _05783_ | _04210_;
	assign _05785_ = _05784_ | _04199_;
	assign _05786_ = _04213_ & ~_05785_;
	assign _05787_ = _04197_ & ~_05786_;
	assign _05788_ = _05787_ | _04217_;
	assign _05789_ = _05788_ | _04219_;
	assign _05791_ = _05789_ | _04221_;
	assign _05792_ = _05791_ | _04223_;
	assign _05793_ = _04225_ & ~_05792_;
	assign _05794_ = _04195_ & ~_05793_;
	assign _05795_ = _05794_ | _04192_;
	assign _05796_ = _05795_ | _04190_;
	assign _05797_ = _04038_ & ~_05796_;
	assign _05798_ = _04382_ | _04381_;
	assign _05799_ = ~(_05798_ | _04385_);
	assign _05800_ = _05799_ | _04387_;
	assign _05803_ = _05800_ | _04376_;
	assign _05804_ = _04390_ & ~_05803_;
	assign _05805_ = _04375_ & ~_05804_;
	assign _05806_ = _05805_ | _04394_;
	assign _05807_ = _05806_ | _04396_;
	assign _05808_ = _05807_ | _04398_;
	assign _05809_ = _05808_ | _04400_;
	assign _05810_ = _04402_ & ~_05809_;
	assign _05811_ = _04372_ & ~_05810_;
	assign _05812_ = _05811_ | _04369_;
	assign _05814_ = _05812_ | _04367_;
	assign _05815_ = _04232_ & ~_05814_;
	assign _05816_ = _05815_ | _05797_;
	assign _05817_ = _05816_ | _05781_;
	assign _05818_ = _05817_ | _05747_;
	assign _05819_ = _05818_ | _05675_;
	assign _05820_ = _04441_ | _04440_;
	assign _05821_ = ~(_05820_ | _04444_);
	assign _05822_ = _05821_ | _04446_;
	assign _05823_ = _05822_ | _04434_;
	assign _05825_ = _04432_ & ~_05823_;
	assign _05826_ = _05279_ & ~_05825_;
	assign _05827_ = _05826_ | _04454_;
	assign _05828_ = _05827_ | _04456_;
	assign _05829_ = _05828_ | _04458_;
	assign _05830_ = _05829_ | _04461_;
	assign _05831_ = _04465_ & ~_05830_;
	assign _05832_ = _04769_ & ~_05831_;
	assign _05833_ = _05832_ | _04469_;
	assign _05834_ = _05539_ & ~_05833_;
	assign io_out[5] = (_04428_ ? _05819_ : _05834_);
	assign _05836_ = _06185_ | _06164_;
	assign _05837_ = _05836_ | _06207_;
	assign _05838_ = _05837_ | _06101_;
	assign _05839_ = _06022_ & ~_05838_;
	assign _05840_ = _05089_ & ~_05839_;
	assign _05841_ = _05840_ | _06281_;
	assign _05842_ = _05841_ | _06302_;
	assign _05843_ = _05842_ | _06324_;
	assign _05844_ = _04789_ & ~_05843_;
	assign _05846_ = _06379_ & ~_05844_;
	assign _05847_ = _05846_ | _05581_;
	assign _05848_ = _05847_ | _05360_;
	assign _05849_ = _05848_ | _05141_;
	assign _05850_ = _04811_ & ~_05849_;
	assign _05851_ = _00219_ | _00186_;
	assign _05852_ = _05851_ | _00252_;
	assign _05853_ = _05852_ | _00120_;
	assign _05854_ = _00109_ & ~_05853_;
	assign _05855_ = _05101_ & ~_05854_;
	assign _05857_ = _05855_ | _00329_;
	assign _05858_ = _05857_ | _00350_;
	assign _05859_ = _05858_ | _00372_;
	assign _05860_ = _04807_ & ~_05859_;
	assign _05861_ = _00426_ & ~_05860_;
	assign _05862_ = _05861_ | _00065_;
	assign _05863_ = _05862_ | _00043_;
	assign _05864_ = _05863_ | _00021_;
	assign _05865_ = _06455_ & ~_05864_;
	assign _05866_ = _00734_ | _00701_;
	assign _05868_ = _05866_ | _00767_;
	assign _05869_ = _05868_ | _00635_;
	assign _05870_ = _00624_ & ~_05869_;
	assign _05871_ = _05113_ & ~_05870_;
	assign _05872_ = _05871_ | _00844_;
	assign _05873_ = _05872_ | _00866_;
	assign _05874_ = _05873_ | _00888_;
	assign _05875_ = _04827_ & ~_05874_;
	assign _05876_ = _00943_ & ~_05875_;
	assign _05877_ = _05876_ | _00580_;
	assign _05879_ = _05877_ | _00558_;
	assign _05880_ = _05879_ | _00536_;
	assign _05881_ = _00503_ & ~_05880_;
	assign _05882_ = _05881_ | _05865_;
	assign _05883_ = _05882_ | _05850_;
	assign _05884_ = _01273_ | _01251_;
	assign _05885_ = _05884_ | _01295_;
	assign _05886_ = _05885_ | _01185_;
	assign _05887_ = _01174_ & ~_05886_;
	assign _05888_ = _05127_ & ~_05887_;
	assign _05890_ = _05888_ | _01372_;
	assign _05891_ = _05890_ | _01394_;
	assign _05892_ = _05891_ | _01416_;
	assign _05893_ = _04848_ & ~_05892_;
	assign _05894_ = _01471_ & ~_05893_;
	assign _05895_ = _05894_ | _01130_;
	assign _05896_ = _05895_ | _01108_;
	assign _05897_ = _05896_ | _01086_;
	assign _05898_ = _01053_ & ~_05897_;
	assign _05899_ = _01756_ | _01734_;
	assign _05901_ = _05899_ | _01778_;
	assign _05902_ = _05901_ | _01668_;
	assign _05903_ = _01657_ & ~_05902_;
	assign _05904_ = _05139_ & ~_05903_;
	assign _05905_ = _05904_ | _01855_;
	assign _05906_ = _05905_ | _01877_;
	assign _05907_ = _05906_ | _01899_;
	assign _05908_ = _04867_ & ~_05907_;
	assign _05909_ = _01954_ & ~_05908_;
	assign _05910_ = _05909_ | _01614_;
	assign _05913_ = _05910_ | _01592_;
	assign _05914_ = _05913_ | _01570_;
	assign _05915_ = _01537_ & ~_05914_;
	assign _05916_ = _05915_ | _05898_;
	assign _05917_ = _02238_ | _02216_;
	assign _05918_ = _05917_ | _02260_;
	assign _05919_ = _05918_ | _02152_;
	assign _05920_ = _02141_ & ~_05919_;
	assign _05921_ = _05154_ & ~_05920_;
	assign _05922_ = _05921_ | _02337_;
	assign _05924_ = _05922_ | _02359_;
	assign _05925_ = _05924_ | _02381_;
	assign _05926_ = _04885_ & ~_05925_;
	assign _05927_ = _02436_ & ~_05926_;
	assign _05928_ = _05927_ | _02099_;
	assign _05929_ = _05928_ | _02079_;
	assign _05930_ = _05929_ | _02059_;
	assign _05931_ = _02028_ & ~_05930_;
	assign _05932_ = _02722_ | _02700_;
	assign _05933_ = _05932_ | _02744_;
	assign _05935_ = _05933_ | _02634_;
	assign _05936_ = _02623_ & ~_05935_;
	assign _05937_ = _05166_ & ~_05936_;
	assign _05938_ = _05937_ | _02821_;
	assign _05939_ = _05938_ | _02843_;
	assign _05940_ = _05939_ | _02865_;
	assign _05941_ = _04904_ & ~_05940_;
	assign _05942_ = _02920_ & ~_05941_;
	assign _05943_ = _05942_ | _02579_;
	assign _05944_ = _05943_ | _02557_;
	assign _05946_ = _05944_ | _02535_;
	assign _05947_ = _02502_ & ~_05946_;
	assign _05948_ = _05947_ | _05931_;
	assign _05949_ = _05948_ | _05916_;
	assign _05950_ = _05949_ | _05883_;
	assign _05951_ = _01694_ | _01692_;
	assign _05952_ = _05951_ | _01696_;
	assign _05953_ = _05952_ | _01685_;
	assign _05954_ = _01699_ & ~_05953_;
	assign _05955_ = _01684_ & ~_05954_;
	assign _05957_ = _05955_ | _01704_;
	assign _05958_ = _05957_ | _01706_;
	assign _05959_ = _05958_ | _01708_;
	assign _05960_ = ~(_05959_ | _01710_);
	assign _05961_ = _01713_ & ~_05960_;
	assign _05962_ = _05961_ | ~_01682_;
	assign _05963_ = _05962_ | _01680_;
	assign _05964_ = _05963_ | _01677_;
	assign _05965_ = _03030_ & ~_05964_;
	assign _05966_ = _01872_ | _01870_;
	assign _05967_ = _05966_ | _01874_;
	assign _05968_ = _05967_ | _01863_;
	assign _05969_ = _01878_ & ~_05968_;
	assign _05970_ = _01862_ & ~_05969_;
	assign _05971_ = _05970_ | _01882_;
	assign _05972_ = _05971_ | _01884_;
	assign _05973_ = _05972_ | _01886_;
	assign _05974_ = ~(_05973_ | _01889_);
	assign _05975_ = _01891_ & ~_05974_;
	assign _05976_ = _05975_ | ~_01860_;
	assign _05978_ = _05976_ | _01858_;
	assign _05979_ = _05978_ | _01856_;
	assign _05980_ = _01719_ & ~_05979_;
	assign _05981_ = _05980_ | _05965_;
	assign _05982_ = _01913_ | _01911_;
	assign _05983_ = _05982_ | _01915_;
	assign _05984_ = _05983_ | _01905_;
	assign _05985_ = _01904_ & ~_05984_;
	assign _05986_ = _05204_ & ~_05985_;
	assign _05987_ = _05986_ | _01922_;
	assign _05989_ = _05987_ | _01924_;
	assign _05990_ = _05989_ | _01926_;
	assign _05991_ = _04960_ & ~_05990_;
	assign _05992_ = _01931_ & ~_05991_;
	assign _05993_ = _05992_ | _01902_;
	assign _05994_ = _05993_ | _01901_;
	assign _05995_ = _05994_ | _01900_;
	assign _05996_ = _01898_ & ~_05995_;
	assign _05997_ = _01948_ | _04979_;
	assign _05998_ = _05997_ | _01950_;
	assign _06000_ = _05998_ | _01946_;
	assign _06001_ = _01945_ & ~_06000_;
	assign _06002_ = _05216_ & ~_06001_;
	assign _06003_ = _06002_ | _01957_;
	assign _06004_ = _06003_ | _01959_;
	assign _06005_ = _06004_ | _01961_;
	assign _06006_ = _04978_ & ~_06005_;
	assign _06007_ = _01966_ & ~_06006_;
	assign _06008_ = _06007_ | _01941_;
	assign _06009_ = _06008_ | _01940_;
	assign _06011_ = _06009_ | _01939_;
	assign _06012_ = _01938_ & ~_06011_;
	assign _06013_ = _06012_ | _05996_;
	assign _06014_ = _06013_ | _05981_;
	assign _06015_ = _03831_ | _03829_;
	assign _06016_ = _06015_ | _03834_;
	assign _06017_ = _06016_ | _03823_;
	assign _06018_ = _03822_ & ~_06017_;
	assign _06019_ = ~(_06018_ | _03838_);
	assign _06020_ = _06019_ | _03841_;
	assign _06023_ = _06020_ | _03844_;
	assign _06024_ = _06023_ | _03846_;
	assign _06025_ = ~(_06024_ | _03848_);
	assign _06026_ = _03851_ & ~_06025_;
	assign _06027_ = _06026_ | _03818_;
	assign _06028_ = _06027_ | _03816_;
	assign _06029_ = _06028_ | _03814_;
	assign _06030_ = _01975_ & ~_06029_;
	assign _06031_ = _04011_ | _04009_;
	assign _06032_ = _06031_ | _04013_;
	assign _06033_ = _06032_ | _04003_;
	assign _06034_ = _04002_ & ~_06033_;
	assign _06035_ = ~(_06034_ | _04018_);
	assign _06036_ = _06035_ | _04021_;
	assign _06037_ = _06036_ | _04023_;
	assign _06038_ = _06037_ | _04025_;
	assign _06039_ = ~(_06038_ | _04028_);
	assign _06040_ = _04031_ & ~_06039_;
	assign _06041_ = _06040_ | _03999_;
	assign _06042_ = _06041_ | _03997_;
	assign _06043_ = _06042_ | _03995_;
	assign _06044_ = _03858_ & ~_06043_;
	assign _06045_ = _06044_ | _06030_;
	assign _06046_ = _04207_ | _04205_;
	assign _06047_ = _06046_ | _04210_;
	assign _06048_ = _06047_ | _04199_;
	assign _06049_ = _04213_ & ~_06048_;
	assign _06050_ = _04197_ & ~_06049_;
	assign _06051_ = _06050_ | _04217_;
	assign _06052_ = _06051_ | _04219_;
	assign _06053_ = _06052_ | _04221_;
	assign _06054_ = ~(_06053_ | _04223_);
	assign _06055_ = _04225_ & ~_06054_;
	assign _06056_ = _06055_ | ~_04195_;
	assign _06057_ = _06056_ | _04192_;
	assign _06058_ = _06057_ | _04190_;
	assign _06059_ = _04038_ & ~_06058_;
	assign _06060_ = _04385_ | _04382_;
	assign _06061_ = _06060_ | _04387_;
	assign _06062_ = _06061_ | _04376_;
	assign _06064_ = _04390_ & ~_06062_;
	assign _06065_ = _04375_ & ~_06064_;
	assign _06066_ = _06065_ | _04394_;
	assign _06067_ = _06066_ | _04396_;
	assign _06068_ = _06067_ | _04398_;
	assign _06069_ = ~(_06068_ | _04400_);
	assign _06070_ = _04402_ & ~_06069_;
	assign _06071_ = _06070_ | ~_04372_;
	assign _06072_ = _06071_ | _04369_;
	assign _06073_ = _06072_ | _04367_;
	assign _06075_ = _04232_ & ~_06073_;
	assign _06076_ = _06075_ | _06059_;
	assign _06077_ = _06076_ | _06045_;
	assign _06078_ = _06077_ | _06014_;
	assign _06079_ = _06078_ | _05950_;
	assign _06080_ = _04444_ | _04441_;
	assign _06081_ = _06080_ | _04446_;
	assign _06082_ = _06081_ | _04434_;
	assign _06083_ = _04432_ & ~_06082_;
	assign _06084_ = _05279_ & ~_06083_;
	assign _06086_ = _06084_ | _04454_;
	assign _06087_ = _06086_ | _04456_;
	assign _06088_ = _06087_ | _04458_;
	assign _06089_ = _05072_ & ~_06088_;
	assign _06090_ = _04465_ & ~_06089_;
	assign _06091_ = _06090_ | _04467_;
	assign _06092_ = _06091_ | _04469_;
	assign _06093_ = _05539_ & ~_06092_;
	assign io_out[6] = (_04428_ ? _06079_ : _06093_);
	assign \mchip.wrapper.nextState  = ~io_in[7];
	assign _06095_ = \mchip.wrapper.currState  & io_in[7];
	assign _06096_ = io_in[1] | ~io_in[0];
	assign \mchip.wrapper.keyReg.en  = _06095_ & ~_06096_;
	assign _06097_ = io_in[0] | ~io_in[1];
	assign \mchip.wrapper.intxtReg.en  = _06095_ & ~_06097_;
	always @(posedge io_in[12])
		if (\mchip.wrapper.intxtReg.en )
			\mchip.wrapper.intxtReg.Q [0] <= io_in[6];
	always @(posedge io_in[12])
		if (\mchip.wrapper.intxtReg.en )
			\mchip.wrapper.intxtReg.Q [1] <= \mchip.wrapper.intxtReg.Q [0];
	always @(posedge io_in[12])
		if (\mchip.wrapper.intxtReg.en )
			\mchip.wrapper.intxtReg.Q [2] <= \mchip.wrapper.intxtReg.Q [1];
	always @(posedge io_in[12])
		if (\mchip.wrapper.intxtReg.en )
			\mchip.wrapper.intxtReg.Q [3] <= \mchip.wrapper.intxtReg.Q [2];
	always @(posedge io_in[12])
		if (\mchip.wrapper.intxtReg.en )
			\mchip.wrapper.intxtReg.Q [4] <= \mchip.wrapper.intxtReg.Q [3];
	always @(posedge io_in[12])
		if (\mchip.wrapper.intxtReg.en )
			\mchip.wrapper.intxtReg.Q [5] <= \mchip.wrapper.intxtReg.Q [4];
	always @(posedge io_in[12])
		if (\mchip.wrapper.intxtReg.en )
			\mchip.wrapper.intxtReg.Q [6] <= \mchip.wrapper.intxtReg.Q [5];
	always @(posedge io_in[12])
		if (\mchip.wrapper.intxtReg.en )
			\mchip.wrapper.intxtReg.Q [7] <= \mchip.wrapper.intxtReg.Q [6];
	always @(posedge io_in[12])
		if (\mchip.wrapper.intxtReg.en )
			\mchip.wrapper.intxtReg.Q [8] <= \mchip.wrapper.intxtReg.Q [7];
	always @(posedge io_in[12])
		if (\mchip.wrapper.intxtReg.en )
			\mchip.wrapper.intxtReg.Q [9] <= \mchip.wrapper.intxtReg.Q [8];
	always @(posedge io_in[12])
		if (\mchip.wrapper.intxtReg.en )
			\mchip.wrapper.intxtReg.Q [10] <= \mchip.wrapper.intxtReg.Q [9];
	always @(posedge io_in[12])
		if (\mchip.wrapper.intxtReg.en )
			\mchip.wrapper.intxtReg.Q [11] <= \mchip.wrapper.intxtReg.Q [10];
	always @(posedge io_in[12])
		if (\mchip.wrapper.intxtReg.en )
			\mchip.wrapper.intxtReg.Q [12] <= \mchip.wrapper.intxtReg.Q [11];
	always @(posedge io_in[12])
		if (\mchip.wrapper.intxtReg.en )
			\mchip.wrapper.intxtReg.Q [13] <= \mchip.wrapper.intxtReg.Q [12];
	always @(posedge io_in[12])
		if (\mchip.wrapper.intxtReg.en )
			\mchip.wrapper.intxtReg.Q [14] <= \mchip.wrapper.intxtReg.Q [13];
	always @(posedge io_in[12])
		if (\mchip.wrapper.intxtReg.en )
			\mchip.wrapper.intxtReg.Q [15] <= \mchip.wrapper.intxtReg.Q [14];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.wrapper.currState  <= 1'h1;
		else
			\mchip.wrapper.currState  <= \mchip.wrapper.nextState ;
	always @(posedge io_in[12])
		if (\mchip.wrapper.keyReg.en )
			\mchip.wrapper.keyReg.Q [0] <= io_in[6];
	always @(posedge io_in[12])
		if (\mchip.wrapper.keyReg.en )
			\mchip.wrapper.keyReg.Q [1] <= \mchip.wrapper.keyReg.Q [0];
	always @(posedge io_in[12])
		if (\mchip.wrapper.keyReg.en )
			\mchip.wrapper.keyReg.Q [2] <= \mchip.wrapper.keyReg.Q [1];
	always @(posedge io_in[12])
		if (\mchip.wrapper.keyReg.en )
			\mchip.wrapper.keyReg.Q [3] <= \mchip.wrapper.keyReg.Q [2];
	always @(posedge io_in[12])
		if (\mchip.wrapper.keyReg.en )
			\mchip.wrapper.keyReg.Q [4] <= \mchip.wrapper.keyReg.Q [3];
	always @(posedge io_in[12])
		if (\mchip.wrapper.keyReg.en )
			\mchip.wrapper.keyReg.Q [5] <= \mchip.wrapper.keyReg.Q [4];
	always @(posedge io_in[12])
		if (\mchip.wrapper.keyReg.en )
			\mchip.wrapper.keyReg.Q [6] <= \mchip.wrapper.keyReg.Q [5];
	always @(posedge io_in[12])
		if (\mchip.wrapper.keyReg.en )
			\mchip.wrapper.keyReg.Q [7] <= \mchip.wrapper.keyReg.Q [6];
	always @(posedge io_in[12])
		if (\mchip.wrapper.keyReg.en )
			\mchip.wrapper.keyReg.Q [8] <= \mchip.wrapper.keyReg.Q [7];
	always @(posedge io_in[12])
		if (\mchip.wrapper.keyReg.en )
			\mchip.wrapper.keyReg.Q [9] <= \mchip.wrapper.keyReg.Q [8];
	always @(posedge io_in[12])
		if (\mchip.wrapper.keyReg.en )
			\mchip.wrapper.keyReg.Q [10] <= \mchip.wrapper.keyReg.Q [9];
	always @(posedge io_in[12])
		if (\mchip.wrapper.keyReg.en )
			\mchip.wrapper.keyReg.Q [11] <= \mchip.wrapper.keyReg.Q [10];
	always @(posedge io_in[12])
		if (\mchip.wrapper.keyReg.en )
			\mchip.wrapper.keyReg.Q [12] <= \mchip.wrapper.keyReg.Q [11];
	always @(posedge io_in[12])
		if (\mchip.wrapper.keyReg.en )
			\mchip.wrapper.keyReg.Q [13] <= \mchip.wrapper.keyReg.Q [12];
	always @(posedge io_in[12])
		if (\mchip.wrapper.keyReg.en )
			\mchip.wrapper.keyReg.Q [14] <= \mchip.wrapper.keyReg.Q [13];
	always @(posedge io_in[12])
		if (\mchip.wrapper.keyReg.en )
			\mchip.wrapper.keyReg.Q [15] <= \mchip.wrapper.keyReg.Q [14];
	assign io_out[13:7] = 7'h01;
	assign \mchip.clock  = io_in[12];
	assign \mchip.io_in  = io_in[11:0];
	assign \mchip.io_out  = {5'h01, io_out[6:0]};
	assign \mchip.reset  = io_in[13];
	assign \mchip.wrapper.clock  = io_in[12];
	assign \mchip.wrapper.de.KEY  = \mchip.wrapper.keyReg.Q ;
	assign \mchip.wrapper.de.P1  = {\mchip.wrapper.keyReg.Q [7:6], 1'h0, \mchip.wrapper.keyReg.Q [4:3], 1'h0, \mchip.wrapper.keyReg.Q [1:0]};
	assign \mchip.wrapper.de.intxt  = \mchip.wrapper.intxtReg.Q ;
	assign \mchip.wrapper.de.p1start  = 8'h24;
	assign \mchip.wrapper.de.p2start  = 8'h3f;
	assign \mchip.wrapper.de.p3start  = 8'h6a;
	assign \mchip.wrapper.de.p4start  = 8'h88;
	assign \mchip.wrapper.de.p5start  = 8'h85;
	assign \mchip.wrapper.de.p6start  = 8'ha3;
	assign \mchip.wrapper.de.p7start  = 8'h08;
	assign \mchip.wrapper.de.p8start  = 8'hd3;
	assign \mchip.wrapper.de.s11  = {\mchip.wrapper.keyReg.Q [7:5], 1'h0, \mchip.wrapper.keyReg.Q [3:2], 2'h0};
	assign \mchip.wrapper.de.sub1.s1  = {\mchip.wrapper.keyReg.Q [7:5], 1'h0, \mchip.wrapper.keyReg.Q [3:2], 2'h0};
	assign \mchip.wrapper.de.sub17.s1  = {\mchip.wrapper.keyReg.Q [7:5], 1'h0, \mchip.wrapper.keyReg.Q [3:2], 2'h0};
	assign \mchip.wrapper.de.sub25.s1  = {\mchip.wrapper.keyReg.Q [7:5], 1'h0, \mchip.wrapper.keyReg.Q [3:2], 2'h0};
	assign \mchip.wrapper.de.sub29.s1  = {\mchip.wrapper.keyReg.Q [7:5], 1'h0, \mchip.wrapper.keyReg.Q [3:2], 2'h0};
	assign \mchip.wrapper.de.sub37.s1  = {\mchip.wrapper.keyReg.Q [7:5], 1'h0, \mchip.wrapper.keyReg.Q [3:2], 2'h0};
	assign \mchip.wrapper.de.sub45.s1  = {\mchip.wrapper.keyReg.Q [7:5], 1'h0, \mchip.wrapper.keyReg.Q [3:2], 2'h0};
	assign \mchip.wrapper.de.sub5.s1  = {\mchip.wrapper.keyReg.Q [7:5], 1'h0, \mchip.wrapper.keyReg.Q [3:2], 2'h0};
	assign \mchip.wrapper.de.sub9.s1  = {\mchip.wrapper.keyReg.Q [7:5], 1'h0, \mchip.wrapper.keyReg.Q [3:2], 2'h0};
	assign \mchip.wrapper.de.temp8  = \mchip.wrapper.intxtReg.Q ;
	assign \mchip.wrapper.display_sel  = io_in[5:2];
	assign \mchip.wrapper.en.KEY  = \mchip.wrapper.keyReg.Q ;
	assign \mchip.wrapper.en.P1  = {\mchip.wrapper.keyReg.Q [7:6], 1'h0, \mchip.wrapper.keyReg.Q [4:3], 1'h0, \mchip.wrapper.keyReg.Q [1:0]};
	assign \mchip.wrapper.en.intxt  = \mchip.wrapper.intxtReg.Q ;
	assign \mchip.wrapper.en.p1start  = 8'h24;
	assign \mchip.wrapper.en.p2start  = 8'h3f;
	assign \mchip.wrapper.en.p3start  = 8'h6a;
	assign \mchip.wrapper.en.p4start  = 8'h88;
	assign \mchip.wrapper.en.p5start  = 8'h85;
	assign \mchip.wrapper.en.p6start  = 8'ha3;
	assign \mchip.wrapper.en.p7start  = 8'h08;
	assign \mchip.wrapper.en.p8start  = 8'hd3;
	assign \mchip.wrapper.en.s11  = {\mchip.wrapper.keyReg.Q [7:5], 1'h0, \mchip.wrapper.keyReg.Q [3:2], 2'h0};
	assign \mchip.wrapper.en.sub1.s1  = {\mchip.wrapper.keyReg.Q [7:5], 1'h0, \mchip.wrapper.keyReg.Q [3:2], 2'h0};
	assign \mchip.wrapper.en.sub1.sel  = \mchip.wrapper.intxtReg.Q [15:14];
	assign \mchip.wrapper.en.sub17.s1  = {\mchip.wrapper.keyReg.Q [7:5], 1'h0, \mchip.wrapper.keyReg.Q [3:2], 2'h0};
	assign \mchip.wrapper.en.sub2.sel  = \mchip.wrapper.intxtReg.Q [13:12];
	assign \mchip.wrapper.en.sub25.s1  = {\mchip.wrapper.keyReg.Q [7:5], 1'h0, \mchip.wrapper.keyReg.Q [3:2], 2'h0};
	assign \mchip.wrapper.en.sub29.s1  = {\mchip.wrapper.keyReg.Q [7:5], 1'h0, \mchip.wrapper.keyReg.Q [3:2], 2'h0};
	assign \mchip.wrapper.en.sub3.sel  = \mchip.wrapper.intxtReg.Q [11:10];
	assign \mchip.wrapper.en.sub37.s1  = {\mchip.wrapper.keyReg.Q [7:5], 1'h0, \mchip.wrapper.keyReg.Q [3:2], 2'h0};
	assign \mchip.wrapper.en.sub4.sel  = \mchip.wrapper.intxtReg.Q [9:8];
	assign \mchip.wrapper.en.sub45.s1  = {\mchip.wrapper.keyReg.Q [7:5], 1'h0, \mchip.wrapper.keyReg.Q [3:2], 2'h0};
	assign \mchip.wrapper.en.sub5.s1  = {\mchip.wrapper.keyReg.Q [7:5], 1'h0, \mchip.wrapper.keyReg.Q [3:2], 2'h0};
	assign \mchip.wrapper.en.sub9.s1  = {\mchip.wrapper.keyReg.Q [7:5], 1'h0, \mchip.wrapper.keyReg.Q [3:2], 2'h0};
	assign \mchip.wrapper.hex_out  = {1'h1, io_out[6:0]};
	assign \mchip.wrapper.i1.hexdigit  = \mchip.wrapper.intxtReg.Q [3:0];
	assign \mchip.wrapper.i1.seg  = 8'h80;
	assign \mchip.wrapper.i10.seg  = 8'h80;
	assign \mchip.wrapper.i11.seg  = 8'h80;
	assign \mchip.wrapper.i12.seg  = 8'h80;
	assign \mchip.wrapper.i13.seg  = 8'h80;
	assign \mchip.wrapper.i14.seg  = 8'h80;
	assign \mchip.wrapper.i15.seg  = 8'h80;
	assign \mchip.wrapper.i16.seg  = 8'h80;
	assign \mchip.wrapper.i2.hexdigit  = \mchip.wrapper.intxtReg.Q [7:4];
	assign \mchip.wrapper.i2.seg  = 8'h80;
	assign \mchip.wrapper.i3.hexdigit  = \mchip.wrapper.intxtReg.Q [11:8];
	assign \mchip.wrapper.i3.seg  = 8'h80;
	assign \mchip.wrapper.i4.hexdigit  = \mchip.wrapper.intxtReg.Q [15:12];
	assign \mchip.wrapper.i4.seg  = 8'h80;
	assign \mchip.wrapper.i5.hexdigit  = \mchip.wrapper.keyReg.Q [3:0];
	assign \mchip.wrapper.i5.seg  = 8'h80;
	assign \mchip.wrapper.i6.hexdigit  = \mchip.wrapper.keyReg.Q [7:4];
	assign \mchip.wrapper.i6.seg  = 8'h80;
	assign \mchip.wrapper.i7.hexdigit  = \mchip.wrapper.keyReg.Q [11:8];
	assign \mchip.wrapper.i7.seg  = 8'h80;
	assign \mchip.wrapper.i8.hexdigit  = \mchip.wrapper.keyReg.Q [15:12];
	assign \mchip.wrapper.i8.seg  = 8'h80;
	assign \mchip.wrapper.i9.seg  = 8'h80;
	assign \mchip.wrapper.in_bit  = io_in[6];
	assign \mchip.wrapper.intxt  = \mchip.wrapper.intxtReg.Q ;
	assign \mchip.wrapper.intxtReg.clock  = io_in[12];
	assign \mchip.wrapper.intxtReg.left  = 1'h1;
	assign \mchip.wrapper.intxtReg.serial  = io_in[6];
	assign \mchip.wrapper.intxt_hex1  = 8'h80;
	assign \mchip.wrapper.intxt_hex2  = 8'h80;
	assign \mchip.wrapper.intxt_hex3  = 8'h80;
	assign \mchip.wrapper.intxt_hex4  = 8'h80;
	assign \mchip.wrapper.key  = \mchip.wrapper.keyReg.Q ;
	assign \mchip.wrapper.keyReg.clock  = io_in[12];
	assign \mchip.wrapper.keyReg.left  = 1'h1;
	assign \mchip.wrapper.keyReg.serial  = io_in[6];
	assign \mchip.wrapper.key_hex1  = 8'h80;
	assign \mchip.wrapper.key_hex2  = 8'h80;
	assign \mchip.wrapper.key_hex3  = 8'h80;
	assign \mchip.wrapper.key_hex4  = 8'h80;
	assign \mchip.wrapper.mode_sel  = io_in[1:0];
	assign \mchip.wrapper.outtxt_de_hex1  = 8'h80;
	assign \mchip.wrapper.outtxt_de_hex2  = 8'h80;
	assign \mchip.wrapper.outtxt_de_hex3  = 8'h80;
	assign \mchip.wrapper.outtxt_de_hex4  = 8'h80;
	assign \mchip.wrapper.outtxt_hex1  = 8'h80;
	assign \mchip.wrapper.outtxt_hex2  = 8'h80;
	assign \mchip.wrapper.outtxt_hex3  = 8'h80;
	assign \mchip.wrapper.outtxt_hex4  = 8'h80;
	assign \mchip.wrapper.ready  = io_in[7];
	assign \mchip.wrapper.reset  = io_in[13];
endmodule
module d20_rashik_tetris (
	io_in,
	io_out
);
	wire _0000_;
	wire _0001_;
	wire _0002_;
	wire _0003_;
	wire _0004_;
	wire _0005_;
	wire _0006_;
	wire _0007_;
	wire _0008_;
	wire _0009_;
	wire _0010_;
	wire _0011_;
	wire _0012_;
	wire _0013_;
	wire _0014_;
	wire _0015_;
	wire _0016_;
	wire _0017_;
	wire _0018_;
	wire _0019_;
	wire _0020_;
	wire _0021_;
	wire _0022_;
	wire _0023_;
	wire _0024_;
	wire _0025_;
	wire _0026_;
	wire _0027_;
	wire _0028_;
	wire _0029_;
	wire _0030_;
	wire _0031_;
	wire _0032_;
	wire _0033_;
	wire _0034_;
	wire _0035_;
	wire _0036_;
	wire _0037_;
	wire _0038_;
	wire _0039_;
	wire _0040_;
	wire _0041_;
	wire _0042_;
	wire _0043_;
	wire _0044_;
	wire _0045_;
	wire _0046_;
	wire _0047_;
	wire _0048_;
	wire _0049_;
	wire _0050_;
	wire _0051_;
	wire _0052_;
	wire _0053_;
	wire _0054_;
	wire _0055_;
	wire _0056_;
	wire _0057_;
	wire _0058_;
	wire _0059_;
	wire _0060_;
	wire _0061_;
	wire _0062_;
	wire _0063_;
	wire _0064_;
	wire _0065_;
	wire _0066_;
	wire _0067_;
	wire _0068_;
	wire _0069_;
	wire _0070_;
	wire _0071_;
	wire _0072_;
	wire _0073_;
	wire _0074_;
	wire _0075_;
	wire _0076_;
	wire _0077_;
	wire _0078_;
	wire _0079_;
	wire _0080_;
	wire _0081_;
	wire _0082_;
	wire _0083_;
	wire _0084_;
	wire _0085_;
	wire _0086_;
	wire _0087_;
	wire _0088_;
	wire _0089_;
	wire _0090_;
	wire _0091_;
	wire _0092_;
	wire _0093_;
	wire _0094_;
	wire _0095_;
	wire _0096_;
	wire _0097_;
	wire _0098_;
	wire _0099_;
	wire _0100_;
	wire _0101_;
	wire _0102_;
	wire _0103_;
	wire _0104_;
	wire _0105_;
	wire _0106_;
	wire _0107_;
	wire _0108_;
	wire _0109_;
	wire _0110_;
	wire _0111_;
	wire _0112_;
	wire _0113_;
	wire _0114_;
	wire _0115_;
	wire _0116_;
	wire _0117_;
	wire _0118_;
	wire _0119_;
	wire _0120_;
	wire _0121_;
	wire _0122_;
	wire _0123_;
	wire _0124_;
	wire _0125_;
	wire _0126_;
	wire _0127_;
	wire _0128_;
	wire _0129_;
	wire _0130_;
	wire _0131_;
	wire _0132_;
	wire _0133_;
	wire _0134_;
	wire _0135_;
	wire _0136_;
	wire _0137_;
	wire _0138_;
	wire _0139_;
	wire _0140_;
	wire _0141_;
	wire _0142_;
	wire _0143_;
	wire _0144_;
	wire _0145_;
	wire _0146_;
	wire _0147_;
	wire _0148_;
	wire _0149_;
	wire _0150_;
	wire _0151_;
	wire _0152_;
	wire _0153_;
	wire _0154_;
	wire _0155_;
	wire _0156_;
	wire _0157_;
	wire _0158_;
	wire _0159_;
	wire _0160_;
	wire _0161_;
	wire _0162_;
	wire _0163_;
	wire _0164_;
	wire _0165_;
	wire _0166_;
	wire _0167_;
	wire _0168_;
	wire _0169_;
	wire _0170_;
	wire _0171_;
	wire _0172_;
	wire _0173_;
	wire _0174_;
	wire _0175_;
	wire _0176_;
	wire _0177_;
	wire _0178_;
	wire _0179_;
	wire _0180_;
	wire _0181_;
	wire _0182_;
	wire _0183_;
	wire _0184_;
	wire _0185_;
	wire _0186_;
	wire _0187_;
	wire _0188_;
	wire _0189_;
	wire _0190_;
	wire _0191_;
	wire _0192_;
	wire _0193_;
	wire _0194_;
	wire _0195_;
	wire _0196_;
	wire _0197_;
	wire _0198_;
	wire _0199_;
	wire _0200_;
	wire _0201_;
	wire _0202_;
	wire _0203_;
	wire _0204_;
	wire _0205_;
	wire _0206_;
	wire _0207_;
	wire _0208_;
	wire _0209_;
	wire _0210_;
	wire _0211_;
	wire _0212_;
	wire _0213_;
	wire _0214_;
	wire _0215_;
	wire _0216_;
	wire _0217_;
	wire _0218_;
	wire _0219_;
	wire _0220_;
	wire _0221_;
	wire _0222_;
	wire _0223_;
	wire _0224_;
	wire _0225_;
	wire _0226_;
	wire _0227_;
	wire _0228_;
	wire _0229_;
	wire _0230_;
	wire _0231_;
	wire _0232_;
	wire _0233_;
	wire _0234_;
	wire _0235_;
	wire _0236_;
	wire _0237_;
	wire _0238_;
	wire _0239_;
	wire _0240_;
	wire _0241_;
	wire _0242_;
	wire _0243_;
	wire _0244_;
	wire _0245_;
	wire _0246_;
	wire _0247_;
	wire _0248_;
	wire _0249_;
	wire _0250_;
	wire _0251_;
	wire _0252_;
	wire _0253_;
	wire _0254_;
	wire _0255_;
	wire _0256_;
	wire _0257_;
	wire _0258_;
	wire _0259_;
	wire _0260_;
	wire _0261_;
	wire _0262_;
	wire _0263_;
	wire _0264_;
	wire _0265_;
	wire _0266_;
	wire _0267_;
	wire _0268_;
	wire _0269_;
	wire _0270_;
	wire _0271_;
	wire _0272_;
	wire _0273_;
	wire _0274_;
	wire _0275_;
	wire _0276_;
	wire _0277_;
	wire _0278_;
	wire _0279_;
	wire _0280_;
	wire _0281_;
	wire _0282_;
	wire _0283_;
	wire _0284_;
	wire _0285_;
	wire _0286_;
	wire _0287_;
	wire _0288_;
	wire _0289_;
	wire _0290_;
	wire _0291_;
	wire _0292_;
	wire _0293_;
	wire _0294_;
	wire _0295_;
	wire _0296_;
	wire _0297_;
	wire _0298_;
	wire _0299_;
	wire _0300_;
	wire _0301_;
	wire _0302_;
	wire _0303_;
	wire _0304_;
	wire _0305_;
	wire _0306_;
	wire _0307_;
	wire _0308_;
	wire _0309_;
	wire _0310_;
	wire _0311_;
	wire _0312_;
	wire _0313_;
	wire _0314_;
	wire _0315_;
	wire _0316_;
	wire _0317_;
	wire _0318_;
	wire _0319_;
	wire _0320_;
	wire _0321_;
	wire _0322_;
	wire _0323_;
	wire _0324_;
	wire _0325_;
	wire _0326_;
	wire _0327_;
	wire _0328_;
	wire _0329_;
	wire _0330_;
	wire _0331_;
	wire _0332_;
	wire _0333_;
	wire _0334_;
	wire _0335_;
	wire _0336_;
	wire _0337_;
	wire _0338_;
	wire _0339_;
	wire _0340_;
	wire _0341_;
	wire _0342_;
	wire _0343_;
	wire _0344_;
	wire _0345_;
	wire _0346_;
	wire _0347_;
	wire _0348_;
	wire _0349_;
	wire _0350_;
	wire _0351_;
	wire _0352_;
	wire _0353_;
	wire _0354_;
	wire _0355_;
	wire _0356_;
	wire _0357_;
	wire _0358_;
	wire _0359_;
	wire _0360_;
	wire _0361_;
	wire _0362_;
	wire _0363_;
	wire _0364_;
	wire _0365_;
	wire _0366_;
	wire _0367_;
	wire _0368_;
	wire _0369_;
	wire _0370_;
	wire _0371_;
	wire _0372_;
	wire _0373_;
	wire _0374_;
	wire _0375_;
	wire _0376_;
	wire _0377_;
	wire _0378_;
	wire _0379_;
	wire _0380_;
	wire _0381_;
	wire _0382_;
	wire _0383_;
	wire _0384_;
	wire _0385_;
	wire _0386_;
	wire _0387_;
	wire _0388_;
	wire _0389_;
	wire _0390_;
	wire _0391_;
	wire _0392_;
	wire _0393_;
	wire _0394_;
	wire _0395_;
	wire _0396_;
	wire _0397_;
	wire _0398_;
	wire _0399_;
	wire _0400_;
	wire _0401_;
	wire _0402_;
	wire _0403_;
	wire _0404_;
	wire _0405_;
	wire _0406_;
	wire _0407_;
	wire _0408_;
	wire _0409_;
	wire _0410_;
	wire _0411_;
	wire _0412_;
	wire _0413_;
	wire _0414_;
	wire _0415_;
	wire _0416_;
	wire _0417_;
	wire _0418_;
	wire _0419_;
	wire _0420_;
	wire _0421_;
	wire _0422_;
	wire _0423_;
	wire _0424_;
	wire _0425_;
	wire _0426_;
	wire _0427_;
	wire _0428_;
	wire _0429_;
	wire _0430_;
	wire _0431_;
	wire _0432_;
	wire _0433_;
	wire _0434_;
	wire _0435_;
	wire _0436_;
	wire _0437_;
	wire _0438_;
	wire _0439_;
	wire _0440_;
	wire _0441_;
	wire _0442_;
	wire _0443_;
	wire _0444_;
	wire _0445_;
	wire _0446_;
	wire _0447_;
	wire _0448_;
	wire _0449_;
	wire _0450_;
	wire _0451_;
	wire _0452_;
	wire _0453_;
	wire _0454_;
	wire _0455_;
	wire _0456_;
	wire _0457_;
	wire _0458_;
	wire _0459_;
	wire _0460_;
	wire _0461_;
	wire _0462_;
	wire _0463_;
	wire _0464_;
	wire _0465_;
	wire _0466_;
	wire _0467_;
	wire _0468_;
	wire _0469_;
	wire _0470_;
	wire _0471_;
	wire _0472_;
	wire _0473_;
	wire _0474_;
	wire _0475_;
	wire _0476_;
	wire _0477_;
	wire _0478_;
	wire _0479_;
	wire _0480_;
	wire _0481_;
	wire _0482_;
	wire _0483_;
	wire _0484_;
	wire _0485_;
	wire _0486_;
	wire _0487_;
	wire _0488_;
	wire _0489_;
	wire _0490_;
	wire _0491_;
	wire _0492_;
	wire _0493_;
	wire _0494_;
	wire _0495_;
	wire _0496_;
	wire _0497_;
	wire _0498_;
	wire _0499_;
	wire _0500_;
	wire _0501_;
	wire _0502_;
	wire _0503_;
	wire _0504_;
	wire _0505_;
	wire _0506_;
	wire _0507_;
	wire _0508_;
	wire _0509_;
	wire _0510_;
	wire _0511_;
	wire _0512_;
	wire _0513_;
	wire _0514_;
	wire _0515_;
	wire _0516_;
	wire _0517_;
	wire _0518_;
	wire _0519_;
	wire _0520_;
	wire _0521_;
	wire _0522_;
	wire _0523_;
	wire _0524_;
	wire _0525_;
	wire _0526_;
	wire _0527_;
	wire _0528_;
	wire _0529_;
	wire _0530_;
	wire _0531_;
	wire _0532_;
	wire _0533_;
	wire _0534_;
	wire _0535_;
	wire _0536_;
	wire _0537_;
	wire _0538_;
	wire _0539_;
	wire _0540_;
	wire _0541_;
	wire _0542_;
	wire _0543_;
	wire _0544_;
	wire _0545_;
	wire _0546_;
	wire _0547_;
	wire _0548_;
	wire _0549_;
	wire _0550_;
	wire _0551_;
	wire _0552_;
	wire _0553_;
	wire _0554_;
	wire _0555_;
	wire _0556_;
	wire _0557_;
	wire _0558_;
	wire _0559_;
	wire _0560_;
	wire _0561_;
	wire _0562_;
	wire _0563_;
	wire _0564_;
	wire _0565_;
	wire _0566_;
	wire _0567_;
	wire _0568_;
	wire _0569_;
	wire _0570_;
	wire _0571_;
	wire _0572_;
	wire _0573_;
	wire _0574_;
	wire _0575_;
	wire _0576_;
	wire _0577_;
	wire _0578_;
	wire _0579_;
	wire _0580_;
	wire _0581_;
	wire _0582_;
	wire _0583_;
	wire _0584_;
	wire _0585_;
	wire _0586_;
	wire _0587_;
	wire _0588_;
	wire _0589_;
	wire _0590_;
	wire _0591_;
	wire _0592_;
	wire _0593_;
	wire _0594_;
	wire _0595_;
	wire _0596_;
	wire _0597_;
	wire _0598_;
	wire _0599_;
	wire _0600_;
	wire _0601_;
	wire _0602_;
	wire _0603_;
	wire _0604_;
	wire _0605_;
	wire _0606_;
	wire _0607_;
	wire _0608_;
	wire _0609_;
	wire _0610_;
	wire _0611_;
	wire _0612_;
	wire _0613_;
	wire _0614_;
	wire _0615_;
	wire _0616_;
	wire _0617_;
	wire _0618_;
	wire _0619_;
	wire _0620_;
	wire _0621_;
	wire _0622_;
	wire _0623_;
	wire _0624_;
	wire _0625_;
	wire _0626_;
	wire _0627_;
	wire _0628_;
	wire _0629_;
	wire _0630_;
	wire _0631_;
	wire _0632_;
	wire _0633_;
	wire _0634_;
	wire _0635_;
	wire _0636_;
	wire _0637_;
	wire _0638_;
	wire _0639_;
	wire _0640_;
	wire _0641_;
	wire _0642_;
	wire _0643_;
	wire _0644_;
	wire _0645_;
	wire _0646_;
	wire _0647_;
	wire _0648_;
	wire _0649_;
	wire _0650_;
	wire _0651_;
	wire _0652_;
	wire _0653_;
	wire _0654_;
	wire _0655_;
	wire _0656_;
	wire _0657_;
	wire _0658_;
	wire _0659_;
	wire _0660_;
	wire _0661_;
	wire _0662_;
	wire _0663_;
	wire _0664_;
	wire _0665_;
	wire _0666_;
	wire _0667_;
	wire _0668_;
	wire _0669_;
	wire _0670_;
	wire _0671_;
	wire _0672_;
	wire _0673_;
	wire _0674_;
	wire _0675_;
	wire _0676_;
	wire _0677_;
	wire _0678_;
	wire _0679_;
	wire _0680_;
	wire _0681_;
	wire _0682_;
	wire _0683_;
	wire _0684_;
	wire _0685_;
	wire _0686_;
	wire _0687_;
	wire _0688_;
	wire _0689_;
	wire _0690_;
	wire _0691_;
	wire _0692_;
	wire _0693_;
	wire _0694_;
	wire _0695_;
	wire _0696_;
	wire _0697_;
	wire _0698_;
	wire _0699_;
	wire _0700_;
	wire _0701_;
	wire _0702_;
	wire _0703_;
	wire _0704_;
	wire _0705_;
	wire _0706_;
	wire _0707_;
	wire _0708_;
	wire _0709_;
	wire _0710_;
	wire _0711_;
	wire _0712_;
	wire _0713_;
	wire _0714_;
	wire _0715_;
	wire _0716_;
	wire _0717_;
	wire _0718_;
	wire _0719_;
	wire _0720_;
	wire _0721_;
	wire _0722_;
	wire _0723_;
	wire _0724_;
	wire _0725_;
	wire _0726_;
	wire _0727_;
	wire _0728_;
	wire _0729_;
	wire _0730_;
	wire _0731_;
	wire _0732_;
	wire _0733_;
	wire _0734_;
	wire _0735_;
	wire _0736_;
	wire _0737_;
	wire _0738_;
	wire _0739_;
	wire _0740_;
	wire _0741_;
	wire _0742_;
	wire _0743_;
	wire _0744_;
	wire _0745_;
	wire _0746_;
	wire _0747_;
	wire _0748_;
	wire _0749_;
	wire _0750_;
	wire _0751_;
	wire _0752_;
	wire _0753_;
	wire _0754_;
	wire _0755_;
	wire _0756_;
	wire _0757_;
	wire _0758_;
	wire _0759_;
	wire _0760_;
	wire _0761_;
	wire _0762_;
	wire _0763_;
	wire _0764_;
	wire _0765_;
	wire _0766_;
	wire _0767_;
	wire _0768_;
	wire _0769_;
	wire _0770_;
	wire _0771_;
	wire _0772_;
	wire _0773_;
	wire _0774_;
	wire _0775_;
	wire _0776_;
	wire _0777_;
	wire _0778_;
	wire _0779_;
	wire _0780_;
	wire _0781_;
	wire _0782_;
	wire _0783_;
	wire _0784_;
	wire _0785_;
	wire _0786_;
	wire _0787_;
	wire _0788_;
	wire _0789_;
	wire _0790_;
	wire _0791_;
	wire _0792_;
	wire _0793_;
	wire _0794_;
	wire _0795_;
	wire _0796_;
	wire _0797_;
	wire _0798_;
	wire _0799_;
	wire _0800_;
	wire _0801_;
	wire _0802_;
	wire _0803_;
	wire _0804_;
	wire _0805_;
	wire _0806_;
	wire _0807_;
	wire _0808_;
	wire _0809_;
	wire _0810_;
	wire _0811_;
	wire _0812_;
	wire _0813_;
	wire _0814_;
	wire _0815_;
	wire _0816_;
	wire _0817_;
	wire _0818_;
	wire _0819_;
	wire _0820_;
	wire _0821_;
	wire _0822_;
	wire _0823_;
	wire _0824_;
	wire _0825_;
	wire _0826_;
	wire _0827_;
	wire _0828_;
	wire _0829_;
	wire _0830_;
	wire _0831_;
	wire _0832_;
	wire _0833_;
	wire _0834_;
	wire _0835_;
	wire _0836_;
	wire _0837_;
	wire _0838_;
	wire _0839_;
	wire _0840_;
	wire _0841_;
	wire _0842_;
	wire _0843_;
	wire _0844_;
	wire _0845_;
	wire _0846_;
	wire _0847_;
	wire _0848_;
	wire _0849_;
	wire _0850_;
	wire _0851_;
	wire _0852_;
	wire _0853_;
	wire _0854_;
	wire _0855_;
	wire _0856_;
	wire _0857_;
	wire _0858_;
	wire _0859_;
	wire _0860_;
	wire _0861_;
	wire _0862_;
	wire _0863_;
	wire _0864_;
	wire _0865_;
	wire _0866_;
	wire _0867_;
	wire _0868_;
	wire _0869_;
	wire _0870_;
	wire _0871_;
	wire _0872_;
	wire _0873_;
	wire _0874_;
	wire _0875_;
	wire _0876_;
	wire _0877_;
	wire _0878_;
	wire _0879_;
	wire _0880_;
	wire _0881_;
	wire _0882_;
	wire _0883_;
	wire _0884_;
	wire _0885_;
	wire _0886_;
	wire _0887_;
	wire _0888_;
	wire _0889_;
	wire _0890_;
	wire _0891_;
	wire _0892_;
	wire _0893_;
	wire _0894_;
	wire _0895_;
	wire _0896_;
	wire _0897_;
	wire _0898_;
	wire _0899_;
	wire _0900_;
	wire _0901_;
	wire _0902_;
	wire _0903_;
	wire _0904_;
	wire _0905_;
	wire _0906_;
	wire _0907_;
	wire _0908_;
	wire _0909_;
	wire _0910_;
	wire _0911_;
	wire _0912_;
	wire _0913_;
	wire _0914_;
	wire _0915_;
	wire _0916_;
	wire _0917_;
	wire _0918_;
	wire _0919_;
	wire _0920_;
	wire _0921_;
	wire _0922_;
	wire _0923_;
	wire _0924_;
	wire _0925_;
	wire _0926_;
	wire _0927_;
	wire _0928_;
	wire _0929_;
	wire _0930_;
	wire _0931_;
	wire _0932_;
	wire _0933_;
	wire _0934_;
	wire _0935_;
	wire _0936_;
	wire _0937_;
	wire _0938_;
	wire _0939_;
	wire _0940_;
	wire _0941_;
	wire _0942_;
	wire _0943_;
	wire _0944_;
	wire _0945_;
	wire _0946_;
	wire _0947_;
	wire _0948_;
	wire _0949_;
	wire _0950_;
	wire _0951_;
	wire _0952_;
	wire _0953_;
	wire _0954_;
	wire _0955_;
	wire _0956_;
	wire _0957_;
	wire _0958_;
	wire _0959_;
	wire _0960_;
	wire _0961_;
	wire _0962_;
	wire _0963_;
	wire _0964_;
	wire _0965_;
	wire _0966_;
	wire _0967_;
	wire _0968_;
	wire _0969_;
	wire _0970_;
	wire _0971_;
	wire _0972_;
	wire _0973_;
	wire _0974_;
	wire _0975_;
	wire _0976_;
	wire _0977_;
	wire _0978_;
	wire _0979_;
	wire _0980_;
	wire _0981_;
	wire _0982_;
	wire _0983_;
	wire _0984_;
	wire _0985_;
	wire _0986_;
	wire _0987_;
	wire _0988_;
	wire _0989_;
	wire _0990_;
	wire _0991_;
	wire _0992_;
	wire _0993_;
	wire _0994_;
	wire _0995_;
	wire _0996_;
	wire _0997_;
	wire _0998_;
	wire _0999_;
	wire _1000_;
	wire _1001_;
	wire _1002_;
	wire _1003_;
	wire _1004_;
	wire _1005_;
	wire _1006_;
	wire _1007_;
	wire _1008_;
	wire _1009_;
	wire _1010_;
	wire _1011_;
	wire _1012_;
	wire _1013_;
	wire _1014_;
	wire _1015_;
	wire _1016_;
	wire _1017_;
	wire _1018_;
	wire _1019_;
	wire _1020_;
	wire _1021_;
	wire _1022_;
	wire _1023_;
	wire _1024_;
	wire _1025_;
	wire _1026_;
	wire _1027_;
	wire _1028_;
	wire _1029_;
	wire _1030_;
	wire _1031_;
	wire _1032_;
	wire _1033_;
	wire _1034_;
	wire _1035_;
	wire _1036_;
	wire _1037_;
	wire _1038_;
	wire _1039_;
	wire _1040_;
	wire _1041_;
	wire _1042_;
	wire _1043_;
	wire _1044_;
	wire _1045_;
	wire _1046_;
	wire _1047_;
	wire _1048_;
	wire _1049_;
	wire _1050_;
	wire _1051_;
	wire _1052_;
	wire _1053_;
	wire _1054_;
	wire _1055_;
	wire _1056_;
	wire _1057_;
	wire _1058_;
	wire _1059_;
	wire _1060_;
	wire _1061_;
	wire _1062_;
	wire _1063_;
	wire _1064_;
	wire _1065_;
	wire _1066_;
	wire _1067_;
	wire _1068_;
	wire _1069_;
	wire _1070_;
	wire _1071_;
	wire _1072_;
	wire _1073_;
	wire _1074_;
	wire _1075_;
	wire _1076_;
	wire _1077_;
	wire _1078_;
	wire _1079_;
	wire _1080_;
	wire _1081_;
	wire _1082_;
	wire _1083_;
	wire _1084_;
	wire _1085_;
	wire _1086_;
	wire _1087_;
	wire _1088_;
	wire _1089_;
	wire _1090_;
	wire _1091_;
	wire _1092_;
	wire _1093_;
	wire _1094_;
	wire _1095_;
	wire _1096_;
	wire _1097_;
	wire _1098_;
	wire _1099_;
	wire _1100_;
	wire _1101_;
	wire _1102_;
	wire _1103_;
	wire _1104_;
	wire _1105_;
	wire _1106_;
	wire _1107_;
	wire _1108_;
	wire _1109_;
	wire _1110_;
	wire _1111_;
	wire _1112_;
	wire _1113_;
	wire _1114_;
	wire _1115_;
	wire _1116_;
	wire _1117_;
	wire _1118_;
	wire _1119_;
	wire _1120_;
	wire _1121_;
	wire _1122_;
	wire _1123_;
	wire _1124_;
	wire _1125_;
	wire _1126_;
	wire _1127_;
	wire _1128_;
	wire _1129_;
	wire _1130_;
	wire _1131_;
	wire _1132_;
	wire _1133_;
	wire _1134_;
	wire _1135_;
	wire _1136_;
	wire _1137_;
	wire _1138_;
	wire _1139_;
	wire _1140_;
	wire _1141_;
	wire _1142_;
	wire _1143_;
	wire _1144_;
	wire _1145_;
	wire _1146_;
	wire _1147_;
	wire _1148_;
	wire _1149_;
	wire _1150_;
	wire _1151_;
	wire _1152_;
	wire _1153_;
	wire _1154_;
	wire _1155_;
	wire _1156_;
	wire _1157_;
	wire _1158_;
	wire _1159_;
	wire _1160_;
	wire _1161_;
	wire _1162_;
	wire _1163_;
	wire _1164_;
	wire _1165_;
	wire _1166_;
	wire _1167_;
	wire _1168_;
	wire _1169_;
	wire _1170_;
	wire _1171_;
	wire _1172_;
	wire _1173_;
	wire _1174_;
	wire _1175_;
	wire _1176_;
	wire _1177_;
	wire _1178_;
	wire _1179_;
	wire _1180_;
	wire _1181_;
	wire _1182_;
	wire _1183_;
	wire _1184_;
	wire _1185_;
	wire _1186_;
	wire _1187_;
	wire _1188_;
	wire _1189_;
	wire _1190_;
	wire _1191_;
	wire _1192_;
	wire _1193_;
	wire _1194_;
	wire _1195_;
	wire _1196_;
	wire _1197_;
	wire _1198_;
	wire _1199_;
	wire _1200_;
	wire _1201_;
	wire _1202_;
	wire _1203_;
	wire _1204_;
	wire _1205_;
	wire _1206_;
	wire _1207_;
	wire _1208_;
	wire _1209_;
	wire _1210_;
	wire _1211_;
	wire _1212_;
	wire _1213_;
	wire _1214_;
	wire _1215_;
	wire _1216_;
	wire _1217_;
	wire _1218_;
	wire _1219_;
	wire _1220_;
	wire _1221_;
	wire _1222_;
	wire _1223_;
	wire _1224_;
	wire _1225_;
	wire _1226_;
	wire _1227_;
	wire _1228_;
	wire _1229_;
	wire _1230_;
	wire _1231_;
	wire _1232_;
	wire _1233_;
	wire _1234_;
	wire _1235_;
	wire _1236_;
	wire _1237_;
	wire _1238_;
	wire _1239_;
	wire _1240_;
	wire _1241_;
	wire _1242_;
	wire _1243_;
	wire _1244_;
	wire _1245_;
	wire _1246_;
	wire _1247_;
	wire _1248_;
	wire _1249_;
	wire _1250_;
	wire _1251_;
	wire _1252_;
	wire _1253_;
	wire _1254_;
	wire _1255_;
	wire _1256_;
	wire _1257_;
	wire _1258_;
	wire _1259_;
	wire _1260_;
	wire _1261_;
	wire _1262_;
	wire _1263_;
	wire _1264_;
	wire _1265_;
	wire _1266_;
	wire _1267_;
	wire _1268_;
	wire _1269_;
	wire _1270_;
	wire _1271_;
	wire _1272_;
	wire _1273_;
	wire _1274_;
	wire _1275_;
	wire _1276_;
	wire _1277_;
	wire _1278_;
	wire _1279_;
	wire _1280_;
	wire _1281_;
	wire _1282_;
	wire _1283_;
	wire _1284_;
	wire _1285_;
	wire _1286_;
	wire _1287_;
	wire _1288_;
	wire _1289_;
	wire _1290_;
	wire _1291_;
	wire _1292_;
	wire _1293_;
	wire _1294_;
	wire _1295_;
	wire _1296_;
	wire _1297_;
	wire _1298_;
	wire _1299_;
	wire _1300_;
	wire _1301_;
	wire _1302_;
	wire _1303_;
	wire _1304_;
	wire _1305_;
	wire _1306_;
	wire _1307_;
	wire _1308_;
	wire _1309_;
	wire _1310_;
	wire _1311_;
	wire _1312_;
	wire _1313_;
	wire _1314_;
	wire _1315_;
	wire _1316_;
	wire _1317_;
	wire _1318_;
	wire _1319_;
	wire _1320_;
	wire _1321_;
	wire _1322_;
	wire _1323_;
	wire _1324_;
	wire _1325_;
	wire _1326_;
	wire _1327_;
	wire _1328_;
	wire _1329_;
	wire _1330_;
	wire _1331_;
	wire _1332_;
	wire _1333_;
	wire _1334_;
	wire _1335_;
	wire _1336_;
	wire _1337_;
	wire _1338_;
	wire _1339_;
	wire _1340_;
	wire _1341_;
	wire _1342_;
	wire _1343_;
	wire _1344_;
	wire _1345_;
	wire _1346_;
	wire _1347_;
	wire _1348_;
	wire _1349_;
	wire _1350_;
	wire _1351_;
	wire _1352_;
	wire _1353_;
	wire _1354_;
	wire _1355_;
	wire _1356_;
	wire _1357_;
	wire _1358_;
	wire _1359_;
	wire _1360_;
	wire _1361_;
	wire _1362_;
	wire _1363_;
	wire _1364_;
	wire _1365_;
	wire _1366_;
	wire _1367_;
	wire _1368_;
	wire _1369_;
	wire _1370_;
	wire _1371_;
	wire _1372_;
	wire _1373_;
	wire _1374_;
	wire _1375_;
	wire _1376_;
	wire _1377_;
	wire _1378_;
	wire _1379_;
	wire _1380_;
	wire _1381_;
	wire _1382_;
	wire _1383_;
	wire _1384_;
	wire _1385_;
	wire _1386_;
	wire _1387_;
	wire _1388_;
	wire _1389_;
	wire _1390_;
	wire _1391_;
	wire _1392_;
	wire _1393_;
	wire _1394_;
	wire _1395_;
	wire _1396_;
	wire _1397_;
	wire _1398_;
	wire _1399_;
	wire _1400_;
	wire _1401_;
	wire _1402_;
	wire _1403_;
	wire _1404_;
	wire _1405_;
	wire _1406_;
	wire _1407_;
	wire _1408_;
	wire _1409_;
	wire _1410_;
	wire _1411_;
	wire _1412_;
	wire _1413_;
	wire _1414_;
	wire _1415_;
	wire _1416_;
	wire _1417_;
	wire _1418_;
	wire _1419_;
	wire _1420_;
	wire _1421_;
	wire _1422_;
	wire _1423_;
	wire _1424_;
	wire _1425_;
	wire _1426_;
	wire _1427_;
	wire _1428_;
	wire _1429_;
	wire _1430_;
	wire _1431_;
	wire _1432_;
	wire _1433_;
	wire _1434_;
	wire _1435_;
	wire _1436_;
	wire _1437_;
	wire _1438_;
	wire _1439_;
	wire _1440_;
	wire _1441_;
	wire _1442_;
	wire _1443_;
	wire _1444_;
	wire _1445_;
	wire _1446_;
	wire _1447_;
	wire _1448_;
	wire _1449_;
	wire _1450_;
	wire _1451_;
	wire _1452_;
	wire _1453_;
	wire _1454_;
	wire _1455_;
	wire _1456_;
	wire _1457_;
	wire _1458_;
	wire _1459_;
	wire _1460_;
	wire _1461_;
	wire _1462_;
	wire _1463_;
	wire _1464_;
	wire _1465_;
	wire _1466_;
	wire _1467_;
	wire _1468_;
	wire _1469_;
	wire _1470_;
	wire _1471_;
	wire _1472_;
	wire _1473_;
	wire _1474_;
	wire _1475_;
	wire _1476_;
	wire _1477_;
	wire _1478_;
	wire _1479_;
	wire _1480_;
	wire _1481_;
	wire _1482_;
	wire _1483_;
	wire _1484_;
	wire _1485_;
	wire _1486_;
	wire _1487_;
	wire _1488_;
	wire _1489_;
	wire _1490_;
	wire _1491_;
	wire _1492_;
	wire _1493_;
	wire _1494_;
	wire _1495_;
	wire _1496_;
	wire _1497_;
	wire _1498_;
	wire _1499_;
	wire _1500_;
	wire _1501_;
	wire _1502_;
	wire _1503_;
	wire _1504_;
	wire _1505_;
	wire _1506_;
	wire _1507_;
	wire _1508_;
	wire _1509_;
	wire _1510_;
	wire _1511_;
	wire _1512_;
	wire _1513_;
	wire _1514_;
	wire _1515_;
	wire _1516_;
	wire _1517_;
	wire _1518_;
	wire _1519_;
	wire _1520_;
	wire _1521_;
	wire _1522_;
	wire _1523_;
	wire _1524_;
	wire _1525_;
	wire _1526_;
	wire _1527_;
	wire _1528_;
	wire _1529_;
	wire _1530_;
	wire _1531_;
	wire _1532_;
	wire _1533_;
	wire _1534_;
	wire _1535_;
	wire _1536_;
	wire _1537_;
	wire _1538_;
	wire _1539_;
	wire _1540_;
	wire _1541_;
	wire _1542_;
	wire _1543_;
	wire _1544_;
	wire _1545_;
	wire _1546_;
	wire _1547_;
	wire _1548_;
	wire _1549_;
	wire _1550_;
	wire _1551_;
	wire _1552_;
	wire _1553_;
	wire _1554_;
	wire _1555_;
	wire _1556_;
	wire _1557_;
	wire _1558_;
	wire _1559_;
	wire _1560_;
	wire _1561_;
	wire _1562_;
	wire _1563_;
	wire _1564_;
	wire _1565_;
	wire _1566_;
	wire _1567_;
	wire _1568_;
	wire _1569_;
	wire _1570_;
	wire _1571_;
	wire _1572_;
	wire _1573_;
	wire _1574_;
	wire _1575_;
	wire _1576_;
	wire _1577_;
	wire _1578_;
	wire _1579_;
	wire _1580_;
	wire _1581_;
	wire _1582_;
	wire _1583_;
	wire _1584_;
	wire _1585_;
	wire _1586_;
	wire _1587_;
	wire _1588_;
	wire _1589_;
	wire _1590_;
	wire _1591_;
	wire _1592_;
	wire _1593_;
	wire _1594_;
	wire _1595_;
	wire _1596_;
	wire _1597_;
	wire _1598_;
	wire _1599_;
	wire _1600_;
	wire _1601_;
	wire _1602_;
	wire _1603_;
	wire _1604_;
	wire _1605_;
	wire _1606_;
	wire _1607_;
	wire _1608_;
	wire _1609_;
	wire _1610_;
	wire _1611_;
	wire _1612_;
	wire _1613_;
	wire _1614_;
	wire _1615_;
	wire _1616_;
	wire _1617_;
	wire _1618_;
	wire _1619_;
	wire _1620_;
	wire _1621_;
	wire _1622_;
	wire _1623_;
	wire _1624_;
	wire _1625_;
	wire _1626_;
	wire _1627_;
	wire _1628_;
	wire _1629_;
	wire _1630_;
	wire _1631_;
	wire _1632_;
	wire _1633_;
	wire _1634_;
	wire _1635_;
	wire _1636_;
	wire _1637_;
	wire _1638_;
	wire _1639_;
	wire _1640_;
	wire _1641_;
	wire _1642_;
	wire _1643_;
	wire _1644_;
	wire _1645_;
	wire _1646_;
	wire _1647_;
	wire _1648_;
	wire _1649_;
	wire _1650_;
	wire _1651_;
	wire _1652_;
	wire _1653_;
	wire _1654_;
	wire _1655_;
	wire _1656_;
	wire _1657_;
	wire _1658_;
	wire _1659_;
	wire _1660_;
	wire _1661_;
	wire _1662_;
	wire _1663_;
	wire _1664_;
	wire _1665_;
	wire _1666_;
	wire _1667_;
	wire _1668_;
	wire _1669_;
	wire _1670_;
	wire _1671_;
	wire _1672_;
	wire _1673_;
	wire _1674_;
	wire _1675_;
	wire _1676_;
	wire _1677_;
	wire _1678_;
	wire _1679_;
	wire _1680_;
	wire _1681_;
	wire _1682_;
	wire _1683_;
	wire _1684_;
	wire _1685_;
	wire _1686_;
	wire _1687_;
	wire _1688_;
	wire _1689_;
	wire _1690_;
	wire _1691_;
	wire _1692_;
	wire _1693_;
	wire _1694_;
	wire _1695_;
	wire _1696_;
	wire _1697_;
	wire _1698_;
	wire _1699_;
	wire _1700_;
	wire _1701_;
	wire _1702_;
	wire _1703_;
	wire _1704_;
	wire _1705_;
	wire _1706_;
	wire _1707_;
	wire _1708_;
	wire _1709_;
	wire _1710_;
	wire _1711_;
	wire _1712_;
	wire _1713_;
	wire _1714_;
	wire _1715_;
	wire _1716_;
	wire _1717_;
	wire _1718_;
	wire _1719_;
	wire _1720_;
	wire _1721_;
	wire _1722_;
	wire _1723_;
	wire _1724_;
	wire _1725_;
	wire _1726_;
	wire _1727_;
	wire _1728_;
	wire _1729_;
	wire _1730_;
	wire _1731_;
	wire _1732_;
	wire _1733_;
	wire _1734_;
	wire _1735_;
	wire _1736_;
	wire _1737_;
	wire _1738_;
	wire _1739_;
	wire _1740_;
	wire _1741_;
	wire _1742_;
	wire _1743_;
	wire _1744_;
	wire _1745_;
	wire _1746_;
	wire _1747_;
	wire _1748_;
	wire _1749_;
	wire _1750_;
	wire _1751_;
	wire _1752_;
	wire _1753_;
	wire _1754_;
	wire _1755_;
	wire _1756_;
	wire _1757_;
	wire _1758_;
	wire _1759_;
	wire _1760_;
	wire _1761_;
	wire _1762_;
	wire _1763_;
	wire _1764_;
	wire _1765_;
	wire _1766_;
	wire _1767_;
	wire _1768_;
	wire _1769_;
	wire _1770_;
	wire _1771_;
	wire _1772_;
	wire _1773_;
	wire _1774_;
	wire _1775_;
	wire _1776_;
	wire _1777_;
	wire _1778_;
	wire _1779_;
	wire _1780_;
	wire _1781_;
	wire _1782_;
	wire _1783_;
	wire _1784_;
	wire _1785_;
	wire _1786_;
	wire _1787_;
	wire _1788_;
	wire _1789_;
	wire _1790_;
	wire _1791_;
	wire _1792_;
	wire _1793_;
	wire _1794_;
	wire _1795_;
	wire _1796_;
	wire _1797_;
	wire _1798_;
	wire _1799_;
	wire _1800_;
	wire _1801_;
	wire _1802_;
	wire _1803_;
	wire _1804_;
	wire _1805_;
	wire _1806_;
	wire _1807_;
	wire _1808_;
	wire _1809_;
	wire _1810_;
	wire _1811_;
	wire _1812_;
	wire _1813_;
	wire _1814_;
	wire _1815_;
	wire _1816_;
	wire _1817_;
	wire _1818_;
	wire _1819_;
	wire _1820_;
	wire _1821_;
	wire _1822_;
	wire _1823_;
	wire _1824_;
	wire _1825_;
	wire _1826_;
	wire _1827_;
	wire _1828_;
	wire _1829_;
	wire _1830_;
	wire _1831_;
	wire _1832_;
	wire _1833_;
	wire _1834_;
	wire _1835_;
	wire _1836_;
	wire _1837_;
	wire _1838_;
	wire _1839_;
	wire _1840_;
	wire _1841_;
	wire _1842_;
	wire _1843_;
	wire _1844_;
	wire _1845_;
	wire _1846_;
	wire _1847_;
	wire _1848_;
	wire _1849_;
	wire _1850_;
	wire _1851_;
	wire _1852_;
	wire _1853_;
	wire _1854_;
	wire _1855_;
	wire _1856_;
	wire _1857_;
	wire _1858_;
	wire _1859_;
	wire _1860_;
	wire _1861_;
	wire _1862_;
	wire _1863_;
	wire _1864_;
	wire _1865_;
	wire _1866_;
	wire _1867_;
	wire _1868_;
	wire _1869_;
	wire _1870_;
	wire _1871_;
	wire _1872_;
	wire _1873_;
	wire _1874_;
	wire _1875_;
	wire _1876_;
	wire _1877_;
	wire _1878_;
	wire _1879_;
	wire _1880_;
	wire _1881_;
	wire _1882_;
	wire _1883_;
	wire _1884_;
	wire _1885_;
	wire _1886_;
	wire _1887_;
	wire _1888_;
	wire _1889_;
	wire _1890_;
	wire _1891_;
	wire _1892_;
	wire _1893_;
	wire _1894_;
	wire _1895_;
	wire _1896_;
	wire _1897_;
	wire _1898_;
	wire _1899_;
	wire _1900_;
	wire _1901_;
	wire _1902_;
	wire _1903_;
	wire _1904_;
	wire _1905_;
	wire _1906_;
	wire _1907_;
	wire _1908_;
	wire _1909_;
	wire _1910_;
	wire _1911_;
	wire _1912_;
	wire _1913_;
	wire _1914_;
	wire _1915_;
	wire _1916_;
	wire _1917_;
	wire _1918_;
	wire _1919_;
	wire _1920_;
	wire _1921_;
	wire _1922_;
	wire _1923_;
	wire _1924_;
	wire _1925_;
	wire _1926_;
	wire _1927_;
	wire _1928_;
	wire _1929_;
	wire _1930_;
	wire _1931_;
	wire _1932_;
	wire _1933_;
	wire _1934_;
	wire _1935_;
	wire _1936_;
	wire _1937_;
	wire _1938_;
	wire _1939_;
	wire _1940_;
	wire _1941_;
	wire _1942_;
	wire _1943_;
	wire _1944_;
	wire _1945_;
	wire _1946_;
	wire _1947_;
	wire _1948_;
	wire _1949_;
	wire _1950_;
	wire _1951_;
	wire _1952_;
	wire _1953_;
	wire _1954_;
	wire _1955_;
	wire _1956_;
	wire _1957_;
	wire _1958_;
	wire _1959_;
	wire _1960_;
	wire _1961_;
	wire _1962_;
	wire _1963_;
	wire _1964_;
	wire _1965_;
	wire _1966_;
	wire _1967_;
	wire _1968_;
	wire _1969_;
	wire _1970_;
	wire _1971_;
	wire _1972_;
	wire _1973_;
	wire _1974_;
	wire _1975_;
	wire _1976_;
	wire _1977_;
	wire _1978_;
	wire _1979_;
	wire _1980_;
	wire _1981_;
	wire _1982_;
	wire _1983_;
	wire _1984_;
	wire _1985_;
	wire _1986_;
	wire _1987_;
	wire _1988_;
	wire _1989_;
	wire _1990_;
	wire _1991_;
	wire _1992_;
	wire _1993_;
	wire _1994_;
	wire _1995_;
	wire _1996_;
	wire _1997_;
	wire _1998_;
	wire _1999_;
	wire _2000_;
	wire _2001_;
	wire _2002_;
	wire _2003_;
	wire _2004_;
	wire _2005_;
	wire _2006_;
	wire _2007_;
	wire _2008_;
	wire _2009_;
	wire _2010_;
	wire _2011_;
	wire _2012_;
	wire _2013_;
	wire _2014_;
	wire _2015_;
	wire _2016_;
	wire _2017_;
	wire _2018_;
	wire _2019_;
	wire _2020_;
	wire _2021_;
	wire _2022_;
	wire _2023_;
	wire _2024_;
	wire _2025_;
	wire _2026_;
	wire _2027_;
	wire _2028_;
	wire _2029_;
	wire _2030_;
	wire _2031_;
	wire _2032_;
	wire _2033_;
	wire _2034_;
	wire _2035_;
	wire _2036_;
	wire _2037_;
	wire _2038_;
	wire _2039_;
	wire _2040_;
	wire _2041_;
	wire _2042_;
	wire _2043_;
	wire _2044_;
	wire _2045_;
	wire _2046_;
	wire _2047_;
	wire _2048_;
	wire _2049_;
	wire _2050_;
	wire _2051_;
	wire _2052_;
	wire _2053_;
	wire _2054_;
	wire _2055_;
	wire _2056_;
	wire _2057_;
	wire _2058_;
	wire _2059_;
	wire _2060_;
	wire _2061_;
	wire _2062_;
	wire _2063_;
	wire _2064_;
	wire _2065_;
	wire _2066_;
	wire _2067_;
	wire _2068_;
	wire _2069_;
	wire _2070_;
	wire _2071_;
	wire _2072_;
	wire _2073_;
	wire _2074_;
	wire _2075_;
	wire _2076_;
	wire _2077_;
	wire _2078_;
	wire _2079_;
	wire _2080_;
	wire _2081_;
	wire _2082_;
	wire _2083_;
	wire _2084_;
	wire _2085_;
	wire _2086_;
	wire _2087_;
	wire _2088_;
	wire _2089_;
	wire _2090_;
	wire _2091_;
	wire _2092_;
	wire _2093_;
	wire _2094_;
	wire _2095_;
	wire _2096_;
	wire _2097_;
	wire _2098_;
	wire _2099_;
	wire _2100_;
	wire _2101_;
	wire _2102_;
	wire _2103_;
	wire _2104_;
	wire _2105_;
	wire _2106_;
	wire _2107_;
	wire _2108_;
	wire _2109_;
	wire _2110_;
	wire _2111_;
	wire _2112_;
	wire _2113_;
	wire _2114_;
	wire _2115_;
	wire _2116_;
	wire _2117_;
	wire _2118_;
	wire _2119_;
	wire _2120_;
	wire _2121_;
	wire _2122_;
	wire _2123_;
	wire _2124_;
	wire _2125_;
	wire _2126_;
	wire _2127_;
	wire _2128_;
	wire _2129_;
	wire _2130_;
	wire _2131_;
	wire _2132_;
	wire _2133_;
	wire _2134_;
	wire _2135_;
	wire _2136_;
	wire _2137_;
	wire _2138_;
	wire _2139_;
	wire _2140_;
	wire _2141_;
	wire _2142_;
	wire _2143_;
	wire _2144_;
	wire _2145_;
	wire _2146_;
	wire _2147_;
	wire _2148_;
	wire _2149_;
	wire _2150_;
	wire _2151_;
	wire _2152_;
	wire _2153_;
	wire _2154_;
	wire _2155_;
	wire _2156_;
	wire _2157_;
	wire _2158_;
	wire _2159_;
	wire _2160_;
	wire _2161_;
	wire _2162_;
	wire _2163_;
	wire _2164_;
	wire _2165_;
	wire _2166_;
	wire _2167_;
	wire _2168_;
	wire _2169_;
	wire _2170_;
	wire _2171_;
	wire _2172_;
	wire _2173_;
	wire _2174_;
	wire _2175_;
	wire _2176_;
	wire _2177_;
	wire _2178_;
	wire _2179_;
	wire _2180_;
	wire _2181_;
	wire [6:0] _2182_;
	wire [6:0] _2183_;
	wire [3:0] _2184_;
	wire [3:0] _2185_;
	input wire [13:0] io_in;
	output wire [13:0] io_out;
	wire \mchip.clk ;
	wire \mchip.clock ;
	wire [127:0] \mchip.fallen_state ;
	wire [6:0] \mchip.idx ;
	wire [11:0] \mchip.io_in ;
	wire [11:0] \mchip.io_out ;
	wire [7:0] \mchip.iout ;
	wire \mchip.left ;
	wire [15:0] \mchip.rand_piece ;
	wire \mchip.read_gs ;
	wire \mchip.reset ;
	wire \mchip.right ;
	reg [6:0] \mchip.x ;
	wire [6:0] \mchip.y ;
	assign _0001_ = io_in[0] & ~io_in[13];
	assign _0000_ = io_in[1] | io_in[2];
	assign _1639_ = io_in[2] & ~\mchip.x [0];
	assign _1650_ = ~(\mchip.x [0] | io_in[2]);
	assign _0002_ = _1650_ | _1639_;
	assign _1670_ = ~io_in[2];
	assign _1681_ = ~(\mchip.x [1] | \mchip.x [0]);
	assign _0033_ = ~(\mchip.x [1] & \mchip.x [0]);
	assign _1697_ = _0033_ & ~_1681_;
	assign _0003_ = _1697_ ^ _1670_;
	assign _1717_ = ~\mchip.x [2];
	assign _1728_ = _1681_ ^ _1717_;
	assign _1739_ = ~_1728_;
	assign _1750_ = _0033_ ^ _1717_;
	assign _0004_ = (io_in[2] ? _1750_ : _1739_);
	assign _1771_ = _1681_ & ~\mchip.x [2];
	assign _1782_ = _1771_ ^ \mchip.x [3];
	assign _0384_ = \mchip.x [2] & ~_0033_;
	assign _1803_ = ~(_0384_ ^ \mchip.x [3]);
	assign _1814_ = ~_1803_;
	assign _0005_ = (io_in[2] ? _1814_ : _1782_);
	assign _1835_ = \mchip.x [3] | \mchip.x [2];
	assign _1846_ = _1681_ & ~_1835_;
	assign _1857_ = _1846_ ^ \mchip.x [4];
	assign _1868_ = ~(\mchip.x [3] & \mchip.x [2]);
	assign _1879_ = ~(_1868_ | _0033_);
	assign _1890_ = _1879_ ^ \mchip.x [4];
	assign _0006_ = (io_in[2] ? _1890_ : _1857_);
	assign _1911_ = _1846_ & ~\mchip.x [4];
	assign _1922_ = _1911_ ^ \mchip.x [5];
	assign _1933_ = ~\mchip.x [4];
	assign _1943_ = _1879_ & ~_1933_;
	assign _1953_ = _1943_ ^ \mchip.x [5];
	assign _0007_ = (io_in[2] ? _1953_ : _1922_);
	assign _1970_ = \mchip.x [5] | \mchip.x [4];
	assign _1981_ = _1846_ & ~_1970_;
	assign _1991_ = _1981_ ^ \mchip.x [6];
	assign _2002_ = ~\mchip.x [6];
	assign _2013_ = ~(\mchip.x [5] & \mchip.x [4]);
	assign _2024_ = _1879_ & ~_2013_;
	assign _2035_ = _2024_ ^ _2002_;
	assign _2046_ = ~_2035_;
	assign _0008_ = (io_in[2] ? _2046_ : _1991_);
	assign _2184_[0] = ~\mchip.idx [3];
	assign _2182_[0] = ~\mchip.y [0];
	assign _2185_[1] = \mchip.idx [4] ^ \mchip.idx [3];
	assign _2097_ = \mchip.idx [4] & \mchip.idx [3];
	assign _2185_[2] = _2097_ ^ \mchip.idx [5];
	assign _2118_ = ~\mchip.idx [5];
	assign _2129_ = _2097_ & ~_2118_;
	assign _2185_[3] = _2129_ ^ \mchip.idx [6];
	assign _2183_[1] = \mchip.y [1] ^ \mchip.y [0];
	assign _2160_ = \mchip.y [1] & \mchip.y [0];
	assign _2183_[2] = _2160_ ^ \mchip.y [2];
	assign _2181_ = ~(_2160_ & \mchip.y [2]);
	assign _2183_[3] = ~(_2181_ ^ \mchip.y [3]);
	assign _0048_ = \mchip.y [1] | ~_1890_;
	assign _0056_ = _1803_ | _2182_[0];
	assign _0067_ = _1890_ ^ \mchip.y [1];
	assign _0077_ = ~(_0067_ | _0056_);
	assign _0088_ = _0048_ & ~_0077_;
	assign _0099_ = \mchip.y [2] ^ \mchip.y [1];
	assign _0110_ = ~_0099_;
	assign _0121_ = _0110_ ^ _1953_;
	assign _0132_ = _0121_ | _0088_;
	assign _0143_ = _1953_ & ~_0110_;
	assign _0154_ = _0132_ & ~_0143_;
	assign _0165_ = \mchip.y [2] & \mchip.y [1];
	assign _0176_ = _0165_ ^ \mchip.y [3];
	assign _0187_ = _0176_ ^ _2035_;
	assign _0198_ = _0187_ ^ _0154_;
	assign _0209_ = _0121_ ^ _0088_;
	assign _0220_ = _0067_ ^ _0056_;
	assign _0231_ = _0220_ | _0209_;
	assign _0242_ = _1803_ ^ _2182_[0];
	assign _0253_ = _0242_ | _1750_;
	assign _0264_ = _0253_ | _0033_;
	assign _0275_ = ~(_0264_ | _0231_);
	assign _0286_ = _0198_ | ~_0275_;
	assign _0297_ = _0231_ | _0198_;
	assign _0307_ = ~(_0297_ | _0264_);
	assign _0318_ = ~(_0307_ & \mchip.x [0]);
	assign _0329_ = ~\mchip.x [0];
	assign _0340_ = _1697_ ^ _0329_;
	assign _0351_ = _0340_ | _0318_;
	assign _0362_ = _1750_ ^ _0033_;
	assign _0373_ = _0362_ | _0351_;
	assign _0395_ = ~(_0384_ ^ _0242_);
	assign _0406_ = _0395_ | _0373_;
	assign _0417_ = _0264_ ^ _0220_;
	assign _0428_ = _0417_ | _0406_;
	assign _0439_ = ~(_0264_ | _0220_);
	assign _0450_ = ~(_0439_ ^ _0209_);
	assign _0461_ = _0450_ | _0428_;
	assign _0472_ = _0198_ & ~_0275_;
	assign _0483_ = ~(_0461_ | _0286_);
	assign _0494_ = \mchip.x [4] & ~\mchip.y [1];
	assign _0505_ = \mchip.y [0] & \mchip.x [3];
	assign _0516_ = \mchip.y [1] ^ \mchip.x [4];
	assign _0527_ = _0505_ & ~_0516_;
	assign _0538_ = _0527_ | _0494_;
	assign _0549_ = ~\mchip.x [5];
	assign _0560_ = _0099_ ^ _0549_;
	assign _0571_ = _0538_ & ~_0560_;
	assign _0581_ = _0099_ & ~_0549_;
	assign _0591_ = _0581_ | _0571_;
	assign _0600_ = _0176_ ^ \mchip.x [6];
	assign _0611_ = _0600_ ^ _0591_;
	assign _0621_ = ~_1681_;
	assign _0632_ = \mchip.y [0] ^ \mchip.x [3];
	assign _0643_ = _0632_ | \mchip.x [2];
	assign _0654_ = ~(_0643_ | _0621_);
	assign _0665_ = ~(_0560_ ^ _0538_);
	assign _0676_ = _0516_ ^ _0505_;
	assign _0687_ = ~_0676_;
	assign _0698_ = _0687_ | _0665_;
	assign _0709_ = _0654_ & ~_0698_;
	assign _0720_ = _0611_ | ~_0709_;
	assign _0731_ = ~(_0632_ ^ _1771_);
	assign _0742_ = ~(_0698_ | _0611_);
	assign _0753_ = _0742_ & _0654_;
	assign _0764_ = ~(_0753_ & _0329_);
	assign _0775_ = _0764_ | _1697_;
	assign _0786_ = _0775_ | _1728_;
	assign _0797_ = _0786_ | _0731_;
	assign _0808_ = _0676_ ^ _0654_;
	assign _0819_ = _0808_ | _0797_;
	assign _0830_ = _0654_ & ~_0687_;
	assign _0841_ = ~(_0830_ ^ _0665_);
	assign _0851_ = _0841_ | _0819_;
	assign _0861_ = _0611_ & ~_0709_;
	assign _0870_ = ~(_0851_ | _0720_);
	assign _0881_ = _0870_ | _0483_;
	assign _0891_ = ~(_2183_[1] & \mchip.x [4]);
	assign _0902_ = \mchip.x [3] & ~\mchip.y [0];
	assign _0913_ = _2183_[1] ^ _1933_;
	assign _0924_ = _0902_ & ~_0913_;
	assign _0935_ = _0891_ & ~_0924_;
	assign _0946_ = _2183_[2] ^ _0549_;
	assign _0957_ = _0946_ | _0935_;
	assign _0968_ = _2183_[2] & ~_0549_;
	assign _0979_ = _0957_ & ~_0968_;
	assign _0990_ = _2183_[3] ^ _2002_;
	assign _1001_ = _0990_ ^ _0979_;
	assign _1012_ = _0946_ ^ _0935_;
	assign _1023_ = ~(_0913_ ^ _0902_);
	assign _1034_ = _1023_ | _1012_;
	assign _1045_ = ~(\mchip.y [0] ^ \mchip.x [3]);
	assign _1056_ = _1045_ | \mchip.x [2];
	assign _1067_ = _1056_ | _0621_;
	assign _1078_ = ~(_1067_ | _1034_);
	assign _1089_ = _1001_ | ~_1078_;
	assign _1100_ = _1034_ | _1001_;
	assign _1111_ = ~(_1100_ | _1067_);
	assign _1121_ = ~(_1111_ & _0329_);
	assign _1131_ = _1121_ | _1697_;
	assign _1140_ = _1131_ | _1728_;
	assign _1151_ = ~(_1045_ ^ _1771_);
	assign _1161_ = _1151_ | _1140_;
	assign _1172_ = _1067_ ^ _1023_;
	assign _1183_ = _1172_ | _1161_;
	assign _1194_ = ~(_1067_ | _1023_);
	assign _1205_ = ~(_1194_ ^ _1012_);
	assign _1216_ = _1205_ | _1183_;
	assign _1227_ = _1001_ & ~_1078_;
	assign _1238_ = ~(_1216_ | _1089_);
	assign _1249_ = _1238_ | _0881_;
	assign _1260_ = \mchip.y [2] & \mchip.x [5];
	assign _1271_ = \mchip.y [1] & \mchip.x [4];
	assign _1292_ = _0516_ & _0505_;
	assign _1303_ = _1292_ | _1271_;
	assign _1314_ = \mchip.y [2] ^ \mchip.x [5];
	assign _1325_ = _1314_ & _1303_;
	assign _1336_ = _1325_ | _1260_;
	assign _1347_ = \mchip.y [3] ^ \mchip.x [6];
	assign _1358_ = _1347_ ^ _1336_;
	assign _1369_ = _1314_ ^ _1303_;
	assign _1380_ = ~(_0516_ ^ _0505_);
	assign _1386_ = ~_1380_;
	assign _1387_ = _1386_ | _1369_;
	assign _1388_ = _0654_ & ~_1387_;
	assign _1389_ = _1358_ | ~_1388_;
	assign _1390_ = ~(_1387_ | _1358_);
	assign _1391_ = _1390_ & _0654_;
	assign _1392_ = ~(_1391_ & _0329_);
	assign _1393_ = _1392_ | _1697_;
	assign _1394_ = _1393_ | _1728_;
	assign _1395_ = _1394_ | _0731_;
	assign _1396_ = _1380_ ^ _0654_;
	assign _1397_ = _1396_ | _1395_;
	assign _1398_ = _0654_ & ~_1386_;
	assign _1399_ = ~(_1398_ ^ _1369_);
	assign _1400_ = _1399_ | _1397_;
	assign _1401_ = _1358_ & ~_1388_;
	assign _1402_ = ~(_1400_ | _1389_);
	assign _1403_ = _1402_ | _1249_;
	assign _1404_ = _0286_ & ~_0472_;
	assign _1405_ = ~_1404_;
	assign _1406_ = ~_0450_;
	assign _1407_ = ~_0417_;
	assign _1408_ = _0307_ | _0329_;
	assign _1409_ = _1408_ | _0340_;
	assign _1410_ = _1409_ | _0362_;
	assign _1411_ = _1410_ | ~_0395_;
	assign _1412_ = _1411_ | _1407_;
	assign _1413_ = _1412_ | _1406_;
	assign _1414_ = _1413_ | _1405_;
	assign _1415_ = _0286_ & ~_1414_;
	assign _1416_ = _0720_ & ~_0861_;
	assign _1417_ = ~_1416_;
	assign _1418_ = ~_0841_;
	assign _1419_ = ~_0808_;
	assign _1420_ = ~_0731_;
	assign _1421_ = _0753_ | \mchip.x [0];
	assign _1422_ = _1421_ | _1697_;
	assign _1423_ = _1422_ | _1728_;
	assign _1424_ = _1423_ | _1420_;
	assign _1425_ = _1424_ | _1419_;
	assign _1426_ = _1425_ | _1418_;
	assign _1427_ = _1426_ | _1417_;
	assign _1428_ = _0720_ & ~_1427_;
	assign _1429_ = _1428_ | _1415_;
	assign _1430_ = _1089_ & ~_1227_;
	assign _1431_ = ~_1430_;
	assign _1432_ = ~_1205_;
	assign _1433_ = ~_1172_;
	assign _1434_ = _1111_ | \mchip.x [0];
	assign _1435_ = _1434_ | _1697_;
	assign _1436_ = _1435_ | _1728_;
	assign _1437_ = _1436_ | ~_1151_;
	assign _1438_ = _1437_ | _1433_;
	assign _1439_ = _1438_ | _1432_;
	assign _1440_ = _1439_ | _1431_;
	assign _1441_ = _1089_ & ~_1440_;
	assign _1442_ = _1441_ | _1429_;
	assign _1443_ = _1389_ & ~_1401_;
	assign _1444_ = ~_1443_;
	assign _1445_ = ~_1399_;
	assign _1446_ = ~_1396_;
	assign _1447_ = _1391_ | \mchip.x [0];
	assign _1448_ = _1447_ | _1697_;
	assign _1449_ = _1448_ | _1728_;
	assign _1450_ = _1449_ | _1420_;
	assign _1451_ = _1450_ | _1446_;
	assign _1452_ = _1451_ | _1445_;
	assign _1453_ = _1452_ | _1444_;
	assign _1454_ = _1389_ & ~_1453_;
	assign _1455_ = _1454_ | _1442_;
	assign _1456_ = (\mchip.idx [3] ? _1455_ : _1403_);
	assign _1457_ = _1410_ | _0395_;
	assign _1458_ = _1457_ | _1407_;
	assign _1459_ = _1458_ | _1406_;
	assign _1460_ = _1459_ | _1405_;
	assign _1461_ = _0286_ & ~_1460_;
	assign _1462_ = _1423_ | _0731_;
	assign _1463_ = _1462_ | _1419_;
	assign _1464_ = _1463_ | _1418_;
	assign _1465_ = _1464_ | _1417_;
	assign _1466_ = _0720_ & ~_1465_;
	assign _1467_ = _1466_ | _1461_;
	assign _1468_ = _1436_ | _1151_;
	assign _1469_ = _1468_ | _1433_;
	assign _1470_ = _1469_ | _1432_;
	assign _1471_ = _1470_ | _1431_;
	assign _1472_ = _1089_ & ~_1471_;
	assign _1473_ = _1472_ | _1467_;
	assign _1474_ = _1449_ | _0731_;
	assign _1475_ = _1474_ | _1446_;
	assign _1476_ = _1475_ | _1445_;
	assign _1477_ = _1476_ | _1444_;
	assign _1478_ = _1389_ & ~_1477_;
	assign _1479_ = _1478_ | _1473_;
	assign _1480_ = _1411_ | _0417_;
	assign _1481_ = _1480_ | _1406_;
	assign _1482_ = _1481_ | _1405_;
	assign _1483_ = _0286_ & ~_1482_;
	assign _1484_ = _1424_ | _0808_;
	assign _1485_ = _1484_ | _1418_;
	assign _1486_ = _1485_ | _1417_;
	assign _1487_ = _0720_ & ~_1486_;
	assign _1488_ = _1487_ | _1483_;
	assign _1489_ = _1437_ | _1172_;
	assign _1490_ = _1489_ | _1432_;
	assign _1491_ = _1490_ | _1431_;
	assign _1492_ = _1089_ & ~_1491_;
	assign _1493_ = _1492_ | _1488_;
	assign _1494_ = _1450_ | _1396_;
	assign _1495_ = _1494_ | _1445_;
	assign _1496_ = _1495_ | _1444_;
	assign _1497_ = _1389_ & ~_1496_;
	assign _1498_ = _1497_ | _1493_;
	assign _1499_ = (\mchip.idx [3] ? _1498_ : _1479_);
	assign _1500_ = (\mchip.idx [4] ? _1499_ : _1456_);
	assign _1501_ = _1457_ | _0417_;
	assign _1502_ = _1501_ | _1406_;
	assign _1503_ = _1502_ | _1405_;
	assign _1504_ = _0286_ & ~_1503_;
	assign _1505_ = _1462_ | _0808_;
	assign _1506_ = _1505_ | _1418_;
	assign _1507_ = _1506_ | _1417_;
	assign _1508_ = _0720_ & ~_1507_;
	assign _1509_ = _1508_ | _1504_;
	assign _1510_ = _1468_ | _1172_;
	assign _1511_ = _1510_ | _1432_;
	assign _1512_ = _1511_ | _1431_;
	assign _1513_ = _1089_ & ~_1512_;
	assign _1514_ = _1513_ | _1509_;
	assign _1515_ = _1474_ | _1396_;
	assign _1516_ = _1515_ | _1445_;
	assign _1517_ = _1516_ | _1444_;
	assign _1518_ = _1389_ & ~_1517_;
	assign _1519_ = _1518_ | _1514_;
	assign _1520_ = _1412_ | _0450_;
	assign _1521_ = _1520_ | _1405_;
	assign _1522_ = _0286_ & ~_1521_;
	assign _1523_ = _1425_ | _0841_;
	assign _1524_ = _1523_ | _1417_;
	assign _1525_ = _0720_ & ~_1524_;
	assign _1526_ = _1525_ | _1522_;
	assign _1527_ = _1438_ | _1205_;
	assign _1528_ = _1527_ | _1431_;
	assign _1529_ = _1089_ & ~_1528_;
	assign _1530_ = _1529_ | _1526_;
	assign _1531_ = _1451_ | _1399_;
	assign _1532_ = _1531_ | _1444_;
	assign _1533_ = _1389_ & ~_1532_;
	assign _1534_ = _1533_ | _1530_;
	assign _1535_ = (\mchip.idx [3] ? _1534_ : _1519_);
	assign _1536_ = _1458_ | _0450_;
	assign _1537_ = _1536_ | _1405_;
	assign _1538_ = _0286_ & ~_1537_;
	assign _1539_ = _1463_ | _0841_;
	assign _1540_ = _1539_ | _1417_;
	assign _1541_ = _0720_ & ~_1540_;
	assign _1542_ = _1541_ | _1538_;
	assign _1543_ = _1469_ | _1205_;
	assign _1544_ = _1543_ | _1431_;
	assign _1545_ = _1089_ & ~_1544_;
	assign _1546_ = _1545_ | _1542_;
	assign _1547_ = _1475_ | _1399_;
	assign _1548_ = _1547_ | _1444_;
	assign _1549_ = _1389_ & ~_1548_;
	assign _1550_ = _1549_ | _1546_;
	assign _1551_ = _1480_ | _0450_;
	assign _1552_ = _1551_ | _1405_;
	assign _1553_ = _0286_ & ~_1552_;
	assign _1554_ = _1484_ | _0841_;
	assign _1555_ = _1554_ | _1417_;
	assign _1556_ = _0720_ & ~_1555_;
	assign _1557_ = _1556_ | _1553_;
	assign _1558_ = _1489_ | _1205_;
	assign _1559_ = _1558_ | _1431_;
	assign _1560_ = _1089_ & ~_1559_;
	assign _1561_ = _1560_ | _1557_;
	assign _1562_ = _1494_ | _1399_;
	assign _1563_ = _1562_ | _1444_;
	assign _1564_ = _1389_ & ~_1563_;
	assign _1565_ = _1564_ | _1561_;
	assign _1566_ = (\mchip.idx [3] ? _1565_ : _1550_);
	assign _1567_ = (\mchip.idx [4] ? _1566_ : _1535_);
	assign _1568_ = (\mchip.idx [5] ? _1567_ : _1500_);
	assign _1569_ = _1501_ | _0450_;
	assign _1570_ = _1569_ | _1405_;
	assign _1571_ = _0286_ & ~_1570_;
	assign _1572_ = _1505_ | _0841_;
	assign _1573_ = _1572_ | _1417_;
	assign _1574_ = _0720_ & ~_1573_;
	assign _1575_ = _1574_ | _1571_;
	assign _1576_ = _1510_ | _1205_;
	assign _1577_ = _1576_ | _1431_;
	assign _1578_ = _1089_ & ~_1577_;
	assign _1579_ = _1578_ | _1575_;
	assign _1580_ = _1515_ | _1399_;
	assign _1581_ = _1580_ | _1444_;
	assign _1582_ = _1389_ & ~_1581_;
	assign _1583_ = _1582_ | _1579_;
	assign _1584_ = _1413_ | _1404_;
	assign _1585_ = _0286_ & ~_1584_;
	assign _1586_ = _1426_ | _1416_;
	assign _1587_ = _0720_ & ~_1586_;
	assign _1588_ = _1587_ | _1585_;
	assign _1589_ = _1439_ | _1430_;
	assign _1590_ = _1089_ & ~_1589_;
	assign _1591_ = _1590_ | _1588_;
	assign _1592_ = _1452_ | _1443_;
	assign _1593_ = _1389_ & ~_1592_;
	assign _1594_ = _1593_ | _1591_;
	assign _1595_ = (\mchip.idx [3] ? _1594_ : _1583_);
	assign _1596_ = _1459_ | _1404_;
	assign _1597_ = _0286_ & ~_1596_;
	assign _1598_ = _1464_ | _1416_;
	assign _1599_ = _0720_ & ~_1598_;
	assign _1600_ = _1599_ | _1597_;
	assign _1601_ = _1470_ | _1430_;
	assign _1602_ = _1089_ & ~_1601_;
	assign _1603_ = _1602_ | _1600_;
	assign _1604_ = _1476_ | _1443_;
	assign _1605_ = _1389_ & ~_1604_;
	assign _1606_ = _1605_ | _1603_;
	assign _1607_ = _1481_ | _1404_;
	assign _1608_ = _0286_ & ~_1607_;
	assign _1609_ = _1485_ | _1416_;
	assign _1610_ = _0720_ & ~_1609_;
	assign _1611_ = _1610_ | _1608_;
	assign _1612_ = _1490_ | _1430_;
	assign _1613_ = _1089_ & ~_1612_;
	assign _1614_ = _1613_ | _1611_;
	assign _1615_ = _1495_ | _1443_;
	assign _1616_ = _1389_ & ~_1615_;
	assign _1617_ = _1616_ | _1614_;
	assign _1618_ = (\mchip.idx [3] ? _1617_ : _1606_);
	assign _1619_ = (\mchip.idx [4] ? _1618_ : _1595_);
	assign _1620_ = _1502_ | _1404_;
	assign _1621_ = _0286_ & ~_1620_;
	assign _1622_ = _1506_ | _1416_;
	assign _1623_ = _0720_ & ~_1622_;
	assign _1624_ = _1623_ | _1621_;
	assign _1625_ = _1511_ | _1430_;
	assign _1626_ = _1089_ & ~_1625_;
	assign _1627_ = _1626_ | _1624_;
	assign _1628_ = _1516_ | _1443_;
	assign _1629_ = _1389_ & ~_1628_;
	assign _1630_ = _1629_ | _1627_;
	assign _1631_ = _1520_ | _1404_;
	assign _1632_ = _0286_ & ~_1631_;
	assign _1633_ = _1523_ | _1416_;
	assign _1634_ = _0720_ & ~_1633_;
	assign _1635_ = _1634_ | _1632_;
	assign _1636_ = _1527_ | _1430_;
	assign _1637_ = _1089_ & ~_1636_;
	assign _1638_ = _1637_ | _1635_;
	assign _1640_ = _1531_ | _1443_;
	assign _1641_ = _1389_ & ~_1640_;
	assign _1642_ = _1641_ | _1638_;
	assign _1643_ = (\mchip.idx [3] ? _1642_ : _1630_);
	assign _1644_ = _1536_ | _1404_;
	assign _1645_ = _0286_ & ~_1644_;
	assign _1646_ = _1539_ | _1416_;
	assign _1647_ = _0720_ & ~_1646_;
	assign _1648_ = _1647_ | _1645_;
	assign _1649_ = _1543_ | _1430_;
	assign _1651_ = _1089_ & ~_1649_;
	assign _1652_ = _1651_ | _1648_;
	assign _1653_ = _1547_ | _1443_;
	assign _1654_ = _1389_ & ~_1653_;
	assign _1655_ = _1654_ | _1652_;
	assign _1656_ = _1551_ | _1404_;
	assign _1657_ = _0286_ & ~_1656_;
	assign _1658_ = _1554_ | _1416_;
	assign _1659_ = _0720_ & ~_1658_;
	assign _1660_ = _1659_ | _1657_;
	assign _1661_ = _1558_ | _1430_;
	assign _1662_ = _1089_ & ~_1661_;
	assign _1663_ = _1662_ | _1660_;
	assign _1664_ = _1562_ | _1443_;
	assign _1665_ = _1389_ & ~_1664_;
	assign _1666_ = _1665_ | _1663_;
	assign _1667_ = (\mchip.idx [3] ? _1666_ : _1655_);
	assign _1668_ = (\mchip.idx [4] ? _1667_ : _1643_);
	assign _1669_ = (\mchip.idx [5] ? _1668_ : _1619_);
	assign \mchip.iout [0] = (\mchip.idx [6] ? _1669_ : _1568_);
	assign _1671_ = ~_0033_;
	assign _1672_ = ~(_1681_ & _1717_);
	assign _1673_ = _1672_ | ~_0395_;
	assign _1674_ = _1673_ | ~_0417_;
	assign _1675_ = _1674_ | ~_0450_;
	assign _1676_ = _1675_ | ~_1404_;
	assign _1677_ = _0286_ & ~_1676_;
	assign _1678_ = \mchip.x [1] | ~\mchip.x [0];
	assign _1679_ = _1678_ | ~_1728_;
	assign _1680_ = _1679_ | ~_0731_;
	assign _1682_ = _1680_ | ~_0808_;
	assign _1683_ = _1682_ | ~_0841_;
	assign _1684_ = _1683_ | ~_1416_;
	assign _1685_ = _0720_ & ~_1684_;
	assign _1686_ = _1685_ | _1677_;
	assign _1687_ = _1679_ | ~_1151_;
	assign _1688_ = _1687_ | ~_1172_;
	assign _1689_ = _1688_ | ~_1205_;
	assign _1690_ = _1689_ | ~_1430_;
	assign _1691_ = _1089_ & ~_1690_;
	assign _1692_ = _1691_ | _1686_;
	assign _1693_ = _1680_ | ~_1396_;
	assign _1694_ = _1693_ | ~_1399_;
	assign _1695_ = _1694_ | ~_1443_;
	assign _1696_ = _1389_ & ~_1695_;
	assign _1698_ = _1696_ | _1692_;
	assign _1699_ = _1672_ | _0395_;
	assign _1700_ = _1699_ | ~_0417_;
	assign _1701_ = _1700_ | ~_0450_;
	assign _1702_ = _1701_ | ~_1404_;
	assign _1703_ = _0286_ & ~_1702_;
	assign _1704_ = _1679_ | _0731_;
	assign _1705_ = _1704_ | ~_0808_;
	assign _1706_ = _1705_ | ~_0841_;
	assign _1707_ = _1706_ | ~_1416_;
	assign _1708_ = _0720_ & ~_1707_;
	assign _1709_ = _1708_ | _1703_;
	assign _1710_ = _1679_ | _1151_;
	assign _1711_ = _1710_ | ~_1172_;
	assign _1712_ = _1711_ | ~_1205_;
	assign _1713_ = _1712_ | ~_1430_;
	assign _1714_ = _1089_ & ~_1713_;
	assign _1715_ = _1714_ | _1709_;
	assign _1716_ = _1704_ | ~_1396_;
	assign _1718_ = _1716_ | ~_1399_;
	assign _1719_ = _1718_ | ~_1443_;
	assign _1720_ = _1389_ & ~_1719_;
	assign _1721_ = _1720_ | _1715_;
	assign _1722_ = (\mchip.idx [3] ? _1721_ : _1698_);
	assign _1723_ = _1673_ | _0417_;
	assign _1724_ = _1723_ | ~_0450_;
	assign _1725_ = _1724_ | ~_1404_;
	assign _1726_ = _0286_ & ~_1725_;
	assign _1727_ = _1680_ | _0808_;
	assign _1729_ = _1727_ | ~_0841_;
	assign _1730_ = _1729_ | ~_1416_;
	assign _1731_ = _0720_ & ~_1730_;
	assign _1732_ = _1731_ | _1726_;
	assign _1733_ = _1687_ | _1172_;
	assign _1734_ = _1733_ | ~_1205_;
	assign _1735_ = _1734_ | ~_1430_;
	assign _1736_ = _1089_ & ~_1735_;
	assign _1737_ = _1736_ | _1732_;
	assign _1738_ = _1680_ | _1396_;
	assign _1740_ = _1738_ | ~_1399_;
	assign _1741_ = _1740_ | ~_1443_;
	assign _1742_ = _1389_ & ~_1741_;
	assign _1743_ = _1742_ | _1737_;
	assign _1744_ = _1699_ | _0417_;
	assign _1745_ = _1744_ | ~_0450_;
	assign _1746_ = _1745_ | ~_1404_;
	assign _1747_ = _0286_ & ~_1746_;
	assign _1748_ = _1704_ | _0808_;
	assign _1749_ = _1748_ | ~_0841_;
	assign _1751_ = _1749_ | ~_1416_;
	assign _1752_ = _0720_ & ~_1751_;
	assign _1753_ = _1752_ | _1747_;
	assign _1754_ = _1710_ | _1172_;
	assign _1755_ = _1754_ | ~_1205_;
	assign _1756_ = _1755_ | ~_1430_;
	assign _1757_ = _1089_ & ~_1756_;
	assign _1758_ = _1757_ | _1753_;
	assign _1759_ = _1704_ | _1396_;
	assign _1760_ = _1759_ | ~_1399_;
	assign _1761_ = _1760_ | ~_1443_;
	assign _1762_ = _1389_ & ~_1761_;
	assign _1763_ = _1762_ | _1758_;
	assign _1764_ = (\mchip.idx [3] ? _1763_ : _1743_);
	assign _1765_ = (\mchip.idx [4] ? _1764_ : _1722_);
	assign _1766_ = _1674_ | _0450_;
	assign _1767_ = _1766_ | ~_1404_;
	assign _1768_ = _0286_ & ~_1767_;
	assign _1769_ = _1682_ | _0841_;
	assign _1770_ = _1769_ | ~_1416_;
	assign _1772_ = _0720_ & ~_1770_;
	assign _1773_ = _1772_ | _1768_;
	assign _1774_ = _1688_ | _1205_;
	assign _1775_ = _1774_ | ~_1430_;
	assign _1776_ = _1089_ & ~_1775_;
	assign _1777_ = _1776_ | _1773_;
	assign _1778_ = _1693_ | _1399_;
	assign _1779_ = _1778_ | ~_1443_;
	assign _1780_ = _1389_ & ~_1779_;
	assign _1781_ = _1780_ | _1777_;
	assign _1783_ = _1700_ | _0450_;
	assign _1784_ = _1783_ | ~_1404_;
	assign _1785_ = _0286_ & ~_1784_;
	assign _1786_ = _1705_ | _0841_;
	assign _1787_ = _1786_ | ~_1416_;
	assign _1788_ = _0720_ & ~_1787_;
	assign _1789_ = _1788_ | _1785_;
	assign _1790_ = _1711_ | _1205_;
	assign _1791_ = _1790_ | ~_1430_;
	assign _1792_ = _1089_ & ~_1791_;
	assign _1793_ = _1792_ | _1789_;
	assign _1794_ = _1716_ | _1399_;
	assign _1795_ = _1794_ | ~_1443_;
	assign _1796_ = _1389_ & ~_1795_;
	assign _1797_ = _1796_ | _1793_;
	assign _1798_ = (\mchip.idx [3] ? _1797_ : _1781_);
	assign _1799_ = _1723_ | _0450_;
	assign _1800_ = _1799_ | ~_1404_;
	assign _1801_ = _0286_ & ~_1800_;
	assign _1802_ = _1727_ | _0841_;
	assign _1804_ = _1802_ | ~_1416_;
	assign _1805_ = _0720_ & ~_1804_;
	assign _1806_ = _1805_ | _1801_;
	assign _1807_ = _1733_ | _1205_;
	assign _1808_ = _1807_ | ~_1430_;
	assign _1809_ = _1089_ & ~_1808_;
	assign _1810_ = _1809_ | _1806_;
	assign _1811_ = _1738_ | _1399_;
	assign _1812_ = _1811_ | ~_1443_;
	assign _1813_ = _1389_ & ~_1812_;
	assign _1815_ = _1813_ | _1810_;
	assign _1816_ = _1744_ | _0450_;
	assign _1817_ = _1816_ | ~_1404_;
	assign _1818_ = _0286_ & ~_1817_;
	assign _1819_ = _1748_ | _0841_;
	assign _1820_ = _1819_ | ~_1416_;
	assign _1821_ = _0720_ & ~_1820_;
	assign _1822_ = _1821_ | _1818_;
	assign _1823_ = _1754_ | _1205_;
	assign _1824_ = _1823_ | ~_1430_;
	assign _1825_ = _1089_ & ~_1824_;
	assign _1826_ = _1825_ | _1822_;
	assign _1827_ = _1759_ | _1399_;
	assign _1828_ = _1827_ | ~_1443_;
	assign _1829_ = _1389_ & ~_1828_;
	assign _1830_ = _1829_ | _1826_;
	assign _1831_ = (\mchip.idx [3] ? _1830_ : _1815_);
	assign _1832_ = (\mchip.idx [4] ? _1831_ : _1798_);
	assign _1833_ = (\mchip.idx [5] ? _1832_ : _1765_);
	assign _1834_ = _1675_ | _1404_;
	assign _1836_ = _0286_ & ~_1834_;
	assign _1837_ = _1683_ | _1416_;
	assign _1838_ = _0720_ & ~_1837_;
	assign _1839_ = _1838_ | _1836_;
	assign _1840_ = _1689_ | _1430_;
	assign _1841_ = _1089_ & ~_1840_;
	assign _1842_ = _1841_ | _1839_;
	assign _1843_ = _1694_ | _1443_;
	assign _1844_ = _1389_ & ~_1843_;
	assign _1845_ = _1844_ | _1842_;
	assign _1847_ = _1701_ | _1404_;
	assign _1848_ = _0286_ & ~_1847_;
	assign _1849_ = _1706_ | _1416_;
	assign _1850_ = _0720_ & ~_1849_;
	assign _1851_ = _1850_ | _1848_;
	assign _1852_ = _1712_ | _1430_;
	assign _1853_ = _1089_ & ~_1852_;
	assign _1854_ = _1853_ | _1851_;
	assign _1855_ = _1718_ | _1443_;
	assign _1856_ = _1389_ & ~_1855_;
	assign _1858_ = _1856_ | _1854_;
	assign _1859_ = (\mchip.idx [3] ? _1858_ : _1845_);
	assign _1860_ = _1724_ | _1404_;
	assign _1861_ = _0286_ & ~_1860_;
	assign _1862_ = _1729_ | _1416_;
	assign _1863_ = _0720_ & ~_1862_;
	assign _1864_ = _1863_ | _1861_;
	assign _1865_ = _1734_ | _1430_;
	assign _1866_ = _1089_ & ~_1865_;
	assign _1867_ = _1866_ | _1864_;
	assign _1869_ = _1740_ | _1443_;
	assign _1870_ = _1389_ & ~_1869_;
	assign _1871_ = _1870_ | _1867_;
	assign _1872_ = _1745_ | _1404_;
	assign _1873_ = _0286_ & ~_1872_;
	assign _1874_ = _1749_ | _1416_;
	assign _1875_ = _0720_ & ~_1874_;
	assign _1876_ = _1875_ | _1873_;
	assign _1877_ = _1755_ | _1430_;
	assign _1878_ = _1089_ & ~_1877_;
	assign _1880_ = _1878_ | _1876_;
	assign _1881_ = _1760_ | _1443_;
	assign _1882_ = _1389_ & ~_1881_;
	assign _1883_ = _1882_ | _1880_;
	assign _1884_ = (\mchip.idx [3] ? _1883_ : _1871_);
	assign _1885_ = (\mchip.idx [4] ? _1884_ : _1859_);
	assign _1886_ = _1766_ | _1404_;
	assign _1887_ = _0286_ & ~_1886_;
	assign _1888_ = _1769_ | _1416_;
	assign _1889_ = _0720_ & ~_1888_;
	assign _1891_ = _1889_ | _1887_;
	assign _1892_ = _1774_ | _1430_;
	assign _1893_ = _1089_ & ~_1892_;
	assign _1894_ = _1893_ | _1891_;
	assign _1895_ = _1778_ | _1443_;
	assign _1896_ = _1389_ & ~_1895_;
	assign _1897_ = _1896_ | _1894_;
	assign _1898_ = _1783_ | _1404_;
	assign _1899_ = _0286_ & ~_1898_;
	assign _1900_ = _1786_ | _1416_;
	assign _1901_ = _0720_ & ~_1900_;
	assign _1902_ = _1901_ | _1899_;
	assign _1903_ = _1790_ | _1430_;
	assign _1904_ = _1089_ & ~_1903_;
	assign _1905_ = _1904_ | _1902_;
	assign _1906_ = _1794_ | _1443_;
	assign _1907_ = _1389_ & ~_1906_;
	assign _1908_ = _1907_ | _1905_;
	assign _1909_ = (\mchip.idx [3] ? _1908_ : _1897_);
	assign _1910_ = _1799_ | _1404_;
	assign _1912_ = _0286_ & ~_1910_;
	assign _1913_ = _1802_ | _1416_;
	assign _1914_ = _0720_ & ~_1913_;
	assign _1915_ = _1914_ | _1912_;
	assign _1916_ = _1807_ | _1430_;
	assign _1917_ = _1089_ & ~_1916_;
	assign _1918_ = _1917_ | _1915_;
	assign _1919_ = _1811_ | _1443_;
	assign _1920_ = _1389_ & ~_1919_;
	assign _1921_ = _1920_ | _1918_;
	assign _1923_ = _1816_ | _1404_;
	assign _1924_ = _0286_ & ~_1923_;
	assign _1925_ = _1819_ | _1416_;
	assign _1926_ = _0720_ & ~_1925_;
	assign _1927_ = _1926_ | _1924_;
	assign _1928_ = _1823_ | _1430_;
	assign _1929_ = _1089_ & ~_1928_;
	assign _1930_ = _1929_ | _1927_;
	assign _1931_ = _1827_ | _1443_;
	assign _1932_ = _1389_ & ~_1931_;
	assign _1934_ = _1932_ | _1930_;
	assign _1935_ = (\mchip.idx [3] ? _1934_ : _1921_);
	assign _1936_ = (\mchip.idx [4] ? _1935_ : _1909_);
	assign _1937_ = (\mchip.idx [5] ? _1936_ : _1885_);
	assign \mchip.iout [1] = (\mchip.idx [6] ? _1937_ : _1833_);
	assign _1938_ = _1678_ | ~_0362_;
	assign _1939_ = _1938_ | ~_0395_;
	assign _1940_ = _1939_ | ~_0417_;
	assign _1941_ = _1940_ | ~_0450_;
	assign _1942_ = _1941_ | ~_1404_;
	assign _1944_ = _0286_ & ~_1942_;
	assign _1945_ = \mchip.x [0] | ~\mchip.x [1];
	assign _1946_ = _1945_ | ~_1728_;
	assign _1947_ = _1946_ | ~_0731_;
	assign _1948_ = _1947_ | ~_0808_;
	assign _1949_ = _1948_ | ~_0841_;
	assign _1950_ = _1949_ | ~_1416_;
	assign _1951_ = _0720_ & ~_1950_;
	assign _1952_ = _1951_ | _1944_;
	assign _1954_ = _1946_ | ~_1151_;
	assign _1955_ = _1954_ | ~_1172_;
	assign _1956_ = _1955_ | ~_1205_;
	assign _1957_ = _1956_ | ~_1430_;
	assign _1958_ = _1089_ & ~_1957_;
	assign _1959_ = _1958_ | _1952_;
	assign _1960_ = _1947_ | ~_1396_;
	assign _1961_ = _1960_ | ~_1399_;
	assign _1962_ = _1961_ | ~_1443_;
	assign _1963_ = _1389_ & ~_1962_;
	assign _1964_ = _1963_ | _1959_;
	assign _1965_ = _1938_ | _0395_;
	assign _1966_ = _1965_ | ~_0417_;
	assign _1967_ = _1966_ | ~_0450_;
	assign _1968_ = _1967_ | ~_1404_;
	assign _1969_ = _0286_ & ~_1968_;
	assign _1971_ = _1946_ | _0731_;
	assign _1972_ = _1971_ | ~_0808_;
	assign _1973_ = _1972_ | ~_0841_;
	assign _1974_ = _1973_ | ~_1416_;
	assign _1975_ = _0720_ & ~_1974_;
	assign _1976_ = _1975_ | _1969_;
	assign _1977_ = _1946_ | _1151_;
	assign _1978_ = _1977_ | ~_1172_;
	assign _1979_ = _1978_ | ~_1205_;
	assign _1980_ = _1979_ | ~_1430_;
	assign _1982_ = _1089_ & ~_1980_;
	assign _1983_ = _1982_ | _1976_;
	assign _1984_ = _1971_ | ~_1396_;
	assign _1985_ = _1984_ | ~_1399_;
	assign _1986_ = _1985_ | ~_1443_;
	assign _1987_ = _1389_ & ~_1986_;
	assign _1988_ = _1987_ | _1983_;
	assign _1989_ = (\mchip.idx [3] ? _1988_ : _1964_);
	assign _1990_ = _1939_ | _0417_;
	assign _1992_ = _1990_ | ~_0450_;
	assign _1993_ = _1992_ | ~_1404_;
	assign _1994_ = _0286_ & ~_1993_;
	assign _1995_ = _1947_ | _0808_;
	assign _1996_ = _1995_ | ~_0841_;
	assign _1997_ = _1996_ | ~_1416_;
	assign _1998_ = _0720_ & ~_1997_;
	assign _1999_ = _1998_ | _1994_;
	assign _2000_ = _1954_ | _1172_;
	assign _2001_ = _2000_ | ~_1205_;
	assign _2003_ = _2001_ | ~_1430_;
	assign _2004_ = _1089_ & ~_2003_;
	assign _2005_ = _2004_ | _1999_;
	assign _2006_ = _1947_ | _1396_;
	assign _2007_ = _2006_ | ~_1399_;
	assign _2008_ = _2007_ | ~_1443_;
	assign _2009_ = _1389_ & ~_2008_;
	assign _2010_ = _2009_ | _2005_;
	assign _2011_ = _1965_ | _0417_;
	assign _2012_ = _2011_ | ~_0450_;
	assign _2014_ = _2012_ | ~_1404_;
	assign _2015_ = _0286_ & ~_2014_;
	assign _2016_ = _1971_ | _0808_;
	assign _2017_ = _2016_ | ~_0841_;
	assign _2018_ = _2017_ | ~_1416_;
	assign _2019_ = _0720_ & ~_2018_;
	assign _2020_ = _2019_ | _2015_;
	assign _2021_ = _1977_ | _1172_;
	assign _2022_ = _2021_ | ~_1205_;
	assign _2023_ = _2022_ | ~_1430_;
	assign _2025_ = _1089_ & ~_2023_;
	assign _2026_ = _2025_ | _2020_;
	assign _2027_ = _1971_ | _1396_;
	assign _2028_ = _2027_ | ~_1399_;
	assign _2029_ = _2028_ | ~_1443_;
	assign _2030_ = _1389_ & ~_2029_;
	assign _2031_ = _2030_ | _2026_;
	assign _2032_ = (\mchip.idx [3] ? _2031_ : _2010_);
	assign _2033_ = (\mchip.idx [4] ? _2032_ : _1989_);
	assign _2034_ = _1940_ | _0450_;
	assign _2036_ = _2034_ | ~_1404_;
	assign _2037_ = _0286_ & ~_2036_;
	assign _2038_ = _1948_ | _0841_;
	assign _2039_ = _2038_ | ~_1416_;
	assign _2040_ = _0720_ & ~_2039_;
	assign _2041_ = _2040_ | _2037_;
	assign _2042_ = _1955_ | _1205_;
	assign _2043_ = _2042_ | ~_1430_;
	assign _2044_ = _1089_ & ~_2043_;
	assign _2045_ = _2044_ | _2041_;
	assign _2047_ = _1960_ | _1399_;
	assign _2048_ = _2047_ | ~_1443_;
	assign _2049_ = _1389_ & ~_2048_;
	assign _2050_ = _2049_ | _2045_;
	assign _2051_ = _1966_ | _0450_;
	assign _2052_ = _2051_ | ~_1404_;
	assign _2053_ = _0286_ & ~_2052_;
	assign _2054_ = _1972_ | _0841_;
	assign _2055_ = _2054_ | ~_1416_;
	assign _2056_ = _0720_ & ~_2055_;
	assign _2057_ = _2056_ | _2053_;
	assign _2058_ = _1978_ | _1205_;
	assign _2059_ = _2058_ | ~_1430_;
	assign _2060_ = _1089_ & ~_2059_;
	assign _2061_ = _2060_ | _2057_;
	assign _2062_ = _1984_ | _1399_;
	assign _2063_ = _2062_ | ~_1443_;
	assign _2064_ = _1389_ & ~_2063_;
	assign _2065_ = _2064_ | _2061_;
	assign _2066_ = (\mchip.idx [3] ? _2065_ : _2050_);
	assign _2067_ = _1990_ | _0450_;
	assign _2068_ = _2067_ | ~_1404_;
	assign _2069_ = _0286_ & ~_2068_;
	assign _2070_ = _1995_ | _0841_;
	assign _2071_ = _2070_ | ~_1416_;
	assign _2072_ = _0720_ & ~_2071_;
	assign _2073_ = _2072_ | _2069_;
	assign _2074_ = _2000_ | _1205_;
	assign _2075_ = _2074_ | ~_1430_;
	assign _2076_ = _1089_ & ~_2075_;
	assign _2077_ = _2076_ | _2073_;
	assign _2078_ = _2006_ | _1399_;
	assign _2079_ = _2078_ | ~_1443_;
	assign _2080_ = _1389_ & ~_2079_;
	assign _2081_ = _2080_ | _2077_;
	assign _2082_ = _2011_ | _0450_;
	assign _2083_ = _2082_ | ~_1404_;
	assign _2084_ = _0286_ & ~_2083_;
	assign _2085_ = _2016_ | _0841_;
	assign _2086_ = _2085_ | ~_1416_;
	assign _2087_ = _0720_ & ~_2086_;
	assign _2088_ = _2087_ | _2084_;
	assign _2089_ = _2021_ | _1205_;
	assign _2090_ = _2089_ | ~_1430_;
	assign _2091_ = _1089_ & ~_2090_;
	assign _2092_ = _2091_ | _2088_;
	assign _2093_ = _2027_ | _1399_;
	assign _2094_ = _2093_ | ~_1443_;
	assign _2095_ = _1389_ & ~_2094_;
	assign _2096_ = _2095_ | _2092_;
	assign _2098_ = (\mchip.idx [3] ? _2096_ : _2081_);
	assign _2099_ = (\mchip.idx [4] ? _2098_ : _2066_);
	assign _2100_ = (\mchip.idx [5] ? _2099_ : _2033_);
	assign _2101_ = _1941_ | _1404_;
	assign _2102_ = _0286_ & ~_2101_;
	assign _2103_ = _1949_ | _1416_;
	assign _2104_ = _0720_ & ~_2103_;
	assign _2105_ = _2104_ | _2102_;
	assign _2106_ = _1956_ | _1430_;
	assign _2107_ = _1089_ & ~_2106_;
	assign _2108_ = _2107_ | _2105_;
	assign _2109_ = _1961_ | _1443_;
	assign _2110_ = _1389_ & ~_2109_;
	assign _2111_ = _2110_ | _2108_;
	assign _2112_ = _1967_ | _1404_;
	assign _2113_ = _0286_ & ~_2112_;
	assign _2114_ = _1973_ | _1416_;
	assign _2115_ = _0720_ & ~_2114_;
	assign _2116_ = _2115_ | _2113_;
	assign _2117_ = _1979_ | _1430_;
	assign _2119_ = _1089_ & ~_2117_;
	assign _2120_ = _2119_ | _2116_;
	assign _2121_ = _1985_ | _1443_;
	assign _2122_ = _1389_ & ~_2121_;
	assign _2123_ = _2122_ | _2120_;
	assign _2124_ = (\mchip.idx [3] ? _2123_ : _2111_);
	assign _2125_ = _1992_ | _1404_;
	assign _2126_ = _0286_ & ~_2125_;
	assign _2127_ = _1996_ | _1416_;
	assign _2128_ = _0720_ & ~_2127_;
	assign _2130_ = _2128_ | _2126_;
	assign _2131_ = _2001_ | _1430_;
	assign _2132_ = _1089_ & ~_2131_;
	assign _2133_ = _2132_ | _2130_;
	assign _2134_ = _2007_ | _1443_;
	assign _2135_ = _1389_ & ~_2134_;
	assign _2136_ = _2135_ | _2133_;
	assign _2137_ = _2012_ | _1404_;
	assign _2138_ = _0286_ & ~_2137_;
	assign _2139_ = _2017_ | _1416_;
	assign _2140_ = _0720_ & ~_2139_;
	assign _2141_ = _2140_ | _2138_;
	assign _2142_ = _2022_ | _1430_;
	assign _2143_ = _1089_ & ~_2142_;
	assign _2144_ = _2143_ | _2141_;
	assign _2145_ = _2028_ | _1443_;
	assign _2146_ = _1389_ & ~_2145_;
	assign _2147_ = _2146_ | _2144_;
	assign _2148_ = (\mchip.idx [3] ? _2147_ : _2136_);
	assign _2149_ = (\mchip.idx [4] ? _2148_ : _2124_);
	assign _2150_ = _2034_ | _1404_;
	assign _2151_ = _0286_ & ~_2150_;
	assign _2152_ = _2038_ | _1416_;
	assign _2153_ = _0720_ & ~_2152_;
	assign _2154_ = _2153_ | _2151_;
	assign _2155_ = _2042_ | _1430_;
	assign _2156_ = _1089_ & ~_2155_;
	assign _2157_ = _2156_ | _2154_;
	assign _2158_ = _2047_ | _1443_;
	assign _2159_ = _1389_ & ~_2158_;
	assign _2161_ = _2159_ | _2157_;
	assign _2162_ = _2051_ | _1404_;
	assign _2163_ = _0286_ & ~_2162_;
	assign _2164_ = _2054_ | _1416_;
	assign _2165_ = _0720_ & ~_2164_;
	assign _2166_ = _2165_ | _2163_;
	assign _2167_ = _2058_ | _1430_;
	assign _2168_ = _1089_ & ~_2167_;
	assign _2169_ = _2168_ | _2166_;
	assign _2170_ = _2062_ | _1443_;
	assign _2171_ = _1389_ & ~_2170_;
	assign _2172_ = _2171_ | _2169_;
	assign _2173_ = (\mchip.idx [3] ? _2172_ : _2161_);
	assign _2174_ = _2067_ | _1404_;
	assign _2175_ = _0286_ & ~_2174_;
	assign _2176_ = _2070_ | _1416_;
	assign _2177_ = _0720_ & ~_2176_;
	assign _2178_ = _2177_ | _2175_;
	assign _2179_ = _2074_ | _1430_;
	assign _2180_ = _1089_ & ~_2179_;
	assign _0009_ = _2180_ | _2178_;
	assign _0010_ = _2078_ | _1443_;
	assign _0011_ = _1389_ & ~_0010_;
	assign _0012_ = _0011_ | _0009_;
	assign _0013_ = _2082_ | _1404_;
	assign _0014_ = _0286_ & ~_0013_;
	assign _0015_ = _2085_ | _1416_;
	assign _0016_ = _0720_ & ~_0015_;
	assign _0017_ = _0016_ | _0014_;
	assign _0018_ = _2089_ | _1430_;
	assign _0019_ = _1089_ & ~_0018_;
	assign _0020_ = _0019_ | _0017_;
	assign _0021_ = _2093_ | _1443_;
	assign _0022_ = _1389_ & ~_0021_;
	assign _0023_ = _0022_ | _0020_;
	assign _0024_ = (\mchip.idx [3] ? _0023_ : _0012_);
	assign _0025_ = (\mchip.idx [4] ? _0024_ : _2173_);
	assign _0026_ = (\mchip.idx [5] ? _0025_ : _2149_);
	assign \mchip.iout [2] = (\mchip.idx [6] ? _0026_ : _2100_);
	assign _0027_ = _1945_ | ~_0362_;
	assign _0028_ = _0027_ | ~_0395_;
	assign _0029_ = _0028_ | ~_0417_;
	assign _0030_ = _0029_ | ~_0450_;
	assign _0031_ = _0030_ | ~_1404_;
	assign _0032_ = _0286_ & ~_0031_;
	assign _0034_ = _0033_ | ~_1728_;
	assign _0035_ = _0034_ | ~_0731_;
	assign _0036_ = _0035_ | ~_0808_;
	assign _0037_ = _0036_ | ~_0841_;
	assign _0038_ = _0037_ | ~_1416_;
	assign _0039_ = _0720_ & ~_0038_;
	assign _0040_ = _0039_ | _0032_;
	assign _0041_ = ~(_1728_ & _1671_);
	assign _0042_ = _0041_ | ~_1151_;
	assign _0043_ = _0042_ | ~_1172_;
	assign _0044_ = _0043_ | ~_1205_;
	assign _0045_ = _0044_ | ~_1430_;
	assign _0046_ = _1089_ & ~_0045_;
	assign _0047_ = _0046_ | _0040_;
	assign _0049_ = _0035_ | ~_1396_;
	assign _0050_ = _0049_ | ~_1399_;
	assign _0051_ = _0050_ | ~_1443_;
	assign _0052_ = _1389_ & ~_0051_;
	assign _0053_ = _0052_ | _0047_;
	assign _0054_ = _0027_ | _0395_;
	assign _0055_ = _0054_ | ~_0417_;
	assign _0057_ = _0055_ | ~_0450_;
	assign _0058_ = _0057_ | ~_1404_;
	assign _0059_ = _0286_ & ~_0058_;
	assign _0060_ = _0034_ | _0731_;
	assign _0061_ = _0060_ | ~_0808_;
	assign _0062_ = _0061_ | ~_0841_;
	assign _0063_ = _0062_ | ~_1416_;
	assign _0064_ = _0720_ & ~_0063_;
	assign _0065_ = _0064_ | _0059_;
	assign _0066_ = _0041_ | _1151_;
	assign _0068_ = _0066_ | ~_1172_;
	assign _0069_ = _0068_ | ~_1205_;
	assign _0070_ = _0069_ | ~_1430_;
	assign _0071_ = _1089_ & ~_0070_;
	assign _0072_ = _0071_ | _0065_;
	assign _0073_ = _0060_ | ~_1396_;
	assign _0074_ = _0073_ | ~_1399_;
	assign _0075_ = _0074_ | ~_1443_;
	assign _0076_ = _1389_ & ~_0075_;
	assign _0078_ = _0076_ | _0072_;
	assign _0079_ = (\mchip.idx [3] ? _0078_ : _0053_);
	assign _0080_ = _0028_ | _0417_;
	assign _0081_ = _0080_ | ~_0450_;
	assign _0082_ = _0081_ | ~_1404_;
	assign _0083_ = _0286_ & ~_0082_;
	assign _0084_ = _0035_ | _0808_;
	assign _0085_ = _0084_ | ~_0841_;
	assign _0086_ = _0085_ | ~_1416_;
	assign _0087_ = _0720_ & ~_0086_;
	assign _0089_ = _0087_ | _0083_;
	assign _0090_ = _0042_ | _1172_;
	assign _0091_ = _0090_ | ~_1205_;
	assign _0092_ = _0091_ | ~_1430_;
	assign _0093_ = _1089_ & ~_0092_;
	assign _0094_ = _0093_ | _0089_;
	assign _0095_ = _0035_ | _1396_;
	assign _0096_ = _0095_ | ~_1399_;
	assign _0097_ = _0096_ | ~_1443_;
	assign _0098_ = _1389_ & ~_0097_;
	assign _0100_ = _0098_ | _0094_;
	assign _0101_ = _0054_ | _0417_;
	assign _0102_ = _0101_ | ~_0450_;
	assign _0103_ = _0102_ | ~_1404_;
	assign _0104_ = _0286_ & ~_0103_;
	assign _0105_ = _0060_ | _0808_;
	assign _0106_ = _0105_ | ~_0841_;
	assign _0107_ = _0106_ | ~_1416_;
	assign _0108_ = _0720_ & ~_0107_;
	assign _0109_ = _0108_ | _0104_;
	assign _0111_ = _0066_ | _1172_;
	assign _0112_ = _0111_ | ~_1205_;
	assign _0113_ = _0112_ | ~_1430_;
	assign _0114_ = _1089_ & ~_0113_;
	assign _0115_ = _0114_ | _0109_;
	assign _0116_ = _0060_ | _1396_;
	assign _0117_ = _0116_ | ~_1399_;
	assign _0118_ = _0117_ | ~_1443_;
	assign _0119_ = _1389_ & ~_0118_;
	assign _0120_ = _0119_ | _0115_;
	assign _0122_ = (\mchip.idx [3] ? _0120_ : _0100_);
	assign _0123_ = (\mchip.idx [4] ? _0122_ : _0079_);
	assign _0124_ = _0029_ | _0450_;
	assign _0125_ = _0124_ | ~_1404_;
	assign _0126_ = _0286_ & ~_0125_;
	assign _0127_ = _0036_ | _0841_;
	assign _0128_ = _0127_ | ~_1416_;
	assign _0129_ = _0720_ & ~_0128_;
	assign _0130_ = _0129_ | _0126_;
	assign _0131_ = _0043_ | _1205_;
	assign _0133_ = _0131_ | ~_1430_;
	assign _0134_ = _1089_ & ~_0133_;
	assign _0135_ = _0134_ | _0130_;
	assign _0136_ = _0049_ | _1399_;
	assign _0137_ = _0136_ | ~_1443_;
	assign _0138_ = _1389_ & ~_0137_;
	assign _0139_ = _0138_ | _0135_;
	assign _0140_ = _0055_ | _0450_;
	assign _0141_ = _0140_ | ~_1404_;
	assign _0142_ = _0286_ & ~_0141_;
	assign _0144_ = _0061_ | _0841_;
	assign _0145_ = _0144_ | ~_1416_;
	assign _0146_ = _0720_ & ~_0145_;
	assign _0147_ = _0146_ | _0142_;
	assign _0148_ = _0068_ | _1205_;
	assign _0149_ = _0148_ | ~_1430_;
	assign _0150_ = _1089_ & ~_0149_;
	assign _0151_ = _0150_ | _0147_;
	assign _0152_ = _0073_ | _1399_;
	assign _0153_ = _0152_ | ~_1443_;
	assign _0155_ = _1389_ & ~_0153_;
	assign _0156_ = _0155_ | _0151_;
	assign _0157_ = (\mchip.idx [3] ? _0156_ : _0139_);
	assign _0158_ = _0080_ | _0450_;
	assign _0159_ = _0158_ | ~_1404_;
	assign _0160_ = _0286_ & ~_0159_;
	assign _0161_ = _0084_ | _0841_;
	assign _0162_ = _0161_ | ~_1416_;
	assign _0163_ = _0720_ & ~_0162_;
	assign _0164_ = _0163_ | _0160_;
	assign _0166_ = _0090_ | _1205_;
	assign _0167_ = _0166_ | ~_1430_;
	assign _0168_ = _1089_ & ~_0167_;
	assign _0169_ = _0168_ | _0164_;
	assign _0170_ = _0095_ | _1399_;
	assign _0171_ = _0170_ | ~_1443_;
	assign _0172_ = _1389_ & ~_0171_;
	assign _0173_ = _0172_ | _0169_;
	assign _0174_ = _0101_ | _0450_;
	assign _0175_ = _0174_ | ~_1404_;
	assign _0177_ = _0286_ & ~_0175_;
	assign _0178_ = _0105_ | _0841_;
	assign _0179_ = _0178_ | ~_1416_;
	assign _0180_ = _0720_ & ~_0179_;
	assign _0181_ = _0180_ | _0177_;
	assign _0182_ = _0111_ | _1205_;
	assign _0183_ = _0182_ | ~_1430_;
	assign _0184_ = _1089_ & ~_0183_;
	assign _0185_ = _0184_ | _0181_;
	assign _0186_ = _0116_ | _1399_;
	assign _0188_ = _0186_ | ~_1443_;
	assign _0189_ = _1389_ & ~_0188_;
	assign _0190_ = _0189_ | _0185_;
	assign _0191_ = (\mchip.idx [3] ? _0190_ : _0173_);
	assign _0192_ = (\mchip.idx [4] ? _0191_ : _0157_);
	assign _0193_ = (\mchip.idx [5] ? _0192_ : _0123_);
	assign _0194_ = _0030_ | _1404_;
	assign _0195_ = _0286_ & ~_0194_;
	assign _0196_ = _0037_ | _1416_;
	assign _0197_ = _0720_ & ~_0196_;
	assign _0199_ = _0197_ | _0195_;
	assign _0200_ = _0044_ | _1430_;
	assign _0201_ = _1089_ & ~_0200_;
	assign _0202_ = _0201_ | _0199_;
	assign _0203_ = _0050_ | _1443_;
	assign _0204_ = _1389_ & ~_0203_;
	assign _0205_ = _0204_ | _0202_;
	assign _0206_ = _0057_ | _1404_;
	assign _0207_ = _0286_ & ~_0206_;
	assign _0208_ = _0062_ | _1416_;
	assign _0210_ = _0720_ & ~_0208_;
	assign _0211_ = _0210_ | _0207_;
	assign _0212_ = _0069_ | _1430_;
	assign _0213_ = _1089_ & ~_0212_;
	assign _0214_ = _0213_ | _0211_;
	assign _0215_ = _0074_ | _1443_;
	assign _0216_ = _1389_ & ~_0215_;
	assign _0217_ = _0216_ | _0214_;
	assign _0218_ = (\mchip.idx [3] ? _0217_ : _0205_);
	assign _0219_ = _0081_ | _1404_;
	assign _0221_ = _0286_ & ~_0219_;
	assign _0222_ = _0085_ | _1416_;
	assign _0223_ = _0720_ & ~_0222_;
	assign _0224_ = _0223_ | _0221_;
	assign _0225_ = _0091_ | _1430_;
	assign _0226_ = _1089_ & ~_0225_;
	assign _0227_ = _0226_ | _0224_;
	assign _0228_ = _0096_ | _1443_;
	assign _0229_ = _1389_ & ~_0228_;
	assign _0230_ = _0229_ | _0227_;
	assign _0232_ = _0102_ | _1404_;
	assign _0233_ = _0286_ & ~_0232_;
	assign _0234_ = _0106_ | _1416_;
	assign _0235_ = _0720_ & ~_0234_;
	assign _0236_ = _0235_ | _0233_;
	assign _0237_ = _0112_ | _1430_;
	assign _0238_ = _1089_ & ~_0237_;
	assign _0239_ = _0238_ | _0236_;
	assign _0240_ = _0117_ | _1443_;
	assign _0241_ = _1389_ & ~_0240_;
	assign _0243_ = _0241_ | _0239_;
	assign _0244_ = (\mchip.idx [3] ? _0243_ : _0230_);
	assign _0245_ = (\mchip.idx [4] ? _0244_ : _0218_);
	assign _0246_ = _0124_ | _1404_;
	assign _0247_ = _0286_ & ~_0246_;
	assign _0248_ = _0127_ | _1416_;
	assign _0249_ = _0720_ & ~_0248_;
	assign _0250_ = _0249_ | _0247_;
	assign _0251_ = _0131_ | _1430_;
	assign _0252_ = _1089_ & ~_0251_;
	assign _0254_ = _0252_ | _0250_;
	assign _0255_ = _0136_ | _1443_;
	assign _0256_ = _1389_ & ~_0255_;
	assign _0257_ = _0256_ | _0254_;
	assign _0258_ = _0140_ | _1404_;
	assign _0259_ = _0286_ & ~_0258_;
	assign _0260_ = _0144_ | _1416_;
	assign _0261_ = _0720_ & ~_0260_;
	assign _0262_ = _0261_ | _0259_;
	assign _0263_ = _0148_ | _1430_;
	assign _0265_ = _1089_ & ~_0263_;
	assign _0266_ = _0265_ | _0262_;
	assign _0267_ = _0152_ | _1443_;
	assign _0268_ = _1389_ & ~_0267_;
	assign _0269_ = _0268_ | _0266_;
	assign _0270_ = (\mchip.idx [3] ? _0269_ : _0257_);
	assign _0271_ = _0158_ | _1404_;
	assign _0272_ = _0286_ & ~_0271_;
	assign _0273_ = _0161_ | _1416_;
	assign _0274_ = _0720_ & ~_0273_;
	assign _0276_ = _0274_ | _0272_;
	assign _0277_ = _0166_ | _1430_;
	assign _0278_ = _1089_ & ~_0277_;
	assign _0279_ = _0278_ | _0276_;
	assign _0280_ = _0170_ | _1443_;
	assign _0281_ = _1389_ & ~_0280_;
	assign _0282_ = _0281_ | _0279_;
	assign _0283_ = _0174_ | _1404_;
	assign _0284_ = _0286_ & ~_0283_;
	assign _0285_ = _0178_ | _1416_;
	assign _0287_ = _0720_ & ~_0285_;
	assign _0288_ = _0287_ | _0284_;
	assign _0289_ = _0182_ | _1430_;
	assign _0290_ = _1089_ & ~_0289_;
	assign _0291_ = _0290_ | _0288_;
	assign _0292_ = _0186_ | _1443_;
	assign _0293_ = _1389_ & ~_0292_;
	assign _0294_ = _0293_ | _0291_;
	assign _0295_ = (\mchip.idx [3] ? _0294_ : _0282_);
	assign _0296_ = (\mchip.idx [4] ? _0295_ : _0270_);
	assign _0298_ = (\mchip.idx [5] ? _0296_ : _0245_);
	assign \mchip.iout [3] = (\mchip.idx [6] ? _0298_ : _0193_);
	assign _0299_ = _1409_ | ~_0362_;
	assign _0300_ = _0299_ | ~_0395_;
	assign _0301_ = _0300_ | _1407_;
	assign _0302_ = _0301_ | _1406_;
	assign _0303_ = _0302_ | _1405_;
	assign _0304_ = _0286_ & ~_0303_;
	assign _0305_ = _1422_ | _1739_;
	assign _0306_ = _0305_ | _1420_;
	assign _0308_ = _0306_ | _1419_;
	assign _0309_ = _0308_ | _1418_;
	assign _0310_ = _0309_ | _1417_;
	assign _0311_ = _0720_ & ~_0310_;
	assign _0312_ = _0311_ | _0304_;
	assign _0313_ = _1435_ | ~_1728_;
	assign _0314_ = _0313_ | ~_1151_;
	assign _0315_ = _0314_ | _1433_;
	assign _0316_ = _0315_ | _1432_;
	assign _0317_ = _0316_ | _1431_;
	assign _0319_ = _1089_ & ~_0317_;
	assign _0320_ = _0319_ | _0312_;
	assign _0321_ = _1448_ | _1739_;
	assign _0322_ = _0321_ | _1420_;
	assign _0323_ = _0322_ | _1446_;
	assign _0324_ = _0323_ | _1445_;
	assign _0325_ = _0324_ | _1444_;
	assign _0326_ = _1389_ & ~_0325_;
	assign _0327_ = _0326_ | _0320_;
	assign _0328_ = _0299_ | _0395_;
	assign _0330_ = _0328_ | _1407_;
	assign _0331_ = _0330_ | _1406_;
	assign _0332_ = _0331_ | _1405_;
	assign _0333_ = _0286_ & ~_0332_;
	assign _0334_ = _0305_ | _0731_;
	assign _0335_ = _0334_ | _1419_;
	assign _0336_ = _0335_ | _1418_;
	assign _0337_ = _0336_ | _1417_;
	assign _0338_ = _0720_ & ~_0337_;
	assign _0339_ = _0338_ | _0333_;
	assign _0341_ = _0313_ | _1151_;
	assign _0342_ = _0341_ | _1433_;
	assign _0343_ = _0342_ | _1432_;
	assign _0344_ = _0343_ | _1431_;
	assign _0345_ = _1089_ & ~_0344_;
	assign _0346_ = _0345_ | _0339_;
	assign _0347_ = _0321_ | _0731_;
	assign _0348_ = _0347_ | _1446_;
	assign _0349_ = _0348_ | _1445_;
	assign _0350_ = _0349_ | _1444_;
	assign _0352_ = _1389_ & ~_0350_;
	assign _0353_ = _0352_ | _0346_;
	assign _0354_ = (\mchip.idx [3] ? _0353_ : _0327_);
	assign _0355_ = _0300_ | _0417_;
	assign _0356_ = _0355_ | _1406_;
	assign _0357_ = _0356_ | _1405_;
	assign _0358_ = _0286_ & ~_0357_;
	assign _0359_ = _0306_ | _0808_;
	assign _0360_ = _0359_ | _1418_;
	assign _0361_ = _0360_ | _1417_;
	assign _0363_ = _0720_ & ~_0361_;
	assign _0364_ = _0363_ | _0358_;
	assign _0365_ = _0314_ | _1172_;
	assign _0366_ = _0365_ | _1432_;
	assign _0367_ = _0366_ | _1431_;
	assign _0368_ = _1089_ & ~_0367_;
	assign _0369_ = _0368_ | _0364_;
	assign _0370_ = _0322_ | _1396_;
	assign _0371_ = _0370_ | _1445_;
	assign _0372_ = _0371_ | _1444_;
	assign _0374_ = _1389_ & ~_0372_;
	assign _0375_ = _0374_ | _0369_;
	assign _0376_ = _0328_ | _0417_;
	assign _0377_ = _0376_ | _1406_;
	assign _0378_ = _0377_ | _1405_;
	assign _0379_ = _0286_ & ~_0378_;
	assign _0380_ = _0334_ | _0808_;
	assign _0381_ = _0380_ | _1418_;
	assign _0382_ = _0381_ | _1417_;
	assign _0383_ = _0720_ & ~_0382_;
	assign _0385_ = _0383_ | _0379_;
	assign _0386_ = _0341_ | _1172_;
	assign _0387_ = _0386_ | _1432_;
	assign _0388_ = _0387_ | _1431_;
	assign _0389_ = _1089_ & ~_0388_;
	assign _0390_ = _0389_ | _0385_;
	assign _0391_ = _0347_ | _1396_;
	assign _0392_ = _0391_ | _1445_;
	assign _0393_ = _0392_ | _1444_;
	assign _0394_ = _1389_ & ~_0393_;
	assign _0396_ = _0394_ | _0390_;
	assign _0397_ = (\mchip.idx [3] ? _0396_ : _0375_);
	assign _0398_ = (\mchip.idx [4] ? _0397_ : _0354_);
	assign _0399_ = _0301_ | _0450_;
	assign _0400_ = _0399_ | _1405_;
	assign _0401_ = _0286_ & ~_0400_;
	assign _0402_ = _0308_ | _0841_;
	assign _0403_ = _0402_ | _1417_;
	assign _0404_ = _0720_ & ~_0403_;
	assign _0405_ = _0404_ | _0401_;
	assign _0407_ = _0315_ | _1205_;
	assign _0408_ = _0407_ | _1431_;
	assign _0409_ = _1089_ & ~_0408_;
	assign _0410_ = _0409_ | _0405_;
	assign _0411_ = _0323_ | _1399_;
	assign _0412_ = _0411_ | _1444_;
	assign _0413_ = _1389_ & ~_0412_;
	assign _0414_ = _0413_ | _0410_;
	assign _0415_ = _0330_ | _0450_;
	assign _0416_ = _0415_ | _1405_;
	assign _0418_ = _0286_ & ~_0416_;
	assign _0419_ = _0335_ | _0841_;
	assign _0420_ = _0419_ | _1417_;
	assign _0421_ = _0720_ & ~_0420_;
	assign _0422_ = _0421_ | _0418_;
	assign _0423_ = _0342_ | _1205_;
	assign _0424_ = _0423_ | _1431_;
	assign _0425_ = _1089_ & ~_0424_;
	assign _0426_ = _0425_ | _0422_;
	assign _0427_ = _0348_ | _1399_;
	assign _0429_ = _0427_ | _1444_;
	assign _0430_ = _1389_ & ~_0429_;
	assign _0431_ = _0430_ | _0426_;
	assign _0432_ = (\mchip.idx [3] ? _0431_ : _0414_);
	assign _0433_ = _0355_ | _0450_;
	assign _0434_ = _0433_ | _1405_;
	assign _0435_ = _0286_ & ~_0434_;
	assign _0436_ = _0359_ | _0841_;
	assign _0437_ = _0436_ | _1417_;
	assign _0438_ = _0720_ & ~_0437_;
	assign _0440_ = _0438_ | _0435_;
	assign _0441_ = _0365_ | _1205_;
	assign _0442_ = _0441_ | _1431_;
	assign _0443_ = _1089_ & ~_0442_;
	assign _0444_ = _0443_ | _0440_;
	assign _0445_ = _0370_ | _1399_;
	assign _0446_ = _0445_ | _1444_;
	assign _0447_ = _1389_ & ~_0446_;
	assign _0448_ = _0447_ | _0444_;
	assign _0449_ = _0376_ | _0450_;
	assign _0451_ = _0449_ | _1405_;
	assign _0452_ = _0286_ & ~_0451_;
	assign _0453_ = _0380_ | _0841_;
	assign _0454_ = _0453_ | _1417_;
	assign _0455_ = _0720_ & ~_0454_;
	assign _0456_ = _0455_ | _0452_;
	assign _0457_ = _0386_ | _1205_;
	assign _0458_ = _0457_ | _1431_;
	assign _0459_ = _1089_ & ~_0458_;
	assign _0460_ = _0459_ | _0456_;
	assign _0462_ = _0391_ | _1399_;
	assign _0463_ = _0462_ | _1444_;
	assign _0464_ = _1389_ & ~_0463_;
	assign _0465_ = _0464_ | _0460_;
	assign _0466_ = (\mchip.idx [3] ? _0465_ : _0448_);
	assign _0467_ = (\mchip.idx [4] ? _0466_ : _0432_);
	assign _0468_ = (\mchip.idx [5] ? _0467_ : _0398_);
	assign _0469_ = _0302_ | _1404_;
	assign _0470_ = _0286_ & ~_0469_;
	assign _0471_ = _0309_ | _1416_;
	assign _0473_ = _0720_ & ~_0471_;
	assign _0474_ = _0473_ | _0470_;
	assign _0475_ = _0316_ | _1430_;
	assign _0476_ = _1089_ & ~_0475_;
	assign _0477_ = _0476_ | _0474_;
	assign _0478_ = _0324_ | _1443_;
	assign _0479_ = _1389_ & ~_0478_;
	assign _0480_ = _0479_ | _0477_;
	assign _0481_ = _0331_ | _1404_;
	assign _0482_ = _0286_ & ~_0481_;
	assign _0484_ = _0336_ | _1416_;
	assign _0485_ = _0720_ & ~_0484_;
	assign _0486_ = _0485_ | _0482_;
	assign _0487_ = _0343_ | _1430_;
	assign _0488_ = _1089_ & ~_0487_;
	assign _0489_ = _0488_ | _0486_;
	assign _0490_ = _0349_ | _1443_;
	assign _0491_ = _1389_ & ~_0490_;
	assign _0492_ = _0491_ | _0489_;
	assign _0493_ = (\mchip.idx [3] ? _0492_ : _0480_);
	assign _0495_ = _0356_ | _1404_;
	assign _0496_ = _0286_ & ~_0495_;
	assign _0497_ = _0360_ | _1416_;
	assign _0498_ = _0720_ & ~_0497_;
	assign _0499_ = _0498_ | _0496_;
	assign _0500_ = _0366_ | _1430_;
	assign _0501_ = _1089_ & ~_0500_;
	assign _0502_ = _0501_ | _0499_;
	assign _0503_ = _0371_ | _1443_;
	assign _0504_ = _1389_ & ~_0503_;
	assign _0506_ = _0504_ | _0502_;
	assign _0507_ = _0377_ | _1404_;
	assign _0508_ = _0286_ & ~_0507_;
	assign _0509_ = _0381_ | _1416_;
	assign _0510_ = _0720_ & ~_0509_;
	assign _0511_ = _0510_ | _0508_;
	assign _0512_ = _0387_ | _1430_;
	assign _0513_ = _1089_ & ~_0512_;
	assign _0514_ = _0513_ | _0511_;
	assign _0515_ = _0392_ | _1443_;
	assign _0517_ = _1389_ & ~_0515_;
	assign _0518_ = _0517_ | _0514_;
	assign _0519_ = (\mchip.idx [3] ? _0518_ : _0506_);
	assign _0520_ = (\mchip.idx [4] ? _0519_ : _0493_);
	assign _0521_ = _0399_ | _1404_;
	assign _0522_ = _0286_ & ~_0521_;
	assign _0523_ = _0402_ | _1416_;
	assign _0524_ = _0720_ & ~_0523_;
	assign _0525_ = _0524_ | _0522_;
	assign _0526_ = _0407_ | _1430_;
	assign _0528_ = _1089_ & ~_0526_;
	assign _0529_ = _0528_ | _0525_;
	assign _0530_ = _0411_ | _1443_;
	assign _0531_ = _1389_ & ~_0530_;
	assign _0532_ = _0531_ | _0529_;
	assign _0533_ = _0415_ | _1404_;
	assign _0534_ = _0286_ & ~_0533_;
	assign _0535_ = _0419_ | _1416_;
	assign _0536_ = _0720_ & ~_0535_;
	assign _0537_ = _0536_ | _0534_;
	assign _0539_ = _0423_ | _1430_;
	assign _0540_ = _1089_ & ~_0539_;
	assign _0541_ = _0540_ | _0537_;
	assign _0542_ = _0427_ | _1443_;
	assign _0543_ = _1389_ & ~_0542_;
	assign _0544_ = _0543_ | _0541_;
	assign _0545_ = (\mchip.idx [3] ? _0544_ : _0532_);
	assign _0546_ = _0433_ | _1404_;
	assign _0547_ = _0286_ & ~_0546_;
	assign _0548_ = _0436_ | _1416_;
	assign _0550_ = _0720_ & ~_0548_;
	assign _0551_ = _0550_ | _0547_;
	assign _0552_ = _0441_ | _1430_;
	assign _0553_ = _1089_ & ~_0552_;
	assign _0554_ = _0553_ | _0551_;
	assign _0555_ = _0445_ | _1443_;
	assign _0556_ = _1389_ & ~_0555_;
	assign _0557_ = _0556_ | _0554_;
	assign _0558_ = _0449_ | _1404_;
	assign _0559_ = _0286_ & ~_0558_;
	assign _0561_ = _0453_ | _1416_;
	assign _0562_ = _0720_ & ~_0561_;
	assign _0563_ = _0562_ | _0559_;
	assign _0564_ = _0457_ | _1430_;
	assign _0565_ = _1089_ & ~_0564_;
	assign _0566_ = _0565_ | _0563_;
	assign _0567_ = _0462_ | _1443_;
	assign _0568_ = _1389_ & ~_0567_;
	assign _0569_ = _0568_ | _0566_;
	assign _0570_ = (\mchip.idx [3] ? _0569_ : _0557_);
	assign _0572_ = (\mchip.idx [4] ? _0570_ : _0545_);
	assign _0573_ = (\mchip.idx [5] ? _0572_ : _0520_);
	assign \mchip.iout [4] = (\mchip.idx [6] ? _0573_ : _0468_);
	assign _0574_ = ~(_1681_ & \mchip.x [2]);
	assign _0575_ = _0574_ | ~_0395_;
	assign _0576_ = _0575_ | ~_0417_;
	assign _0577_ = _0576_ | ~_0450_;
	assign _0578_ = _0577_ | ~_1404_;
	assign _0579_ = _0286_ & ~_0578_;
	assign _0580_ = _1678_ | _1728_;
	assign _0582_ = _0580_ | ~_0731_;
	assign _0583_ = _0582_ | ~_0808_;
	assign _0584_ = _0583_ | ~_0841_;
	assign _0585_ = _0584_ | ~_1416_;
	assign _0586_ = _0720_ & ~_0585_;
	assign _0587_ = _0586_ | _0579_;
	assign _0588_ = _0580_ | ~_1151_;
	assign _0589_ = _0588_ | ~_1172_;
	assign _0590_ = _0589_ | ~_1205_;
	assign _0592_ = _0590_ | ~_1430_;
	assign _0593_ = _1089_ & ~_0592_;
	assign _0594_ = _0593_ | _0587_;
	assign _0595_ = _0582_ | ~_1396_;
	assign _0596_ = _0595_ | ~_1399_;
	assign _0597_ = _0596_ | ~_1443_;
	assign _0598_ = _1389_ & ~_0597_;
	assign _0599_ = _0598_ | _0594_;
	assign _0601_ = _0574_ | _0395_;
	assign _0602_ = _0601_ | ~_0417_;
	assign _0603_ = _0602_ | ~_0450_;
	assign _0604_ = _0603_ | ~_1404_;
	assign _0605_ = _0286_ & ~_0604_;
	assign _0606_ = _0580_ | _0731_;
	assign _0607_ = _0606_ | ~_0808_;
	assign _0608_ = _0607_ | ~_0841_;
	assign _0609_ = _0608_ | ~_1416_;
	assign _0610_ = _0720_ & ~_0609_;
	assign _0612_ = _0610_ | _0605_;
	assign _0613_ = _0580_ | _1151_;
	assign _0614_ = _0613_ | ~_1172_;
	assign _0615_ = _0614_ | ~_1205_;
	assign _0616_ = _0615_ | ~_1430_;
	assign _0617_ = _1089_ & ~_0616_;
	assign _0618_ = _0617_ | _0612_;
	assign _0619_ = _0606_ | ~_1396_;
	assign _0620_ = _0619_ | ~_1399_;
	assign _0622_ = _0620_ | ~_1443_;
	assign _0623_ = _1389_ & ~_0622_;
	assign _0624_ = _0623_ | _0618_;
	assign _0625_ = (\mchip.idx [3] ? _0624_ : _0599_);
	assign _0626_ = _0575_ | _0417_;
	assign _0627_ = _0626_ | ~_0450_;
	assign _0628_ = _0627_ | ~_1404_;
	assign _0629_ = _0286_ & ~_0628_;
	assign _0630_ = _0582_ | _0808_;
	assign _0631_ = _0630_ | ~_0841_;
	assign _0633_ = _0631_ | ~_1416_;
	assign _0634_ = _0720_ & ~_0633_;
	assign _0635_ = _0634_ | _0629_;
	assign _0636_ = _0588_ | _1172_;
	assign _0637_ = _0636_ | ~_1205_;
	assign _0638_ = _0637_ | ~_1430_;
	assign _0639_ = _1089_ & ~_0638_;
	assign _0640_ = _0639_ | _0635_;
	assign _0641_ = _0582_ | _1396_;
	assign _0642_ = _0641_ | ~_1399_;
	assign _0644_ = _0642_ | ~_1443_;
	assign _0645_ = _1389_ & ~_0644_;
	assign _0646_ = _0645_ | _0640_;
	assign _0647_ = _0601_ | _0417_;
	assign _0648_ = _0647_ | ~_0450_;
	assign _0649_ = _0648_ | ~_1404_;
	assign _0650_ = _0286_ & ~_0649_;
	assign _0651_ = _0606_ | _0808_;
	assign _0652_ = _0651_ | ~_0841_;
	assign _0653_ = _0652_ | ~_1416_;
	assign _0655_ = _0720_ & ~_0653_;
	assign _0656_ = _0655_ | _0650_;
	assign _0657_ = _0613_ | _1172_;
	assign _0658_ = _0657_ | ~_1205_;
	assign _0659_ = _0658_ | ~_1430_;
	assign _0660_ = _1089_ & ~_0659_;
	assign _0661_ = _0660_ | _0656_;
	assign _0662_ = _0606_ | _1396_;
	assign _0663_ = _0662_ | ~_1399_;
	assign _0664_ = _0663_ | ~_1443_;
	assign _0666_ = _1389_ & ~_0664_;
	assign _0667_ = _0666_ | _0661_;
	assign _0668_ = (\mchip.idx [3] ? _0667_ : _0646_);
	assign _0669_ = (\mchip.idx [4] ? _0668_ : _0625_);
	assign _0670_ = _0576_ | _0450_;
	assign _0671_ = _0670_ | ~_1404_;
	assign _0672_ = _0286_ & ~_0671_;
	assign _0673_ = _0583_ | _0841_;
	assign _0674_ = _0673_ | ~_1416_;
	assign _0675_ = _0720_ & ~_0674_;
	assign _0677_ = _0675_ | _0672_;
	assign _0678_ = _0589_ | _1205_;
	assign _0679_ = _0678_ | ~_1430_;
	assign _0680_ = _1089_ & ~_0679_;
	assign _0681_ = _0680_ | _0677_;
	assign _0682_ = _0595_ | _1399_;
	assign _0683_ = _0682_ | ~_1443_;
	assign _0684_ = _1389_ & ~_0683_;
	assign _0685_ = _0684_ | _0681_;
	assign _0686_ = _0602_ | _0450_;
	assign _0688_ = _0686_ | ~_1404_;
	assign _0689_ = _0286_ & ~_0688_;
	assign _0690_ = _0607_ | _0841_;
	assign _0691_ = _0690_ | ~_1416_;
	assign _0692_ = _0720_ & ~_0691_;
	assign _0693_ = _0692_ | _0689_;
	assign _0694_ = _0614_ | _1205_;
	assign _0695_ = _0694_ | ~_1430_;
	assign _0696_ = _1089_ & ~_0695_;
	assign _0697_ = _0696_ | _0693_;
	assign _0699_ = _0619_ | _1399_;
	assign _0700_ = _0699_ | ~_1443_;
	assign _0701_ = _1389_ & ~_0700_;
	assign _0702_ = _0701_ | _0697_;
	assign _0703_ = (\mchip.idx [3] ? _0702_ : _0685_);
	assign _0704_ = _0626_ | _0450_;
	assign _0705_ = _0704_ | ~_1404_;
	assign _0706_ = _0286_ & ~_0705_;
	assign _0707_ = _0630_ | _0841_;
	assign _0708_ = _0707_ | ~_1416_;
	assign _0710_ = _0720_ & ~_0708_;
	assign _0711_ = _0710_ | _0706_;
	assign _0712_ = _0636_ | _1205_;
	assign _0713_ = _0712_ | ~_1430_;
	assign _0714_ = _1089_ & ~_0713_;
	assign _0715_ = _0714_ | _0711_;
	assign _0716_ = _0641_ | _1399_;
	assign _0717_ = _0716_ | ~_1443_;
	assign _0718_ = _1389_ & ~_0717_;
	assign _0719_ = _0718_ | _0715_;
	assign _0721_ = _0647_ | _0450_;
	assign _0722_ = _0721_ | ~_1404_;
	assign _0723_ = _0286_ & ~_0722_;
	assign _0724_ = _0651_ | _0841_;
	assign _0725_ = _0724_ | ~_1416_;
	assign _0726_ = _0720_ & ~_0725_;
	assign _0727_ = _0726_ | _0723_;
	assign _0728_ = _0657_ | _1205_;
	assign _0729_ = _0728_ | ~_1430_;
	assign _0730_ = _1089_ & ~_0729_;
	assign _0732_ = _0730_ | _0727_;
	assign _0733_ = _0662_ | _1399_;
	assign _0734_ = _0733_ | ~_1443_;
	assign _0735_ = _1389_ & ~_0734_;
	assign _0736_ = _0735_ | _0732_;
	assign _0737_ = (\mchip.idx [3] ? _0736_ : _0719_);
	assign _0738_ = (\mchip.idx [4] ? _0737_ : _0703_);
	assign _0739_ = (\mchip.idx [5] ? _0738_ : _0669_);
	assign _0740_ = _0577_ | _1404_;
	assign _0741_ = _0286_ & ~_0740_;
	assign _0743_ = _0584_ | _1416_;
	assign _0744_ = _0720_ & ~_0743_;
	assign _0745_ = _0744_ | _0741_;
	assign _0746_ = _0590_ | _1430_;
	assign _0747_ = _1089_ & ~_0746_;
	assign _0748_ = _0747_ | _0745_;
	assign _0749_ = _0596_ | _1443_;
	assign _0750_ = _1389_ & ~_0749_;
	assign _0751_ = _0750_ | _0748_;
	assign _0752_ = _0603_ | _1404_;
	assign _0754_ = _0286_ & ~_0752_;
	assign _0755_ = _0608_ | _1416_;
	assign _0756_ = _0720_ & ~_0755_;
	assign _0757_ = _0756_ | _0754_;
	assign _0758_ = _0615_ | _1430_;
	assign _0759_ = _1089_ & ~_0758_;
	assign _0760_ = _0759_ | _0757_;
	assign _0761_ = _0620_ | _1443_;
	assign _0762_ = _1389_ & ~_0761_;
	assign _0763_ = _0762_ | _0760_;
	assign _0765_ = (\mchip.idx [3] ? _0763_ : _0751_);
	assign _0766_ = _0627_ | _1404_;
	assign _0767_ = _0286_ & ~_0766_;
	assign _0768_ = _0631_ | _1416_;
	assign _0769_ = _0720_ & ~_0768_;
	assign _0770_ = _0769_ | _0767_;
	assign _0771_ = _0637_ | _1430_;
	assign _0772_ = _1089_ & ~_0771_;
	assign _0773_ = _0772_ | _0770_;
	assign _0774_ = _0642_ | _1443_;
	assign _0776_ = _1389_ & ~_0774_;
	assign _0777_ = _0776_ | _0773_;
	assign _0778_ = _0648_ | _1404_;
	assign _0779_ = _0286_ & ~_0778_;
	assign _0780_ = _0652_ | _1416_;
	assign _0781_ = _0720_ & ~_0780_;
	assign _0782_ = _0781_ | _0779_;
	assign _0783_ = _0658_ | _1430_;
	assign _0784_ = _1089_ & ~_0783_;
	assign _0785_ = _0784_ | _0782_;
	assign _0787_ = _0663_ | _1443_;
	assign _0788_ = _1389_ & ~_0787_;
	assign _0789_ = _0788_ | _0785_;
	assign _0790_ = (\mchip.idx [3] ? _0789_ : _0777_);
	assign _0791_ = (\mchip.idx [4] ? _0790_ : _0765_);
	assign _0792_ = _0670_ | _1404_;
	assign _0793_ = _0286_ & ~_0792_;
	assign _0794_ = _0673_ | _1416_;
	assign _0795_ = _0720_ & ~_0794_;
	assign _0796_ = _0795_ | _0793_;
	assign _0798_ = _0678_ | _1430_;
	assign _0799_ = _1089_ & ~_0798_;
	assign _0800_ = _0799_ | _0796_;
	assign _0801_ = _0682_ | _1443_;
	assign _0802_ = _1389_ & ~_0801_;
	assign _0803_ = _0802_ | _0800_;
	assign _0804_ = _0686_ | _1404_;
	assign _0805_ = _0286_ & ~_0804_;
	assign _0806_ = _0690_ | _1416_;
	assign _0807_ = _0720_ & ~_0806_;
	assign _0809_ = _0807_ | _0805_;
	assign _0810_ = _0694_ | _1430_;
	assign _0811_ = _1089_ & ~_0810_;
	assign _0812_ = _0811_ | _0809_;
	assign _0813_ = _0699_ | _1443_;
	assign _0814_ = _1389_ & ~_0813_;
	assign _0815_ = _0814_ | _0812_;
	assign _0816_ = (\mchip.idx [3] ? _0815_ : _0803_);
	assign _0817_ = _0704_ | _1404_;
	assign _0818_ = _0286_ & ~_0817_;
	assign _0820_ = _0707_ | _1416_;
	assign _0821_ = _0720_ & ~_0820_;
	assign _0822_ = _0821_ | _0818_;
	assign _0823_ = _0712_ | _1430_;
	assign _0824_ = _1089_ & ~_0823_;
	assign _0825_ = _0824_ | _0822_;
	assign _0826_ = _0716_ | _1443_;
	assign _0827_ = _1389_ & ~_0826_;
	assign _0828_ = _0827_ | _0825_;
	assign _0829_ = _0721_ | _1404_;
	assign _0831_ = _0286_ & ~_0829_;
	assign _0832_ = _0724_ | _1416_;
	assign _0833_ = _0720_ & ~_0832_;
	assign _0834_ = _0833_ | _0831_;
	assign _0835_ = _0728_ | _1430_;
	assign _0836_ = _1089_ & ~_0835_;
	assign _0837_ = _0836_ | _0834_;
	assign _0838_ = _0733_ | _1443_;
	assign _0839_ = _1389_ & ~_0838_;
	assign _0840_ = _0839_ | _0837_;
	assign _0842_ = (\mchip.idx [3] ? _0840_ : _0828_);
	assign _0843_ = (\mchip.idx [4] ? _0842_ : _0816_);
	assign _0844_ = (\mchip.idx [5] ? _0843_ : _0791_);
	assign \mchip.iout [5] = (\mchip.idx [6] ? _0844_ : _0739_);
	assign _0845_ = _1678_ | _0362_;
	assign _0846_ = _0845_ | ~_0395_;
	assign _0847_ = _0846_ | ~_0417_;
	assign _0848_ = _0847_ | ~_0450_;
	assign _0849_ = _0848_ | ~_1404_;
	assign _0850_ = _0286_ & ~_0849_;
	assign _0852_ = _1945_ | _1728_;
	assign _0853_ = _0852_ | ~_0731_;
	assign _0854_ = _0853_ | ~_0808_;
	assign _0855_ = _0854_ | ~_0841_;
	assign _0856_ = _0855_ | ~_1416_;
	assign _0857_ = _0720_ & ~_0856_;
	assign _0858_ = _0857_ | _0850_;
	assign _0859_ = _0852_ | ~_1151_;
	assign _0860_ = _0859_ | ~_1172_;
	assign _0862_ = _0860_ | ~_1205_;
	assign _0863_ = _0862_ | ~_1430_;
	assign _0864_ = _1089_ & ~_0863_;
	assign _0865_ = _0864_ | _0858_;
	assign _0866_ = _0853_ | ~_1396_;
	assign _0867_ = _0866_ | ~_1399_;
	assign _0868_ = _0867_ | ~_1443_;
	assign _0869_ = _1389_ & ~_0868_;
	assign _0871_ = _0869_ | _0865_;
	assign _0872_ = _0845_ | _0395_;
	assign _0873_ = _0872_ | ~_0417_;
	assign _0874_ = _0873_ | ~_0450_;
	assign _0875_ = _0874_ | ~_1404_;
	assign _0876_ = _0286_ & ~_0875_;
	assign _0877_ = _0852_ | _0731_;
	assign _0878_ = _0877_ | ~_0808_;
	assign _0879_ = _0878_ | ~_0841_;
	assign _0880_ = _0879_ | ~_1416_;
	assign _0882_ = _0720_ & ~_0880_;
	assign _0883_ = _0882_ | _0876_;
	assign _0884_ = _0852_ | _1151_;
	assign _0885_ = _0884_ | ~_1172_;
	assign _0886_ = _0885_ | ~_1205_;
	assign _0887_ = _0886_ | ~_1430_;
	assign _0888_ = _1089_ & ~_0887_;
	assign _0889_ = _0888_ | _0883_;
	assign _0890_ = _0877_ | ~_1396_;
	assign _0892_ = _0890_ | ~_1399_;
	assign _0893_ = _0892_ | ~_1443_;
	assign _0894_ = _1389_ & ~_0893_;
	assign _0895_ = _0894_ | _0889_;
	assign _0896_ = (\mchip.idx [3] ? _0895_ : _0871_);
	assign _0897_ = _0846_ | _0417_;
	assign _0898_ = _0897_ | ~_0450_;
	assign _0899_ = _0898_ | ~_1404_;
	assign _0900_ = _0286_ & ~_0899_;
	assign _0901_ = _0853_ | _0808_;
	assign _0903_ = _0901_ | ~_0841_;
	assign _0904_ = _0903_ | ~_1416_;
	assign _0905_ = _0720_ & ~_0904_;
	assign _0906_ = _0905_ | _0900_;
	assign _0907_ = _0859_ | _1172_;
	assign _0908_ = _0907_ | ~_1205_;
	assign _0909_ = _0908_ | ~_1430_;
	assign _0910_ = _1089_ & ~_0909_;
	assign _0911_ = _0910_ | _0906_;
	assign _0912_ = _0853_ | _1396_;
	assign _0914_ = _0912_ | ~_1399_;
	assign _0915_ = _0914_ | ~_1443_;
	assign _0916_ = _1389_ & ~_0915_;
	assign _0917_ = _0916_ | _0911_;
	assign _0918_ = _0872_ | _0417_;
	assign _0919_ = _0918_ | ~_0450_;
	assign _0920_ = _0919_ | ~_1404_;
	assign _0921_ = _0286_ & ~_0920_;
	assign _0922_ = _0877_ | _0808_;
	assign _0923_ = _0922_ | ~_0841_;
	assign _0925_ = _0923_ | ~_1416_;
	assign _0926_ = _0720_ & ~_0925_;
	assign _0927_ = _0926_ | _0921_;
	assign _0928_ = _0884_ | _1172_;
	assign _0929_ = _0928_ | ~_1205_;
	assign _0930_ = _0929_ | ~_1430_;
	assign _0931_ = _1089_ & ~_0930_;
	assign _0932_ = _0931_ | _0927_;
	assign _0933_ = _0877_ | _1396_;
	assign _0934_ = _0933_ | ~_1399_;
	assign _0936_ = _0934_ | ~_1443_;
	assign _0937_ = _1389_ & ~_0936_;
	assign _0938_ = _0937_ | _0932_;
	assign _0939_ = (\mchip.idx [3] ? _0938_ : _0917_);
	assign _0940_ = (\mchip.idx [4] ? _0939_ : _0896_);
	assign _0941_ = _0847_ | _0450_;
	assign _0942_ = _0941_ | ~_1404_;
	assign _0943_ = _0286_ & ~_0942_;
	assign _0944_ = _0854_ | _0841_;
	assign _0945_ = _0944_ | ~_1416_;
	assign _0947_ = _0720_ & ~_0945_;
	assign _0948_ = _0947_ | _0943_;
	assign _0949_ = _0860_ | _1205_;
	assign _0950_ = _0949_ | ~_1430_;
	assign _0951_ = _1089_ & ~_0950_;
	assign _0952_ = _0951_ | _0948_;
	assign _0953_ = _0866_ | _1399_;
	assign _0954_ = _0953_ | ~_1443_;
	assign _0955_ = _1389_ & ~_0954_;
	assign _0956_ = _0955_ | _0952_;
	assign _0958_ = _0873_ | _0450_;
	assign _0959_ = _0958_ | ~_1404_;
	assign _0960_ = _0286_ & ~_0959_;
	assign _0961_ = _0878_ | _0841_;
	assign _0962_ = _0961_ | ~_1416_;
	assign _0963_ = _0720_ & ~_0962_;
	assign _0964_ = _0963_ | _0960_;
	assign _0965_ = _0885_ | _1205_;
	assign _0966_ = _0965_ | ~_1430_;
	assign _0967_ = _1089_ & ~_0966_;
	assign _0969_ = _0967_ | _0964_;
	assign _0970_ = _0890_ | _1399_;
	assign _0971_ = _0970_ | ~_1443_;
	assign _0972_ = _1389_ & ~_0971_;
	assign _0973_ = _0972_ | _0969_;
	assign _0974_ = (\mchip.idx [3] ? _0973_ : _0956_);
	assign _0975_ = _0897_ | _0450_;
	assign _0976_ = _0975_ | ~_1404_;
	assign _0977_ = _0286_ & ~_0976_;
	assign _0978_ = _0901_ | _0841_;
	assign _0980_ = _0978_ | ~_1416_;
	assign _0981_ = _0720_ & ~_0980_;
	assign _0982_ = _0981_ | _0977_;
	assign _0983_ = _0907_ | _1205_;
	assign _0984_ = _0983_ | ~_1430_;
	assign _0985_ = _1089_ & ~_0984_;
	assign _0986_ = _0985_ | _0982_;
	assign _0987_ = _0912_ | _1399_;
	assign _0988_ = _0987_ | ~_1443_;
	assign _0989_ = _1389_ & ~_0988_;
	assign _0991_ = _0989_ | _0986_;
	assign _0992_ = _0918_ | _0450_;
	assign _0993_ = _0992_ | ~_1404_;
	assign _0994_ = _0286_ & ~_0993_;
	assign _0995_ = _0922_ | _0841_;
	assign _0996_ = _0995_ | ~_1416_;
	assign _0997_ = _0720_ & ~_0996_;
	assign _0998_ = _0997_ | _0994_;
	assign _0999_ = _0928_ | _1205_;
	assign _1000_ = _0999_ | ~_1430_;
	assign _1002_ = _1089_ & ~_1000_;
	assign _1003_ = _1002_ | _0998_;
	assign _1004_ = _0933_ | _1399_;
	assign _1005_ = _1004_ | ~_1443_;
	assign _1006_ = _1389_ & ~_1005_;
	assign _1007_ = _1006_ | _1003_;
	assign _1008_ = (\mchip.idx [3] ? _1007_ : _0991_);
	assign _1009_ = (\mchip.idx [4] ? _1008_ : _0974_);
	assign _1010_ = (\mchip.idx [5] ? _1009_ : _0940_);
	assign _1011_ = _0848_ | _1404_;
	assign _1013_ = _0286_ & ~_1011_;
	assign _1014_ = _0855_ | _1416_;
	assign _1015_ = _0720_ & ~_1014_;
	assign _1016_ = _1015_ | _1013_;
	assign _1017_ = _0862_ | _1430_;
	assign _1018_ = _1089_ & ~_1017_;
	assign _1019_ = _1018_ | _1016_;
	assign _1020_ = _0867_ | _1443_;
	assign _1021_ = _1389_ & ~_1020_;
	assign _1022_ = _1021_ | _1019_;
	assign _1024_ = _0874_ | _1404_;
	assign _1025_ = _0286_ & ~_1024_;
	assign _1026_ = _0879_ | _1416_;
	assign _1027_ = _0720_ & ~_1026_;
	assign _1028_ = _1027_ | _1025_;
	assign _1029_ = _0886_ | _1430_;
	assign _1030_ = _1089_ & ~_1029_;
	assign _1031_ = _1030_ | _1028_;
	assign _1032_ = _0892_ | _1443_;
	assign _1033_ = _1389_ & ~_1032_;
	assign _1035_ = _1033_ | _1031_;
	assign _1036_ = (\mchip.idx [3] ? _1035_ : _1022_);
	assign _1037_ = _0898_ | _1404_;
	assign _1038_ = _0286_ & ~_1037_;
	assign _1039_ = _0903_ | _1416_;
	assign _1040_ = _0720_ & ~_1039_;
	assign _1041_ = _1040_ | _1038_;
	assign _1042_ = _0908_ | _1430_;
	assign _1043_ = _1089_ & ~_1042_;
	assign _1044_ = _1043_ | _1041_;
	assign _1046_ = _0914_ | _1443_;
	assign _1047_ = _1389_ & ~_1046_;
	assign _1048_ = _1047_ | _1044_;
	assign _1049_ = _0919_ | _1404_;
	assign _1050_ = _0286_ & ~_1049_;
	assign _1051_ = _0923_ | _1416_;
	assign _1052_ = _0720_ & ~_1051_;
	assign _1053_ = _1052_ | _1050_;
	assign _1054_ = _0929_ | _1430_;
	assign _1055_ = _1089_ & ~_1054_;
	assign _1057_ = _1055_ | _1053_;
	assign _1058_ = _0934_ | _1443_;
	assign _1059_ = _1389_ & ~_1058_;
	assign _1060_ = _1059_ | _1057_;
	assign _1061_ = (\mchip.idx [3] ? _1060_ : _1048_);
	assign _1062_ = (\mchip.idx [4] ? _1061_ : _1036_);
	assign _1063_ = _0941_ | _1404_;
	assign _1064_ = _0286_ & ~_1063_;
	assign _1065_ = _0944_ | _1416_;
	assign _1066_ = _0720_ & ~_1065_;
	assign _1068_ = _1066_ | _1064_;
	assign _1069_ = _0949_ | _1430_;
	assign _1070_ = _1089_ & ~_1069_;
	assign _1071_ = _1070_ | _1068_;
	assign _1072_ = _0953_ | _1443_;
	assign _1073_ = _1389_ & ~_1072_;
	assign _1074_ = _1073_ | _1071_;
	assign _1075_ = _0958_ | _1404_;
	assign _1076_ = _0286_ & ~_1075_;
	assign _1077_ = _0961_ | _1416_;
	assign _1079_ = _0720_ & ~_1077_;
	assign _1080_ = _1079_ | _1076_;
	assign _1081_ = _0965_ | _1430_;
	assign _1082_ = _1089_ & ~_1081_;
	assign _1083_ = _1082_ | _1080_;
	assign _1084_ = _0970_ | _1443_;
	assign _1085_ = _1389_ & ~_1084_;
	assign _1086_ = _1085_ | _1083_;
	assign _1087_ = (\mchip.idx [3] ? _1086_ : _1074_);
	assign _1088_ = _0975_ | _1404_;
	assign _1090_ = _0286_ & ~_1088_;
	assign _1091_ = _0978_ | _1416_;
	assign _1092_ = _0720_ & ~_1091_;
	assign _1093_ = _1092_ | _1090_;
	assign _1094_ = _0983_ | _1430_;
	assign _1095_ = _1089_ & ~_1094_;
	assign _1096_ = _1095_ | _1093_;
	assign _1097_ = _0987_ | _1443_;
	assign _1098_ = _1389_ & ~_1097_;
	assign _1099_ = _1098_ | _1096_;
	assign _1101_ = _0992_ | _1404_;
	assign _1102_ = _0286_ & ~_1101_;
	assign _1103_ = _0995_ | _1416_;
	assign _1104_ = _0720_ & ~_1103_;
	assign _1105_ = _1104_ | _1102_;
	assign _1106_ = _0999_ | _1430_;
	assign _1107_ = _1089_ & ~_1106_;
	assign _1108_ = _1107_ | _1105_;
	assign _1109_ = _1004_ | _1443_;
	assign _1110_ = _1389_ & ~_1109_;
	assign _1112_ = _1110_ | _1108_;
	assign _1113_ = (\mchip.idx [3] ? _1112_ : _1099_);
	assign _1114_ = (\mchip.idx [4] ? _1113_ : _1087_);
	assign _1115_ = (\mchip.idx [5] ? _1114_ : _1062_);
	assign \mchip.iout [6] = (\mchip.idx [6] ? _1115_ : _1010_);
	assign _1116_ = _1945_ | _0362_;
	assign _1117_ = _1116_ | ~_0395_;
	assign _1118_ = _1117_ | ~_0417_;
	assign _1119_ = _1118_ | ~_0450_;
	assign _1120_ = _1119_ | ~_1404_;
	assign _1122_ = _0286_ & ~_1120_;
	assign _1123_ = _0033_ | _1728_;
	assign _1124_ = _1123_ | ~_0731_;
	assign _1125_ = _1124_ | ~_0808_;
	assign _1126_ = _1125_ | ~_0841_;
	assign _1127_ = _1126_ | ~_1416_;
	assign _1128_ = _0720_ & ~_1127_;
	assign _1129_ = _1128_ | _1122_;
	assign _1130_ = _1123_ | ~_1151_;
	assign _1132_ = _1130_ | ~_1172_;
	assign _1133_ = _1132_ | ~_1205_;
	assign _1134_ = _1133_ | ~_1430_;
	assign _1135_ = _1089_ & ~_1134_;
	assign _1136_ = _1135_ | _1129_;
	assign _1137_ = _1124_ | ~_1396_;
	assign _1138_ = _1137_ | ~_1399_;
	assign _1139_ = _1138_ | ~_1443_;
	assign _1141_ = _1389_ & ~_1139_;
	assign _1142_ = _1141_ | _1136_;
	assign _1143_ = _1116_ | _0395_;
	assign _1144_ = _1143_ | ~_0417_;
	assign _1145_ = _1144_ | ~_0450_;
	assign _1146_ = _1145_ | ~_1404_;
	assign _1147_ = _0286_ & ~_1146_;
	assign _1148_ = _1123_ | _0731_;
	assign _1149_ = _1148_ | ~_0808_;
	assign _1150_ = _1149_ | ~_0841_;
	assign _1152_ = _1150_ | ~_1416_;
	assign _1153_ = _0720_ & ~_1152_;
	assign _1154_ = _1153_ | _1147_;
	assign _1155_ = _1123_ | _1151_;
	assign _1156_ = _1155_ | ~_1172_;
	assign _1157_ = _1156_ | ~_1205_;
	assign _1158_ = _1157_ | ~_1430_;
	assign _1159_ = _1089_ & ~_1158_;
	assign _1160_ = _1159_ | _1154_;
	assign _1162_ = _1148_ | ~_1396_;
	assign _1163_ = _1162_ | ~_1399_;
	assign _1164_ = _1163_ | ~_1443_;
	assign _1165_ = _1389_ & ~_1164_;
	assign _1166_ = _1165_ | _1160_;
	assign _1167_ = (\mchip.idx [3] ? _1166_ : _1142_);
	assign _1168_ = _1117_ | _0417_;
	assign _1169_ = _1168_ | ~_0450_;
	assign _1170_ = _1169_ | ~_1404_;
	assign _1171_ = _0286_ & ~_1170_;
	assign _1173_ = _1124_ | _0808_;
	assign _1174_ = _1173_ | ~_0841_;
	assign _1175_ = _1174_ | ~_1416_;
	assign _1176_ = _0720_ & ~_1175_;
	assign _1177_ = _1176_ | _1171_;
	assign _1178_ = _1130_ | _1172_;
	assign _1179_ = _1178_ | ~_1205_;
	assign _1180_ = _1179_ | ~_1430_;
	assign _1181_ = _1089_ & ~_1180_;
	assign _1182_ = _1181_ | _1177_;
	assign _1184_ = _1124_ | _1396_;
	assign _1185_ = _1184_ | ~_1399_;
	assign _1186_ = _1185_ | ~_1443_;
	assign _1187_ = _1389_ & ~_1186_;
	assign _1188_ = _1187_ | _1182_;
	assign _1189_ = _1143_ | _0417_;
	assign _1190_ = _1189_ | ~_0450_;
	assign _1191_ = _1190_ | ~_1404_;
	assign _1192_ = _0286_ & ~_1191_;
	assign _1193_ = _1148_ | _0808_;
	assign _1195_ = _1193_ | ~_0841_;
	assign _1196_ = _1195_ | ~_1416_;
	assign _1197_ = _0720_ & ~_1196_;
	assign _1198_ = _1197_ | _1192_;
	assign _1199_ = _1155_ | _1172_;
	assign _1200_ = _1199_ | ~_1205_;
	assign _1201_ = _1200_ | ~_1430_;
	assign _1202_ = _1089_ & ~_1201_;
	assign _1203_ = _1202_ | _1198_;
	assign _1204_ = _1148_ | _1396_;
	assign _1206_ = _1204_ | ~_1399_;
	assign _1207_ = _1206_ | ~_1443_;
	assign _1208_ = _1389_ & ~_1207_;
	assign _1209_ = _1208_ | _1203_;
	assign _1210_ = (\mchip.idx [3] ? _1209_ : _1188_);
	assign _1211_ = (\mchip.idx [4] ? _1210_ : _1167_);
	assign _1212_ = _1118_ | _0450_;
	assign _1213_ = _1212_ | ~_1404_;
	assign _1214_ = _0286_ & ~_1213_;
	assign _1215_ = _1125_ | _0841_;
	assign _1217_ = _1215_ | ~_1416_;
	assign _1218_ = _0720_ & ~_1217_;
	assign _1219_ = _1218_ | _1214_;
	assign _1220_ = _1132_ | _1205_;
	assign _1221_ = _1220_ | ~_1430_;
	assign _1222_ = _1089_ & ~_1221_;
	assign _1223_ = _1222_ | _1219_;
	assign _1224_ = _1137_ | _1399_;
	assign _1225_ = _1224_ | ~_1443_;
	assign _1226_ = _1389_ & ~_1225_;
	assign _1228_ = _1226_ | _1223_;
	assign _1229_ = _1144_ | _0450_;
	assign _1230_ = _1229_ | ~_1404_;
	assign _1231_ = _0286_ & ~_1230_;
	assign _1232_ = _1149_ | _0841_;
	assign _1233_ = _1232_ | ~_1416_;
	assign _1234_ = _0720_ & ~_1233_;
	assign _1235_ = _1234_ | _1231_;
	assign _1236_ = _1156_ | _1205_;
	assign _1237_ = _1236_ | ~_1430_;
	assign _1239_ = _1089_ & ~_1237_;
	assign _1240_ = _1239_ | _1235_;
	assign _1241_ = _1162_ | _1399_;
	assign _1242_ = _1241_ | ~_1443_;
	assign _1243_ = _1389_ & ~_1242_;
	assign _1244_ = _1243_ | _1240_;
	assign _1245_ = (\mchip.idx [3] ? _1244_ : _1228_);
	assign _1246_ = _1168_ | _0450_;
	assign _1247_ = _1246_ | ~_1404_;
	assign _1248_ = _0286_ & ~_1247_;
	assign _1250_ = _1173_ | _0841_;
	assign _1251_ = _1250_ | ~_1416_;
	assign _1252_ = _0720_ & ~_1251_;
	assign _1253_ = _1252_ | _1248_;
	assign _1254_ = _1178_ | _1205_;
	assign _1255_ = _1254_ | ~_1430_;
	assign _1256_ = _1089_ & ~_1255_;
	assign _1257_ = _1256_ | _1253_;
	assign _1258_ = _1184_ | _1399_;
	assign _1259_ = _1258_ | ~_1443_;
	assign _1261_ = _1389_ & ~_1259_;
	assign _1262_ = _1261_ | _1257_;
	assign _1263_ = _1189_ | _0450_;
	assign _1264_ = _1263_ | ~_1404_;
	assign _1265_ = _0286_ & ~_1264_;
	assign _1266_ = _1193_ | _0841_;
	assign _1267_ = _1266_ | ~_1416_;
	assign _1268_ = _0720_ & ~_1267_;
	assign _1269_ = _1268_ | _1265_;
	assign _1270_ = _1199_ | _1205_;
	assign _1272_ = _1270_ | ~_1430_;
	assign _1273_ = _1089_ & ~_1272_;
	assign _1274_ = _1273_ | _1269_;
	assign _1275_ = _1204_ | _1399_;
	assign _1276_ = _1275_ | ~_1443_;
	assign _1277_ = _1389_ & ~_1276_;
	assign _1278_ = _1277_ | _1274_;
	assign _1279_ = (\mchip.idx [3] ? _1278_ : _1262_);
	assign _1280_ = (\mchip.idx [4] ? _1279_ : _1245_);
	assign _1281_ = (\mchip.idx [5] ? _1280_ : _1211_);
	assign _1282_ = _1119_ | _1404_;
	assign _1283_ = _0286_ & ~_1282_;
	assign _1284_ = _1126_ | _1416_;
	assign _1285_ = _0720_ & ~_1284_;
	assign _1286_ = _1285_ | _1283_;
	assign _1287_ = _1133_ | _1430_;
	assign _1288_ = _1089_ & ~_1287_;
	assign _1289_ = _1288_ | _1286_;
	assign _1290_ = _1138_ | _1443_;
	assign _1291_ = _1389_ & ~_1290_;
	assign _1293_ = _1291_ | _1289_;
	assign _1294_ = _1145_ | _1404_;
	assign _1295_ = _0286_ & ~_1294_;
	assign _1296_ = _1150_ | _1416_;
	assign _1297_ = _0720_ & ~_1296_;
	assign _1298_ = _1297_ | _1295_;
	assign _1299_ = _1157_ | _1430_;
	assign _1300_ = _1089_ & ~_1299_;
	assign _1301_ = _1300_ | _1298_;
	assign _1302_ = _1163_ | _1443_;
	assign _1304_ = _1389_ & ~_1302_;
	assign _1305_ = _1304_ | _1301_;
	assign _1306_ = (\mchip.idx [3] ? _1305_ : _1293_);
	assign _1307_ = _1169_ | _1404_;
	assign _1308_ = _0286_ & ~_1307_;
	assign _1309_ = _1174_ | _1416_;
	assign _1310_ = _0720_ & ~_1309_;
	assign _1311_ = _1310_ | _1308_;
	assign _1312_ = _1179_ | _1430_;
	assign _1313_ = _1089_ & ~_1312_;
	assign _1315_ = _1313_ | _1311_;
	assign _1316_ = _1185_ | _1443_;
	assign _1317_ = _1389_ & ~_1316_;
	assign _1318_ = _1317_ | _1315_;
	assign _1319_ = _1190_ | _1404_;
	assign _1320_ = _0286_ & ~_1319_;
	assign _1321_ = _1195_ | _1416_;
	assign _1322_ = _0720_ & ~_1321_;
	assign _1323_ = _1322_ | _1320_;
	assign _1324_ = _1200_ | _1430_;
	assign _1326_ = _1089_ & ~_1324_;
	assign _1327_ = _1326_ | _1323_;
	assign _1328_ = _1206_ | _1443_;
	assign _1329_ = _1389_ & ~_1328_;
	assign _1330_ = _1329_ | _1327_;
	assign _1331_ = (\mchip.idx [3] ? _1330_ : _1318_);
	assign _1332_ = (\mchip.idx [4] ? _1331_ : _1306_);
	assign _1333_ = _1212_ | _1404_;
	assign _1334_ = _0286_ & ~_1333_;
	assign _1335_ = _1215_ | _1416_;
	assign _1337_ = _0720_ & ~_1335_;
	assign _1338_ = _1337_ | _1334_;
	assign _1339_ = _1220_ | _1430_;
	assign _1340_ = _1089_ & ~_1339_;
	assign _1341_ = _1340_ | _1338_;
	assign _1342_ = _1224_ | _1443_;
	assign _1343_ = _1389_ & ~_1342_;
	assign _1344_ = _1343_ | _1341_;
	assign _1345_ = _1229_ | _1404_;
	assign _1346_ = _0286_ & ~_1345_;
	assign _1348_ = _1232_ | _1416_;
	assign _1349_ = _0720_ & ~_1348_;
	assign _1350_ = _1349_ | _1346_;
	assign _1351_ = _1236_ | _1430_;
	assign _1352_ = _1089_ & ~_1351_;
	assign _1353_ = _1352_ | _1350_;
	assign _1354_ = _1241_ | _1443_;
	assign _1355_ = _1389_ & ~_1354_;
	assign _1356_ = _1355_ | _1353_;
	assign _1357_ = (\mchip.idx [3] ? _1356_ : _1344_);
	assign _1359_ = _1246_ | _1404_;
	assign _1360_ = _0286_ & ~_1359_;
	assign _1361_ = _1250_ | _1416_;
	assign _1362_ = _0720_ & ~_1361_;
	assign _1363_ = _1362_ | _1360_;
	assign _1364_ = _1254_ | _1430_;
	assign _1365_ = _1089_ & ~_1364_;
	assign _1366_ = _1365_ | _1363_;
	assign _1367_ = _1258_ | _1443_;
	assign _1368_ = _1389_ & ~_1367_;
	assign _1370_ = _1368_ | _1366_;
	assign _1371_ = _1263_ | _1404_;
	assign _1372_ = _0286_ & ~_1371_;
	assign _1373_ = _1266_ | _1416_;
	assign _1374_ = _0720_ & ~_1373_;
	assign _1375_ = _1374_ | _1372_;
	assign _1376_ = _1270_ | _1430_;
	assign _1377_ = _1089_ & ~_1376_;
	assign _1378_ = _1377_ | _1375_;
	assign _1379_ = _1275_ | _1443_;
	assign _1381_ = _1389_ & ~_1379_;
	assign _1382_ = _1381_ | _1378_;
	assign _1383_ = (\mchip.idx [3] ? _1382_ : _1370_);
	assign _1384_ = (\mchip.idx [4] ? _1383_ : _1357_);
	assign _1385_ = (\mchip.idx [5] ? _1384_ : _1332_);
	assign \mchip.iout [7] = (\mchip.idx [6] ? _1385_ : _1281_);
	reg \mchip.idx_reg[3] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.idx_reg[3]  <= 1'h0;
		else if (io_in[0])
			\mchip.idx_reg[3]  <= _2184_[0];
	assign \mchip.idx [3] = \mchip.idx_reg[3] ;
	reg \mchip.idx_reg[4] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.idx_reg[4]  <= 1'h0;
		else if (io_in[0])
			\mchip.idx_reg[4]  <= _2185_[1];
	assign \mchip.idx [4] = \mchip.idx_reg[4] ;
	reg \mchip.idx_reg[5] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.idx_reg[5]  <= 1'h0;
		else if (io_in[0])
			\mchip.idx_reg[5]  <= _2185_[2];
	assign \mchip.idx [5] = \mchip.idx_reg[5] ;
	reg \mchip.idx_reg[6] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.idx_reg[6]  <= 1'h0;
		else if (io_in[0])
			\mchip.idx_reg[6]  <= _2185_[3];
	assign \mchip.idx [6] = \mchip.idx_reg[6] ;
	reg \mchip.y_reg[0] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.y_reg[0]  <= 1'h0;
		else
			\mchip.y_reg[0]  <= _2182_[0];
	assign \mchip.y [0] = \mchip.y_reg[0] ;
	reg \mchip.y_reg[1] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.y_reg[1]  <= 1'h0;
		else
			\mchip.y_reg[1]  <= _2183_[1];
	assign \mchip.y [1] = \mchip.y_reg[1] ;
	reg \mchip.y_reg[2] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.y_reg[2]  <= 1'h0;
		else
			\mchip.y_reg[2]  <= _2183_[2];
	assign \mchip.y [2] = \mchip.y_reg[2] ;
	reg \mchip.y_reg[3] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.y_reg[3]  <= 1'h0;
		else
			\mchip.y_reg[3]  <= _2183_[3];
	assign \mchip.y [3] = \mchip.y_reg[3] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.x [0] <= 1'h0;
		else if (_0000_)
			\mchip.x [0] <= _0002_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.x [1] <= 1'h0;
		else if (_0000_)
			\mchip.x [1] <= _0003_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.x [2] <= 1'h0;
		else if (_0000_)
			\mchip.x [2] <= _0004_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.x [3] <= 1'h0;
		else if (_0000_)
			\mchip.x [3] <= _0005_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.x [4] <= 1'h0;
		else if (_0000_)
			\mchip.x [4] <= _0006_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.x [5] <= 1'h0;
		else if (_0000_)
			\mchip.x [5] <= _0007_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.x [6] <= 1'h0;
		else if (_0000_)
			\mchip.x [6] <= _0008_;
	reg \mchip.io_out_reg[0] ;
	always @(posedge io_in[12])
		if (_0001_)
			\mchip.io_out_reg[0]  <= \mchip.iout [0];
	assign \mchip.io_out [0] = \mchip.io_out_reg[0] ;
	reg \mchip.io_out_reg[1] ;
	always @(posedge io_in[12])
		if (_0001_)
			\mchip.io_out_reg[1]  <= \mchip.iout [1];
	assign \mchip.io_out [1] = \mchip.io_out_reg[1] ;
	reg \mchip.io_out_reg[2] ;
	always @(posedge io_in[12])
		if (_0001_)
			\mchip.io_out_reg[2]  <= \mchip.iout [2];
	assign \mchip.io_out [2] = \mchip.io_out_reg[2] ;
	reg \mchip.io_out_reg[3] ;
	always @(posedge io_in[12])
		if (_0001_)
			\mchip.io_out_reg[3]  <= \mchip.iout [3];
	assign \mchip.io_out [3] = \mchip.io_out_reg[3] ;
	reg \mchip.io_out_reg[4] ;
	always @(posedge io_in[12])
		if (_0001_)
			\mchip.io_out_reg[4]  <= \mchip.iout [4];
	assign \mchip.io_out [4] = \mchip.io_out_reg[4] ;
	reg \mchip.io_out_reg[5] ;
	always @(posedge io_in[12])
		if (_0001_)
			\mchip.io_out_reg[5]  <= \mchip.iout [5];
	assign \mchip.io_out [5] = \mchip.io_out_reg[5] ;
	reg \mchip.io_out_reg[6] ;
	always @(posedge io_in[12])
		if (_0001_)
			\mchip.io_out_reg[6]  <= \mchip.iout [6];
	assign \mchip.io_out [6] = \mchip.io_out_reg[6] ;
	reg \mchip.io_out_reg[7] ;
	always @(posedge io_in[12])
		if (_0001_)
			\mchip.io_out_reg[7]  <= \mchip.iout [7];
	assign \mchip.io_out [7] = \mchip.io_out_reg[7] ;
	assign _2182_[6:1] = {3'h0, \mchip.y [3:1]};
	assign {_2183_[6:4], _2183_[0]} = {3'h0, _2182_[0]};
	assign _2184_[3:1] = \mchip.idx [6:4];
	assign _2185_[0] = _2184_[0];
	assign io_out = {6'h00, \mchip.io_out [7:0]};
	assign \mchip.clk  = io_in[12];
	assign \mchip.clock  = io_in[12];
	assign \mchip.fallen_state  = 128'h00000000000000000000000000000000;
	assign \mchip.idx [2:0] = 3'h0;
	assign \mchip.io_in  = io_in[11:0];
	assign \mchip.io_out [11:8] = 4'h0;
	assign \mchip.left  = io_in[2];
	assign \mchip.rand_piece  = 16'h0126;
	assign \mchip.read_gs  = io_in[0];
	assign \mchip.reset  = io_in[13];
	assign \mchip.right  = io_in[1];
	assign \mchip.y [6:4] = 3'h0;
endmodule
module d21_varunk2_motorctrl (
	io_in,
	io_out
);
	wire _000_;
	wire _001_;
	wire _002_;
	wire _003_;
	wire _004_;
	wire _005_;
	wire _006_;
	wire _007_;
	wire _008_;
	wire _009_;
	wire _010_;
	wire _011_;
	wire _012_;
	wire _013_;
	wire _014_;
	wire _015_;
	wire _016_;
	wire _017_;
	wire _018_;
	wire _019_;
	wire _020_;
	wire _021_;
	wire _022_;
	wire _023_;
	wire _024_;
	wire _025_;
	wire _026_;
	wire _027_;
	wire _028_;
	wire _029_;
	wire _030_;
	wire _031_;
	wire _032_;
	wire _033_;
	wire _034_;
	wire _035_;
	wire _036_;
	wire _037_;
	wire _038_;
	wire _039_;
	wire _040_;
	wire _041_;
	wire _042_;
	wire _043_;
	wire _044_;
	wire _045_;
	wire _046_;
	wire _047_;
	wire _048_;
	wire _049_;
	wire _050_;
	wire _051_;
	wire _052_;
	wire _053_;
	wire _054_;
	wire _055_;
	wire _056_;
	wire _057_;
	wire _058_;
	wire _059_;
	wire _060_;
	wire _061_;
	wire _062_;
	wire _063_;
	wire _064_;
	wire _065_;
	wire _066_;
	wire _067_;
	wire _068_;
	wire _069_;
	wire _070_;
	wire _071_;
	wire _072_;
	wire _073_;
	wire _074_;
	wire _075_;
	wire _076_;
	wire _077_;
	wire _078_;
	wire _079_;
	wire _080_;
	wire _081_;
	wire _082_;
	wire _083_;
	wire _084_;
	wire _085_;
	wire _086_;
	wire _087_;
	wire _088_;
	wire _089_;
	wire _090_;
	wire _091_;
	wire _092_;
	wire _093_;
	wire _094_;
	wire _095_;
	wire _096_;
	wire _097_;
	wire _098_;
	wire _099_;
	wire _100_;
	wire _101_;
	wire _102_;
	wire _103_;
	wire _104_;
	wire _105_;
	wire _106_;
	wire _107_;
	wire _108_;
	wire _109_;
	wire _110_;
	wire _111_;
	wire _112_;
	wire _113_;
	wire _114_;
	wire _115_;
	wire _116_;
	wire _117_;
	wire _118_;
	wire _119_;
	wire _120_;
	wire _121_;
	wire _122_;
	wire _123_;
	wire _124_;
	wire _125_;
	wire _126_;
	wire _127_;
	wire _128_;
	wire _129_;
	wire _130_;
	wire _131_;
	wire _132_;
	wire _133_;
	wire _134_;
	wire _135_;
	wire _136_;
	wire _137_;
	wire _138_;
	wire _139_;
	wire _140_;
	wire _141_;
	wire _142_;
	wire _143_;
	wire _144_;
	wire _145_;
	wire _146_;
	wire _147_;
	wire _148_;
	wire _149_;
	wire _150_;
	wire _151_;
	wire _152_;
	wire _153_;
	wire _154_;
	wire _155_;
	wire _156_;
	wire _157_;
	wire _158_;
	wire _159_;
	wire _160_;
	wire _161_;
	wire _162_;
	wire _163_;
	wire _164_;
	wire _165_;
	wire _166_;
	wire _167_;
	wire _168_;
	wire _169_;
	wire _170_;
	wire _171_;
	wire _172_;
	wire _173_;
	wire _174_;
	wire _175_;
	wire _176_;
	wire _177_;
	wire _178_;
	wire _179_;
	wire _180_;
	wire _181_;
	wire _182_;
	wire _183_;
	wire _184_;
	wire _185_;
	wire _186_;
	wire _187_;
	wire _188_;
	wire _189_;
	wire _190_;
	wire _191_;
	wire _192_;
	wire _193_;
	wire _194_;
	wire _195_;
	wire _196_;
	wire _197_;
	wire _198_;
	wire _199_;
	wire _200_;
	wire _201_;
	wire _202_;
	wire _203_;
	wire _204_;
	wire _205_;
	wire _206_;
	wire _207_;
	wire _208_;
	wire _209_;
	wire _210_;
	wire _211_;
	wire _212_;
	wire _213_;
	wire _214_;
	wire _215_;
	wire _216_;
	wire _217_;
	wire _218_;
	wire _219_;
	wire _220_;
	wire _221_;
	wire _222_;
	wire _223_;
	wire _224_;
	wire _225_;
	wire _226_;
	wire _227_;
	wire _228_;
	wire _229_;
	wire _230_;
	wire _231_;
	wire _232_;
	wire _233_;
	wire _234_;
	wire _235_;
	wire _236_;
	wire _237_;
	wire _238_;
	wire _239_;
	wire _240_;
	wire _241_;
	wire _242_;
	wire _243_;
	wire _244_;
	wire _245_;
	wire _246_;
	wire _247_;
	wire _248_;
	wire _249_;
	wire _250_;
	wire _251_;
	wire _252_;
	wire _253_;
	wire _254_;
	wire _255_;
	wire _256_;
	wire _257_;
	wire _258_;
	wire _259_;
	wire _260_;
	wire _261_;
	wire _262_;
	wire _263_;
	wire _264_;
	wire _265_;
	wire _266_;
	wire _267_;
	wire _268_;
	wire _269_;
	wire _270_;
	wire _271_;
	wire _272_;
	wire _273_;
	wire _274_;
	wire _275_;
	wire _276_;
	wire _277_;
	wire _278_;
	wire _279_;
	wire _280_;
	wire _281_;
	wire _282_;
	wire _283_;
	wire _284_;
	wire _285_;
	wire _286_;
	wire _287_;
	wire _288_;
	wire _289_;
	wire _290_;
	wire _291_;
	wire _292_;
	wire _293_;
	wire _294_;
	wire _295_;
	wire _296_;
	wire _297_;
	wire _298_;
	wire _299_;
	wire _300_;
	wire _301_;
	wire _302_;
	wire _303_;
	wire _304_;
	wire _305_;
	wire _306_;
	wire _307_;
	wire _308_;
	wire _309_;
	wire _310_;
	wire _311_;
	wire _312_;
	wire _313_;
	wire _314_;
	wire _315_;
	wire _316_;
	wire _317_;
	wire _318_;
	wire _319_;
	wire _320_;
	wire _321_;
	wire _322_;
	wire _323_;
	wire _324_;
	wire _325_;
	wire _326_;
	wire _327_;
	wire _328_;
	wire _329_;
	wire _330_;
	wire _331_;
	wire _332_;
	wire _333_;
	wire _334_;
	wire _335_;
	wire _336_;
	wire _337_;
	wire _338_;
	wire _339_;
	wire _340_;
	wire _341_;
	wire _342_;
	wire _343_;
	wire _344_;
	wire _345_;
	wire _346_;
	wire _347_;
	wire _348_;
	wire _349_;
	wire _350_;
	wire _351_;
	wire _352_;
	wire _353_;
	wire _354_;
	wire _355_;
	wire _356_;
	wire _357_;
	wire _358_;
	wire _359_;
	wire _360_;
	wire _361_;
	wire _362_;
	wire _363_;
	wire _364_;
	wire _365_;
	wire _366_;
	wire _367_;
	wire _368_;
	wire _369_;
	wire _370_;
	wire _371_;
	wire _372_;
	wire _373_;
	wire _374_;
	wire _375_;
	wire _376_;
	wire _377_;
	wire _378_;
	wire _379_;
	wire _380_;
	wire _381_;
	wire _382_;
	wire _383_;
	wire _384_;
	wire _385_;
	wire _386_;
	wire _387_;
	wire _388_;
	wire _389_;
	wire _390_;
	wire _391_;
	wire _392_;
	wire _393_;
	wire _394_;
	wire _395_;
	wire _396_;
	wire _397_;
	wire _398_;
	wire _399_;
	wire _400_;
	wire _401_;
	wire _402_;
	wire _403_;
	wire _404_;
	wire _405_;
	wire _406_;
	wire _407_;
	wire _408_;
	wire _409_;
	wire _410_;
	wire _411_;
	wire _412_;
	wire _413_;
	wire _414_;
	wire _415_;
	wire [3:0] _416_;
	wire [3:0] _417_;
	wire [19:0] _418_;
	wire [19:0] _419_;
	wire [3:0] _420_;
	wire [3:0] _421_;
	wire [19:0] _422_;
	wire [19:0] _423_;
	input wire [13:0] io_in;
	output wire [13:0] io_out;
	wire \mchip.DECODE_1.A ;
	reg \mchip.DECODE_1.A_prev ;
	wire \mchip.DECODE_1.B ;
	reg \mchip.DECODE_1.B_prev ;
	wire \mchip.DECODE_1.clock ;
	reg \mchip.DECODE_1.dir ;
	reg \mchip.DECODE_1.p ;
	wire \mchip.DECODE_1.reset ;
	wire \mchip.DECODE_2.A ;
	reg \mchip.DECODE_2.A_prev ;
	wire \mchip.DECODE_2.B ;
	reg \mchip.DECODE_2.B_prev ;
	wire \mchip.DECODE_2.clock ;
	reg \mchip.DECODE_2.dir ;
	reg \mchip.DECODE_2.p ;
	wire \mchip.DECODE_2.reset ;
	wire \mchip.PWM_1.CLK ;
	wire \mchip.PWM_1.M_OUT ;
	wire \mchip.PWM_1.PWM_DUTY ;
	wire \mchip.PWM_1.PWM_PERIOD ;
	wire \mchip.PWM_1.SCL ;
	wire \mchip.PWM_1.reset ;
	wire \mchip.PWM_2.CLK ;
	wire \mchip.PWM_2.M_OUT ;
	wire \mchip.PWM_2.PWM_DUTY ;
	wire \mchip.PWM_2.PWM_PERIOD ;
	wire \mchip.PWM_2.SCL ;
	wire \mchip.PWM_2.reset ;
	wire \mchip.SERVO_1.CLK ;
	wire \mchip.SERVO_1.SCL ;
	wire \mchip.SERVO_1.S_IN ;
	wire \mchip.SERVO_1.S_OUT ;
	reg [3:0] \mchip.SERVO_1.eight_count ;
	reg \mchip.SERVO_1.last_in_clk ;
	reg [7:0] \mchip.SERVO_1.position ;
	wire \mchip.SERVO_1.pwm.clk ;
	reg [19:0] \mchip.SERVO_1.pwm.ctr_d ;
	wire [7:0] \mchip.SERVO_1.pwm.position ;
	wire \mchip.SERVO_1.pwm.rst ;
	reg \mchip.SERVO_1.pwm.servo ;
	wire [19:0] \mchip.SERVO_1.pwm.temp_val ;
	wire \mchip.SERVO_1.reset ;
	reg [7:0] \mchip.SERVO_1.shreg ;
	wire \mchip.SERVO_2.CLK ;
	wire \mchip.SERVO_2.SCL ;
	wire \mchip.SERVO_2.S_IN ;
	wire \mchip.SERVO_2.S_OUT ;
	reg [3:0] \mchip.SERVO_2.eight_count ;
	wire \mchip.SERVO_2.last_in_clk ;
	reg [7:0] \mchip.SERVO_2.position ;
	wire \mchip.SERVO_2.pwm.clk ;
	reg [19:0] \mchip.SERVO_2.pwm.ctr_d ;
	wire [7:0] \mchip.SERVO_2.pwm.position ;
	wire \mchip.SERVO_2.pwm.rst ;
	reg \mchip.SERVO_2.pwm.servo ;
	wire [19:0] \mchip.SERVO_2.pwm.temp_val ;
	wire \mchip.SERVO_2.reset ;
	reg [7:0] \mchip.SERVO_2.shreg ;
	wire \mchip.clock ;
	wire [11:0] \mchip.io_in ;
	wire [11:0] \mchip.io_out ;
	wire \mchip.reset ;
	assign _013_ = ~(\mchip.SERVO_2.eight_count [0] | \mchip.SERVO_2.eight_count [1]);
	assign _014_ = \mchip.SERVO_2.eight_count [2] | ~\mchip.SERVO_2.eight_count [3];
	assign _015_ = _013_ & ~_014_;
	assign _005_ = _015_ | io_in[13];
	assign _016_ = io_in[6] & ~\mchip.DECODE_1.A_prev ;
	assign _007_ = _016_ & ~io_in[7];
	assign _017_ = io_in[7] & ~\mchip.DECODE_1.B_prev ;
	assign _018_ = _017_ & ~io_in[6];
	assign _001_ = _018_ | _007_;
	assign _019_ = io_in[8] & ~\mchip.DECODE_2.A_prev ;
	assign _009_ = _019_ & ~io_in[9];
	assign _020_ = io_in[9] & ~\mchip.DECODE_2.B_prev ;
	assign _021_ = _020_ & ~io_in[8];
	assign _000_ = _021_ | _009_;
	assign _022_ = ~(\mchip.SERVO_1.eight_count [0] | \mchip.SERVO_1.eight_count [1]);
	assign _023_ = \mchip.SERVO_1.eight_count [2] | ~\mchip.SERVO_1.eight_count [3];
	assign _024_ = _022_ & ~_023_;
	assign _004_ = _024_ & ~io_in[13];
	assign _006_ = _024_ | io_in[13];
	assign _025_ = io_in[11] & ~\mchip.SERVO_1.last_in_clk ;
	assign _003_ = _025_ & ~io_in[13];
	assign _002_ = _015_ & ~io_in[13];
	assign _026_ = ~(\mchip.SERVO_2.pwm.ctr_d [0] | \mchip.SERVO_2.pwm.ctr_d [1]);
	assign _027_ = \mchip.SERVO_2.pwm.ctr_d [2] | \mchip.SERVO_2.pwm.ctr_d [3];
	assign _028_ = _026_ & ~_027_;
	assign _029_ = \mchip.SERVO_2.pwm.ctr_d [6] | \mchip.SERVO_2.pwm.ctr_d [7];
	assign _030_ = \mchip.SERVO_2.pwm.ctr_d [4] | ~\mchip.SERVO_2.pwm.ctr_d [5];
	assign _031_ = _030_ | _029_;
	assign _032_ = _028_ & ~_031_;
	assign _033_ = \mchip.SERVO_2.pwm.ctr_d [15] | ~\mchip.SERVO_2.pwm.ctr_d [14];
	assign _034_ = \mchip.SERVO_2.pwm.ctr_d [12] | \mchip.SERVO_2.pwm.ctr_d [13];
	assign _035_ = _034_ | _033_;
	assign _036_ = ~(\mchip.SERVO_2.pwm.ctr_d [10] & \mchip.SERVO_2.pwm.ctr_d [11]);
	assign _037_ = \mchip.SERVO_2.pwm.ctr_d [8] | ~\mchip.SERVO_2.pwm.ctr_d [9];
	assign _038_ = _037_ | _036_;
	assign _039_ = _038_ | _035_;
	assign _040_ = _032_ & ~_039_;
	assign _041_ = \mchip.SERVO_2.pwm.ctr_d [18] | \mchip.SERVO_2.pwm.ctr_d [19];
	assign _042_ = \mchip.SERVO_2.pwm.ctr_d [16] | \mchip.SERVO_2.pwm.ctr_d [17];
	assign _043_ = _042_ | _041_;
	assign _044_ = _040_ & ~_043_;
	assign _045_ = \mchip.SERVO_2.pwm.ctr_d [0] & ~_044_;
	assign _422_[0] = ~_045_;
	assign _416_[0] = ~\mchip.SERVO_1.eight_count [0];
	assign _046_ = ~\mchip.SERVO_2.position [7];
	assign _047_ = ~(\mchip.SERVO_2.position [5] | \mchip.SERVO_2.position [6]);
	assign _048_ = ~(\mchip.SERVO_2.position [3] | \mchip.SERVO_2.position [4]);
	assign _049_ = \mchip.SERVO_2.position [1] & \mchip.SERVO_2.position [2];
	assign _050_ = _049_ | ~_048_;
	assign _051_ = _047_ & ~_050_;
	assign _052_ = _051_ ^ _046_;
	assign _053_ = _048_ & ~_049_;
	assign _054_ = _053_ & ~\mchip.SERVO_2.position [5];
	assign _055_ = _054_ ^ \mchip.SERVO_2.position [6];
	assign _056_ = _052_ & ~_055_;
	assign _057_ = _053_ ^ \mchip.SERVO_2.position [5];
	assign _058_ = ~(_049_ | \mchip.SERVO_2.position [3]);
	assign _059_ = _058_ ^ \mchip.SERVO_2.position [4];
	assign _060_ = _059_ | _057_;
	assign _061_ = _056_ & ~_060_;
	assign _062_ = _049_ ^ \mchip.SERVO_2.position [3];
	assign _063_ = \mchip.SERVO_2.position [1] ^ \mchip.SERVO_2.position [2];
	assign _064_ = _062_ & ~_063_;
	assign _065_ = \mchip.SERVO_2.position [0] & ~\mchip.SERVO_2.position [1];
	assign _066_ = _064_ & ~_065_;
	assign _067_ = _061_ & ~_066_;
	assign _068_ = _067_ | ~_061_;
	assign _069_ = _051_ & ~\mchip.SERVO_2.position [7];
	assign _070_ = ~_069_;
	assign _071_ = _070_ | _068_;
	assign _072_ = \mchip.SERVO_2.pwm.ctr_d [19] & ~_044_;
	assign _073_ = ~(_072_ & _071_);
	assign _074_ = _072_ ^ _071_;
	assign _075_ = \mchip.SERVO_2.pwm.ctr_d [18] & ~_044_;
	assign _076_ = ~(_075_ & _071_);
	assign _077_ = _074_ & ~_076_;
	assign _078_ = _073_ & ~_077_;
	assign _079_ = _069_ & ~_068_;
	assign _080_ = _075_ ^ _079_;
	assign _081_ = _074_ & ~_080_;
	assign _082_ = \mchip.SERVO_2.pwm.ctr_d [17] & ~_044_;
	assign _083_ = ~(_082_ & _071_);
	assign _084_ = _082_ ^ _071_;
	assign _085_ = \mchip.SERVO_2.pwm.ctr_d [16] & ~_044_;
	assign _086_ = ~(_085_ & _071_);
	assign _087_ = _084_ & ~_086_;
	assign _088_ = _083_ & ~_087_;
	assign _089_ = _085_ ^ _079_;
	assign _090_ = _084_ & ~_089_;
	assign _091_ = \mchip.SERVO_2.pwm.ctr_d [15] & ~_044_;
	assign _092_ = ~(_091_ & _071_);
	assign _093_ = _044_ | ~\mchip.SERVO_2.pwm.ctr_d [14];
	assign _094_ = _071_ & ~_093_;
	assign _095_ = _091_ ^ _079_;
	assign _096_ = _094_ & ~_095_;
	assign _097_ = _092_ & ~_096_;
	assign _098_ = _090_ & ~_097_;
	assign _099_ = _088_ & ~_098_;
	assign _100_ = ~_093_;
	assign _101_ = _100_ ^ _079_;
	assign _102_ = _101_ | _095_;
	assign _103_ = _090_ & ~_102_;
	assign _104_ = \mchip.SERVO_2.pwm.ctr_d [13] & ~_044_;
	assign _105_ = ~(_104_ & _071_);
	assign _106_ = _104_ ^ _079_;
	assign _107_ = \mchip.SERVO_2.pwm.ctr_d [12] & ~_044_;
	assign _108_ = ~_107_;
	assign _109_ = _071_ & ~_108_;
	assign _110_ = _109_ & ~_106_;
	assign _111_ = _105_ & ~_110_;
	assign _112_ = \mchip.SERVO_2.pwm.ctr_d [11] & ~_044_;
	assign _113_ = ~_112_;
	assign _114_ = _071_ & ~_113_;
	assign _115_ = _069_ ^ _068_;
	assign _116_ = _044_ | ~\mchip.SERVO_2.pwm.ctr_d [10];
	assign _117_ = ~_116_;
	assign _118_ = _117_ & ~_115_;
	assign _119_ = _112_ ^ _079_;
	assign _120_ = _118_ & ~_119_;
	assign _121_ = _120_ | _114_;
	assign _122_ = _107_ ^ _079_;
	assign _123_ = _122_ | _106_;
	assign _124_ = _121_ & ~_123_;
	assign _125_ = _111_ & ~_124_;
	assign _126_ = _103_ & ~_125_;
	assign _127_ = _099_ & ~_126_;
	assign _128_ = _117_ ^ _115_;
	assign _129_ = _128_ | _119_;
	assign _130_ = _129_ | _123_;
	assign _131_ = _103_ & ~_130_;
	assign _132_ = _066_ & ~_060_;
	assign _133_ = _132_ & ~_055_;
	assign _134_ = _133_ ^ _052_;
	assign _135_ = \mchip.SERVO_2.pwm.ctr_d [9] & ~_044_;
	assign _136_ = ~(_135_ & _134_);
	assign _137_ = _135_ ^ _134_;
	assign _138_ = \mchip.SERVO_2.pwm.ctr_d [8] & ~_044_;
	assign _139_ = _132_ ^ _055_;
	assign _140_ = _139_ | ~_138_;
	assign _141_ = _137_ & ~_140_;
	assign _142_ = _136_ & ~_141_;
	assign _143_ = _139_ ^ _138_;
	assign _144_ = _137_ & ~_143_;
	assign _145_ = _066_ & ~_059_;
	assign _146_ = _145_ ^ _057_;
	assign _147_ = \mchip.SERVO_2.pwm.ctr_d [7] & ~_044_;
	assign _148_ = _146_ | ~_147_;
	assign _149_ = _147_ ^ _146_;
	assign _150_ = _066_ ^ _059_;
	assign _151_ = \mchip.SERVO_2.pwm.ctr_d [6] & ~_044_;
	assign _152_ = _151_ & ~_150_;
	assign _153_ = _152_ & ~_149_;
	assign _154_ = _148_ & ~_153_;
	assign _155_ = _144_ & ~_154_;
	assign _156_ = _142_ & ~_155_;
	assign _157_ = _151_ ^ _150_;
	assign _158_ = _157_ | _149_;
	assign _159_ = _144_ & ~_158_;
	assign _160_ = ~(_065_ | _063_);
	assign _161_ = ~(_160_ ^ _062_);
	assign _162_ = _044_ | ~\mchip.SERVO_2.pwm.ctr_d [5];
	assign _163_ = _162_ | _161_;
	assign _164_ = _162_ ^ _161_;
	assign _165_ = ~(_065_ ^ _063_);
	assign _166_ = \mchip.SERVO_2.pwm.ctr_d [4] & ~_044_;
	assign _167_ = _165_ | ~_166_;
	assign _168_ = _164_ & ~_167_;
	assign _169_ = _163_ & ~_168_;
	assign _170_ = _166_ ^ _165_;
	assign _171_ = _164_ & ~_170_;
	assign _172_ = ~(\mchip.SERVO_2.position [0] ^ \mchip.SERVO_2.position [1]);
	assign _173_ = _044_ | ~\mchip.SERVO_2.pwm.ctr_d [3];
	assign _174_ = _173_ | _172_;
	assign _175_ = _173_ ^ _172_;
	assign _176_ = \mchip.SERVO_2.pwm.ctr_d [2] & ~_044_;
	assign _177_ = ~(_176_ | \mchip.SERVO_2.position [0]);
	assign _178_ = _175_ & ~_177_;
	assign _179_ = _174_ & ~_178_;
	assign _180_ = _171_ & ~_179_;
	assign _181_ = _169_ & ~_180_;
	assign _182_ = _159_ & ~_181_;
	assign _183_ = _156_ & ~_182_;
	assign _184_ = _131_ & ~_183_;
	assign _185_ = _127_ & ~_184_;
	assign _186_ = _081_ & ~_185_;
	assign _012_ = _078_ & ~_186_;
	assign _187_ = ~\mchip.SERVO_1.position [7];
	assign _188_ = ~(\mchip.SERVO_1.position [6] | \mchip.SERVO_1.position [5]);
	assign _189_ = ~(\mchip.SERVO_1.position [3] | \mchip.SERVO_1.position [4]);
	assign _190_ = \mchip.SERVO_1.position [1] & \mchip.SERVO_1.position [2];
	assign _191_ = _190_ | ~_189_;
	assign _192_ = _188_ & ~_191_;
	assign _193_ = _192_ ^ _187_;
	assign _194_ = _189_ & ~_190_;
	assign _195_ = _194_ & ~\mchip.SERVO_1.position [5];
	assign _196_ = _195_ ^ \mchip.SERVO_1.position [6];
	assign _197_ = _193_ & ~_196_;
	assign _198_ = _194_ ^ \mchip.SERVO_1.position [5];
	assign _199_ = ~(_190_ | \mchip.SERVO_1.position [3]);
	assign _200_ = _199_ ^ \mchip.SERVO_1.position [4];
	assign _201_ = _200_ | _198_;
	assign _202_ = _197_ & ~_201_;
	assign _203_ = _190_ ^ \mchip.SERVO_1.position [3];
	assign _204_ = \mchip.SERVO_1.position [1] ^ \mchip.SERVO_1.position [2];
	assign _205_ = _203_ & ~_204_;
	assign _206_ = \mchip.SERVO_1.position [0] & ~\mchip.SERVO_1.position [1];
	assign _207_ = _205_ & ~_206_;
	assign _208_ = _202_ & ~_207_;
	assign _209_ = _208_ | ~_202_;
	assign _210_ = _192_ & ~\mchip.SERVO_1.position [7];
	assign _211_ = ~_210_;
	assign _212_ = _211_ | _209_;
	assign _213_ = ~(\mchip.SERVO_1.pwm.ctr_d [0] | \mchip.SERVO_1.pwm.ctr_d [1]);
	assign _214_ = \mchip.SERVO_1.pwm.ctr_d [2] | \mchip.SERVO_1.pwm.ctr_d [3];
	assign _215_ = _213_ & ~_214_;
	assign _216_ = \mchip.SERVO_1.pwm.ctr_d [6] | \mchip.SERVO_1.pwm.ctr_d [7];
	assign _217_ = \mchip.SERVO_1.pwm.ctr_d [4] | ~\mchip.SERVO_1.pwm.ctr_d [5];
	assign _218_ = _217_ | _216_;
	assign _219_ = _215_ & ~_218_;
	assign _220_ = \mchip.SERVO_1.pwm.ctr_d [15] | ~\mchip.SERVO_1.pwm.ctr_d [14];
	assign _221_ = \mchip.SERVO_1.pwm.ctr_d [12] | \mchip.SERVO_1.pwm.ctr_d [13];
	assign _222_ = _221_ | _220_;
	assign _223_ = ~(\mchip.SERVO_1.pwm.ctr_d [10] & \mchip.SERVO_1.pwm.ctr_d [11]);
	assign _224_ = \mchip.SERVO_1.pwm.ctr_d [8] | ~\mchip.SERVO_1.pwm.ctr_d [9];
	assign _225_ = _224_ | _223_;
	assign _226_ = _225_ | _222_;
	assign _227_ = _219_ & ~_226_;
	assign _228_ = \mchip.SERVO_1.pwm.ctr_d [18] | \mchip.SERVO_1.pwm.ctr_d [19];
	assign _229_ = \mchip.SERVO_1.pwm.ctr_d [16] | \mchip.SERVO_1.pwm.ctr_d [17];
	assign _230_ = _229_ | _228_;
	assign _231_ = _227_ & ~_230_;
	assign _232_ = \mchip.SERVO_1.pwm.ctr_d [19] & ~_231_;
	assign _233_ = ~(_232_ & _212_);
	assign _234_ = _232_ ^ _212_;
	assign _235_ = \mchip.SERVO_1.pwm.ctr_d [18] & ~_231_;
	assign _236_ = ~(_235_ & _212_);
	assign _237_ = _234_ & ~_236_;
	assign _238_ = _233_ & ~_237_;
	assign _239_ = _210_ & ~_209_;
	assign _240_ = _235_ ^ _239_;
	assign _241_ = _234_ & ~_240_;
	assign _242_ = \mchip.SERVO_1.pwm.ctr_d [17] & ~_231_;
	assign _243_ = ~(_242_ & _212_);
	assign _244_ = _242_ ^ _212_;
	assign _245_ = \mchip.SERVO_1.pwm.ctr_d [16] & ~_231_;
	assign _246_ = ~(_245_ & _212_);
	assign _247_ = _244_ & ~_246_;
	assign _248_ = _243_ & ~_247_;
	assign _249_ = _245_ ^ _239_;
	assign _250_ = _244_ & ~_249_;
	assign _251_ = \mchip.SERVO_1.pwm.ctr_d [15] & ~_231_;
	assign _252_ = ~(_251_ & _212_);
	assign _253_ = _231_ | ~\mchip.SERVO_1.pwm.ctr_d [14];
	assign _254_ = _212_ & ~_253_;
	assign _255_ = _251_ ^ _239_;
	assign _256_ = _254_ & ~_255_;
	assign _257_ = _252_ & ~_256_;
	assign _258_ = _250_ & ~_257_;
	assign _259_ = _248_ & ~_258_;
	assign _260_ = ~_253_;
	assign _261_ = _260_ ^ _239_;
	assign _262_ = _261_ | _255_;
	assign _263_ = _250_ & ~_262_;
	assign _264_ = \mchip.SERVO_1.pwm.ctr_d [13] & ~_231_;
	assign _265_ = ~(_264_ & _212_);
	assign _266_ = _264_ ^ _239_;
	assign _267_ = \mchip.SERVO_1.pwm.ctr_d [12] & ~_231_;
	assign _268_ = ~_267_;
	assign _269_ = _212_ & ~_268_;
	assign _270_ = _269_ & ~_266_;
	assign _271_ = _265_ & ~_270_;
	assign _272_ = \mchip.SERVO_1.pwm.ctr_d [11] & ~_231_;
	assign _273_ = ~_272_;
	assign _274_ = _212_ & ~_273_;
	assign _275_ = _210_ ^ _209_;
	assign _276_ = _231_ | ~\mchip.SERVO_1.pwm.ctr_d [10];
	assign _277_ = ~_276_;
	assign _278_ = _277_ & ~_275_;
	assign _279_ = _272_ ^ _239_;
	assign _280_ = _278_ & ~_279_;
	assign _281_ = _280_ | _274_;
	assign _282_ = _267_ ^ _239_;
	assign _283_ = _282_ | _266_;
	assign _284_ = _281_ & ~_283_;
	assign _285_ = _271_ & ~_284_;
	assign _286_ = _263_ & ~_285_;
	assign _287_ = _259_ & ~_286_;
	assign _288_ = _277_ ^ _275_;
	assign _289_ = _288_ | _279_;
	assign _290_ = _289_ | _283_;
	assign _291_ = _263_ & ~_290_;
	assign _292_ = _207_ & ~_201_;
	assign _293_ = _292_ & ~_196_;
	assign _294_ = _293_ ^ _193_;
	assign _295_ = \mchip.SERVO_1.pwm.ctr_d [9] & ~_231_;
	assign _296_ = ~(_295_ & _294_);
	assign _297_ = _295_ ^ _294_;
	assign _298_ = \mchip.SERVO_1.pwm.ctr_d [8] & ~_231_;
	assign _299_ = _292_ ^ _196_;
	assign _300_ = _299_ | ~_298_;
	assign _301_ = _297_ & ~_300_;
	assign _302_ = _296_ & ~_301_;
	assign _303_ = _299_ ^ _298_;
	assign _304_ = _297_ & ~_303_;
	assign _305_ = _207_ & ~_200_;
	assign _306_ = _305_ ^ _198_;
	assign _307_ = \mchip.SERVO_1.pwm.ctr_d [7] & ~_231_;
	assign _308_ = _306_ | ~_307_;
	assign _309_ = _307_ ^ _306_;
	assign _310_ = _207_ ^ _200_;
	assign _311_ = \mchip.SERVO_1.pwm.ctr_d [6] & ~_231_;
	assign _312_ = _311_ & ~_310_;
	assign _313_ = _312_ & ~_309_;
	assign _314_ = _308_ & ~_313_;
	assign _315_ = _304_ & ~_314_;
	assign _316_ = _302_ & ~_315_;
	assign _317_ = _311_ ^ _310_;
	assign _318_ = _317_ | _309_;
	assign _319_ = _304_ & ~_318_;
	assign _320_ = ~(_206_ | _204_);
	assign _321_ = ~(_320_ ^ _203_);
	assign _322_ = _231_ | ~\mchip.SERVO_1.pwm.ctr_d [5];
	assign _323_ = _322_ | _321_;
	assign _324_ = _322_ ^ _321_;
	assign _325_ = ~(_206_ ^ _204_);
	assign _326_ = \mchip.SERVO_1.pwm.ctr_d [4] & ~_231_;
	assign _327_ = _325_ | ~_326_;
	assign _328_ = _324_ & ~_327_;
	assign _329_ = _323_ & ~_328_;
	assign _330_ = _326_ ^ _325_;
	assign _331_ = _324_ & ~_330_;
	assign _332_ = ~(\mchip.SERVO_1.position [0] ^ \mchip.SERVO_1.position [1]);
	assign _333_ = _231_ | ~\mchip.SERVO_1.pwm.ctr_d [3];
	assign _334_ = _333_ | _332_;
	assign _335_ = _333_ ^ _332_;
	assign _336_ = \mchip.SERVO_1.pwm.ctr_d [2] & ~_231_;
	assign _337_ = ~(_336_ | \mchip.SERVO_1.position [0]);
	assign _338_ = _335_ & ~_337_;
	assign _339_ = _334_ & ~_338_;
	assign _340_ = _331_ & ~_339_;
	assign _341_ = _329_ & ~_340_;
	assign _342_ = _319_ & ~_341_;
	assign _343_ = _316_ & ~_342_;
	assign _344_ = _291_ & ~_343_;
	assign _345_ = _287_ & ~_344_;
	assign _346_ = _241_ & ~_345_;
	assign _011_ = _238_ & ~_346_;
	assign _347_ = \mchip.SERVO_1.pwm.ctr_d [0] & ~_231_;
	assign _418_[0] = ~_347_;
	assign _420_[0] = ~\mchip.SERVO_2.eight_count [0];
	assign _348_ = _044_ | ~\mchip.SERVO_2.pwm.ctr_d [1];
	assign _423_[1] = ~(_348_ ^ _045_);
	assign _349_ = _045_ & ~_348_;
	assign _423_[2] = _349_ ^ _176_;
	assign _350_ = ~(_349_ & _176_);
	assign _423_[3] = _350_ ^ _173_;
	assign _351_ = _173_ | ~_176_;
	assign _352_ = _349_ & ~_351_;
	assign _423_[4] = _352_ ^ _166_;
	assign _353_ = ~(_352_ & _166_);
	assign _423_[5] = _353_ ^ _162_;
	assign _354_ = _162_ | ~_166_;
	assign _355_ = _352_ & ~_354_;
	assign _423_[6] = _355_ ^ _151_;
	assign _356_ = ~_151_;
	assign _357_ = _355_ & ~_356_;
	assign _423_[7] = _357_ ^ _147_;
	assign _358_ = ~(_151_ & _147_);
	assign _359_ = _358_ | _354_;
	assign _360_ = _352_ & ~_359_;
	assign _423_[8] = _360_ ^ _138_;
	assign _361_ = _360_ & _138_;
	assign _423_[9] = _361_ ^ _135_;
	assign _362_ = ~(_138_ & _135_);
	assign _363_ = _360_ & ~_362_;
	assign _423_[10] = _363_ ^ _117_;
	assign _364_ = _363_ & ~_116_;
	assign _423_[11] = _364_ ^ _112_;
	assign _365_ = _116_ | ~_112_;
	assign _366_ = _365_ | _362_;
	assign _367_ = _360_ & ~_366_;
	assign _423_[12] = _367_ ^ _107_;
	assign _368_ = _367_ & ~_108_;
	assign _423_[13] = _368_ ^ _104_;
	assign _369_ = ~(_107_ & _104_);
	assign _370_ = _367_ & ~_369_;
	assign _423_[14] = _370_ ^ _100_;
	assign _371_ = _370_ & ~_093_;
	assign _423_[15] = _371_ ^ _091_;
	assign _372_ = _093_ | ~_091_;
	assign _373_ = _372_ | _369_;
	assign _374_ = _373_ | _366_;
	assign _375_ = _360_ & ~_374_;
	assign _423_[16] = _375_ ^ _085_;
	assign _376_ = _375_ & _085_;
	assign _423_[17] = _376_ ^ _082_;
	assign _377_ = ~(\mchip.SERVO_2.pwm.ctr_d [16] & \mchip.SERVO_2.pwm.ctr_d [17]);
	assign _378_ = _375_ & ~_377_;
	assign _423_[18] = _378_ ^ _075_;
	assign _379_ = _378_ & _075_;
	assign _423_[19] = _379_ ^ _072_;
	assign _417_[1] = \mchip.SERVO_1.eight_count [0] ^ \mchip.SERVO_1.eight_count [1];
	assign _380_ = \mchip.SERVO_1.eight_count [0] & \mchip.SERVO_1.eight_count [1];
	assign _417_[2] = _380_ ^ \mchip.SERVO_1.eight_count [2];
	assign _381_ = _380_ & \mchip.SERVO_1.eight_count [2];
	assign _417_[3] = _381_ ^ \mchip.SERVO_1.eight_count [3];
	assign _010_ = io_in[8] & ~io_in[9];
	assign _008_ = io_in[6] & ~io_in[7];
	assign _421_[1] = \mchip.SERVO_2.eight_count [0] ^ \mchip.SERVO_2.eight_count [1];
	assign _382_ = \mchip.SERVO_2.eight_count [0] & \mchip.SERVO_2.eight_count [1];
	assign _421_[2] = _382_ ^ \mchip.SERVO_2.eight_count [2];
	assign _383_ = _382_ & \mchip.SERVO_2.eight_count [2];
	assign _421_[3] = _383_ ^ \mchip.SERVO_2.eight_count [3];
	assign _384_ = _231_ | ~\mchip.SERVO_1.pwm.ctr_d [1];
	assign _419_[1] = ~(_384_ ^ _347_);
	assign _385_ = _347_ & ~_384_;
	assign _419_[2] = _385_ ^ _336_;
	assign _386_ = ~(_385_ & _336_);
	assign _419_[3] = _386_ ^ _333_;
	assign _387_ = _333_ | ~_336_;
	assign _388_ = _385_ & ~_387_;
	assign _419_[4] = _388_ ^ _326_;
	assign _389_ = ~(_388_ & _326_);
	assign _419_[5] = _389_ ^ _322_;
	assign _390_ = _322_ | ~_326_;
	assign _391_ = _388_ & ~_390_;
	assign _419_[6] = _391_ ^ _311_;
	assign _392_ = ~_311_;
	assign _393_ = _391_ & ~_392_;
	assign _419_[7] = _393_ ^ _307_;
	assign _394_ = ~(_311_ & _307_);
	assign _395_ = _394_ | _390_;
	assign _396_ = _388_ & ~_395_;
	assign _419_[8] = _396_ ^ _298_;
	assign _397_ = _396_ & _298_;
	assign _419_[9] = _397_ ^ _295_;
	assign _398_ = ~(_298_ & _295_);
	assign _399_ = _396_ & ~_398_;
	assign _419_[10] = _399_ ^ _277_;
	assign _400_ = _399_ & ~_276_;
	assign _419_[11] = _400_ ^ _272_;
	assign _401_ = _276_ | ~_272_;
	assign _402_ = _401_ | _398_;
	assign _403_ = _396_ & ~_402_;
	assign _419_[12] = _403_ ^ _267_;
	assign _404_ = _403_ & ~_268_;
	assign _419_[13] = _404_ ^ _264_;
	assign _405_ = ~(_267_ & _264_);
	assign _406_ = _403_ & ~_405_;
	assign _419_[14] = _406_ ^ _260_;
	assign _407_ = _406_ & ~_253_;
	assign _419_[15] = _407_ ^ _251_;
	assign _408_ = _253_ | ~_251_;
	assign _409_ = _408_ | _405_;
	assign _410_ = _409_ | _402_;
	assign _411_ = _396_ & ~_410_;
	assign _419_[16] = _411_ ^ _245_;
	assign _412_ = _411_ & _245_;
	assign _419_[17] = _412_ ^ _242_;
	assign _413_ = ~(\mchip.SERVO_1.pwm.ctr_d [16] & \mchip.SERVO_1.pwm.ctr_d [17]);
	assign _414_ = _411_ & ~_413_;
	assign _419_[18] = _414_ ^ _235_;
	assign _415_ = _414_ & _235_;
	assign _419_[19] = _415_ ^ _232_;
	always @(posedge io_in[12])
		if (!io_in[13])
			\mchip.SERVO_2.pwm.servo  <= _012_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DECODE_1.p  <= 1'h0;
		else
			\mchip.DECODE_1.p  <= _008_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DECODE_2.dir  <= 1'h0;
		else if (_000_)
			\mchip.DECODE_2.dir  <= _009_;
	always @(posedge io_in[12]) \mchip.DECODE_2.A_prev  <= io_in[8];
	always @(posedge io_in[12]) \mchip.DECODE_2.B_prev  <= io_in[9];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DECODE_1.dir  <= 1'h0;
		else if (_001_)
			\mchip.DECODE_1.dir  <= _007_;
	always @(posedge io_in[12]) \mchip.DECODE_1.A_prev  <= io_in[6];
	always @(posedge io_in[12]) \mchip.DECODE_1.B_prev  <= io_in[7];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.SERVO_2.pwm.ctr_d [0] <= 1'h0;
		else
			\mchip.SERVO_2.pwm.ctr_d [0] <= _422_[0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.SERVO_2.pwm.ctr_d [1] <= 1'h0;
		else
			\mchip.SERVO_2.pwm.ctr_d [1] <= _423_[1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.SERVO_2.pwm.ctr_d [2] <= 1'h0;
		else
			\mchip.SERVO_2.pwm.ctr_d [2] <= _423_[2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.SERVO_2.pwm.ctr_d [3] <= 1'h0;
		else
			\mchip.SERVO_2.pwm.ctr_d [3] <= _423_[3];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.SERVO_2.pwm.ctr_d [4] <= 1'h0;
		else
			\mchip.SERVO_2.pwm.ctr_d [4] <= _423_[4];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.SERVO_2.pwm.ctr_d [5] <= 1'h0;
		else
			\mchip.SERVO_2.pwm.ctr_d [5] <= _423_[5];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.SERVO_2.pwm.ctr_d [6] <= 1'h0;
		else
			\mchip.SERVO_2.pwm.ctr_d [6] <= _423_[6];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.SERVO_2.pwm.ctr_d [7] <= 1'h0;
		else
			\mchip.SERVO_2.pwm.ctr_d [7] <= _423_[7];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.SERVO_2.pwm.ctr_d [8] <= 1'h0;
		else
			\mchip.SERVO_2.pwm.ctr_d [8] <= _423_[8];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.SERVO_2.pwm.ctr_d [9] <= 1'h0;
		else
			\mchip.SERVO_2.pwm.ctr_d [9] <= _423_[9];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.SERVO_2.pwm.ctr_d [10] <= 1'h0;
		else
			\mchip.SERVO_2.pwm.ctr_d [10] <= _423_[10];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.SERVO_2.pwm.ctr_d [11] <= 1'h0;
		else
			\mchip.SERVO_2.pwm.ctr_d [11] <= _423_[11];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.SERVO_2.pwm.ctr_d [12] <= 1'h0;
		else
			\mchip.SERVO_2.pwm.ctr_d [12] <= _423_[12];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.SERVO_2.pwm.ctr_d [13] <= 1'h0;
		else
			\mchip.SERVO_2.pwm.ctr_d [13] <= _423_[13];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.SERVO_2.pwm.ctr_d [14] <= 1'h0;
		else
			\mchip.SERVO_2.pwm.ctr_d [14] <= _423_[14];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.SERVO_2.pwm.ctr_d [15] <= 1'h0;
		else
			\mchip.SERVO_2.pwm.ctr_d [15] <= _423_[15];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.SERVO_2.pwm.ctr_d [16] <= 1'h0;
		else
			\mchip.SERVO_2.pwm.ctr_d [16] <= _423_[16];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.SERVO_2.pwm.ctr_d [17] <= 1'h0;
		else
			\mchip.SERVO_2.pwm.ctr_d [17] <= _423_[17];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.SERVO_2.pwm.ctr_d [18] <= 1'h0;
		else
			\mchip.SERVO_2.pwm.ctr_d [18] <= _423_[18];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.SERVO_2.pwm.ctr_d [19] <= 1'h0;
		else
			\mchip.SERVO_2.pwm.ctr_d [19] <= _423_[19];
	always @(posedge io_in[12])
		if (!io_in[13])
			\mchip.SERVO_1.pwm.servo  <= _011_;
	always @(posedge io_in[12])
		if (_003_)
			\mchip.SERVO_2.shreg [0] <= io_in[5];
	always @(posedge io_in[12])
		if (_003_)
			\mchip.SERVO_2.shreg [1] <= \mchip.SERVO_2.shreg [0];
	always @(posedge io_in[12])
		if (_003_)
			\mchip.SERVO_2.shreg [2] <= \mchip.SERVO_2.shreg [1];
	always @(posedge io_in[12])
		if (_003_)
			\mchip.SERVO_2.shreg [3] <= \mchip.SERVO_2.shreg [2];
	always @(posedge io_in[12])
		if (_003_)
			\mchip.SERVO_2.shreg [4] <= \mchip.SERVO_2.shreg [3];
	always @(posedge io_in[12])
		if (_003_)
			\mchip.SERVO_2.shreg [5] <= \mchip.SERVO_2.shreg [4];
	always @(posedge io_in[12])
		if (_003_)
			\mchip.SERVO_2.shreg [6] <= \mchip.SERVO_2.shreg [5];
	always @(posedge io_in[12])
		if (_003_)
			\mchip.SERVO_2.shreg [7] <= \mchip.SERVO_2.shreg [6];
	always @(posedge io_in[12])
		if (_002_)
			\mchip.SERVO_2.position [0] <= \mchip.SERVO_2.shreg [0];
	always @(posedge io_in[12])
		if (_002_)
			\mchip.SERVO_2.position [1] <= \mchip.SERVO_2.shreg [1];
	always @(posedge io_in[12])
		if (_002_)
			\mchip.SERVO_2.position [2] <= \mchip.SERVO_2.shreg [2];
	always @(posedge io_in[12])
		if (_002_)
			\mchip.SERVO_2.position [3] <= \mchip.SERVO_2.shreg [3];
	always @(posedge io_in[12])
		if (_002_)
			\mchip.SERVO_2.position [4] <= \mchip.SERVO_2.shreg [4];
	always @(posedge io_in[12])
		if (_002_)
			\mchip.SERVO_2.position [5] <= \mchip.SERVO_2.shreg [5];
	always @(posedge io_in[12])
		if (_002_)
			\mchip.SERVO_2.position [6] <= \mchip.SERVO_2.shreg [6];
	always @(posedge io_in[12])
		if (_002_)
			\mchip.SERVO_2.position [7] <= \mchip.SERVO_2.shreg [7];
	always @(posedge io_in[12])
		if (_005_)
			\mchip.SERVO_2.eight_count [0] <= 1'h0;
		else
			\mchip.SERVO_2.eight_count [0] <= _420_[0];
	always @(posedge io_in[12])
		if (_005_)
			\mchip.SERVO_2.eight_count [1] <= 1'h0;
		else
			\mchip.SERVO_2.eight_count [1] <= _421_[1];
	always @(posedge io_in[12])
		if (_005_)
			\mchip.SERVO_2.eight_count [2] <= 1'h0;
		else
			\mchip.SERVO_2.eight_count [2] <= _421_[2];
	always @(posedge io_in[12])
		if (_005_)
			\mchip.SERVO_2.eight_count [3] <= 1'h0;
		else
			\mchip.SERVO_2.eight_count [3] <= _421_[3];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.SERVO_1.pwm.ctr_d [0] <= 1'h0;
		else
			\mchip.SERVO_1.pwm.ctr_d [0] <= _418_[0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.SERVO_1.pwm.ctr_d [1] <= 1'h0;
		else
			\mchip.SERVO_1.pwm.ctr_d [1] <= _419_[1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.SERVO_1.pwm.ctr_d [2] <= 1'h0;
		else
			\mchip.SERVO_1.pwm.ctr_d [2] <= _419_[2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.SERVO_1.pwm.ctr_d [3] <= 1'h0;
		else
			\mchip.SERVO_1.pwm.ctr_d [3] <= _419_[3];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.SERVO_1.pwm.ctr_d [4] <= 1'h0;
		else
			\mchip.SERVO_1.pwm.ctr_d [4] <= _419_[4];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.SERVO_1.pwm.ctr_d [5] <= 1'h0;
		else
			\mchip.SERVO_1.pwm.ctr_d [5] <= _419_[5];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.SERVO_1.pwm.ctr_d [6] <= 1'h0;
		else
			\mchip.SERVO_1.pwm.ctr_d [6] <= _419_[6];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.SERVO_1.pwm.ctr_d [7] <= 1'h0;
		else
			\mchip.SERVO_1.pwm.ctr_d [7] <= _419_[7];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.SERVO_1.pwm.ctr_d [8] <= 1'h0;
		else
			\mchip.SERVO_1.pwm.ctr_d [8] <= _419_[8];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.SERVO_1.pwm.ctr_d [9] <= 1'h0;
		else
			\mchip.SERVO_1.pwm.ctr_d [9] <= _419_[9];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.SERVO_1.pwm.ctr_d [10] <= 1'h0;
		else
			\mchip.SERVO_1.pwm.ctr_d [10] <= _419_[10];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.SERVO_1.pwm.ctr_d [11] <= 1'h0;
		else
			\mchip.SERVO_1.pwm.ctr_d [11] <= _419_[11];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.SERVO_1.pwm.ctr_d [12] <= 1'h0;
		else
			\mchip.SERVO_1.pwm.ctr_d [12] <= _419_[12];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.SERVO_1.pwm.ctr_d [13] <= 1'h0;
		else
			\mchip.SERVO_1.pwm.ctr_d [13] <= _419_[13];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.SERVO_1.pwm.ctr_d [14] <= 1'h0;
		else
			\mchip.SERVO_1.pwm.ctr_d [14] <= _419_[14];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.SERVO_1.pwm.ctr_d [15] <= 1'h0;
		else
			\mchip.SERVO_1.pwm.ctr_d [15] <= _419_[15];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.SERVO_1.pwm.ctr_d [16] <= 1'h0;
		else
			\mchip.SERVO_1.pwm.ctr_d [16] <= _419_[16];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.SERVO_1.pwm.ctr_d [17] <= 1'h0;
		else
			\mchip.SERVO_1.pwm.ctr_d [17] <= _419_[17];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.SERVO_1.pwm.ctr_d [18] <= 1'h0;
		else
			\mchip.SERVO_1.pwm.ctr_d [18] <= _419_[18];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.SERVO_1.pwm.ctr_d [19] <= 1'h0;
		else
			\mchip.SERVO_1.pwm.ctr_d [19] <= _419_[19];
	always @(posedge io_in[12]) \mchip.SERVO_1.last_in_clk  <= io_in[11];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DECODE_2.p  <= 1'h0;
		else
			\mchip.DECODE_2.p  <= _010_;
	always @(posedge io_in[12])
		if (_003_)
			\mchip.SERVO_1.shreg [0] <= io_in[4];
	always @(posedge io_in[12])
		if (_003_)
			\mchip.SERVO_1.shreg [1] <= \mchip.SERVO_1.shreg [0];
	always @(posedge io_in[12])
		if (_003_)
			\mchip.SERVO_1.shreg [2] <= \mchip.SERVO_1.shreg [1];
	always @(posedge io_in[12])
		if (_003_)
			\mchip.SERVO_1.shreg [3] <= \mchip.SERVO_1.shreg [2];
	always @(posedge io_in[12])
		if (_003_)
			\mchip.SERVO_1.shreg [4] <= \mchip.SERVO_1.shreg [3];
	always @(posedge io_in[12])
		if (_003_)
			\mchip.SERVO_1.shreg [5] <= \mchip.SERVO_1.shreg [4];
	always @(posedge io_in[12])
		if (_003_)
			\mchip.SERVO_1.shreg [6] <= \mchip.SERVO_1.shreg [5];
	always @(posedge io_in[12])
		if (_003_)
			\mchip.SERVO_1.shreg [7] <= \mchip.SERVO_1.shreg [6];
	always @(posedge io_in[12])
		if (_004_)
			\mchip.SERVO_1.position [0] <= \mchip.SERVO_1.shreg [0];
	always @(posedge io_in[12])
		if (_004_)
			\mchip.SERVO_1.position [1] <= \mchip.SERVO_1.shreg [1];
	always @(posedge io_in[12])
		if (_004_)
			\mchip.SERVO_1.position [2] <= \mchip.SERVO_1.shreg [2];
	always @(posedge io_in[12])
		if (_004_)
			\mchip.SERVO_1.position [3] <= \mchip.SERVO_1.shreg [3];
	always @(posedge io_in[12])
		if (_004_)
			\mchip.SERVO_1.position [4] <= \mchip.SERVO_1.shreg [4];
	always @(posedge io_in[12])
		if (_004_)
			\mchip.SERVO_1.position [5] <= \mchip.SERVO_1.shreg [5];
	always @(posedge io_in[12])
		if (_004_)
			\mchip.SERVO_1.position [6] <= \mchip.SERVO_1.shreg [6];
	always @(posedge io_in[12])
		if (_004_)
			\mchip.SERVO_1.position [7] <= \mchip.SERVO_1.shreg [7];
	always @(posedge io_in[12])
		if (_006_)
			\mchip.SERVO_1.eight_count [0] <= 1'h0;
		else
			\mchip.SERVO_1.eight_count [0] <= _416_[0];
	always @(posedge io_in[12])
		if (_006_)
			\mchip.SERVO_1.eight_count [1] <= 1'h0;
		else
			\mchip.SERVO_1.eight_count [1] <= _417_[1];
	always @(posedge io_in[12])
		if (_006_)
			\mchip.SERVO_1.eight_count [2] <= 1'h0;
		else
			\mchip.SERVO_1.eight_count [2] <= _417_[2];
	always @(posedge io_in[12])
		if (_006_)
			\mchip.SERVO_1.eight_count [3] <= 1'h0;
		else
			\mchip.SERVO_1.eight_count [3] <= _417_[3];
	assign _416_[3:1] = \mchip.SERVO_1.eight_count [3:1];
	assign _417_[0] = _416_[0];
	assign _418_[19:1] = 19'h00000;
	assign _419_[0] = _418_[0];
	assign _420_[3:1] = \mchip.SERVO_2.eight_count [3:1];
	assign _421_[0] = _420_[0];
	assign _422_[19:1] = 19'h00000;
	assign _423_[0] = _422_[0];
	assign io_out = {6'h00, \mchip.DECODE_2.dir , \mchip.DECODE_2.p , \mchip.DECODE_1.dir , \mchip.DECODE_1.p , \mchip.SERVO_2.pwm.servo , \mchip.SERVO_1.pwm.servo , 2'h0};
	assign \mchip.DECODE_1.A  = io_in[6];
	assign \mchip.DECODE_1.B  = io_in[7];
	assign \mchip.DECODE_1.clock  = io_in[12];
	assign \mchip.DECODE_1.reset  = io_in[13];
	assign \mchip.DECODE_2.A  = io_in[8];
	assign \mchip.DECODE_2.B  = io_in[9];
	assign \mchip.DECODE_2.clock  = io_in[12];
	assign \mchip.DECODE_2.reset  = io_in[13];
	assign \mchip.PWM_1.CLK  = io_in[12];
	assign \mchip.PWM_1.M_OUT  = 1'h0;
	assign \mchip.PWM_1.PWM_DUTY  = io_in[1];
	assign \mchip.PWM_1.PWM_PERIOD  = io_in[0];
	assign \mchip.PWM_1.SCL  = io_in[11];
	assign \mchip.PWM_1.reset  = io_in[13];
	assign \mchip.PWM_2.CLK  = io_in[12];
	assign \mchip.PWM_2.M_OUT  = 1'h0;
	assign \mchip.PWM_2.PWM_DUTY  = io_in[3];
	assign \mchip.PWM_2.PWM_PERIOD  = io_in[2];
	assign \mchip.PWM_2.SCL  = io_in[11];
	assign \mchip.PWM_2.reset  = io_in[13];
	assign \mchip.SERVO_1.CLK  = io_in[12];
	assign \mchip.SERVO_1.SCL  = io_in[11];
	assign \mchip.SERVO_1.S_IN  = io_in[4];
	assign \mchip.SERVO_1.S_OUT  = \mchip.SERVO_1.pwm.servo ;
	assign \mchip.SERVO_1.pwm.clk  = io_in[12];
	assign \mchip.SERVO_1.pwm.position  = \mchip.SERVO_1.position ;
	assign \mchip.SERVO_1.pwm.rst  = io_in[13];
	assign \mchip.SERVO_1.pwm.temp_val  = 20'h00000;
	assign \mchip.SERVO_1.reset  = io_in[13];
	assign \mchip.SERVO_2.CLK  = io_in[12];
	assign \mchip.SERVO_2.SCL  = io_in[11];
	assign \mchip.SERVO_2.S_IN  = io_in[5];
	assign \mchip.SERVO_2.S_OUT  = \mchip.SERVO_2.pwm.servo ;
	assign \mchip.SERVO_2.last_in_clk  = \mchip.SERVO_1.last_in_clk ;
	assign \mchip.SERVO_2.pwm.clk  = io_in[12];
	assign \mchip.SERVO_2.pwm.position  = \mchip.SERVO_2.position ;
	assign \mchip.SERVO_2.pwm.rst  = io_in[13];
	assign \mchip.SERVO_2.pwm.temp_val  = 20'h00000;
	assign \mchip.SERVO_2.reset  = io_in[13];
	assign \mchip.clock  = io_in[12];
	assign \mchip.io_in  = io_in[11:0];
	assign \mchip.io_out  = {4'h0, \mchip.DECODE_2.dir , \mchip.DECODE_2.p , \mchip.DECODE_1.dir , \mchip.DECODE_1.p , \mchip.SERVO_2.pwm.servo , \mchip.SERVO_1.pwm.servo , 2'h0};
	assign \mchip.reset  = io_in[13];
endmodule
module d22_yushuanl_convolution (
	io_in,
	io_out
);
	wire [2:0] _00_;
	wire _01_;
	wire _02_;
	wire _03_;
	wire _04_;
	wire _05_;
	wire _06_;
	wire _07_;
	wire _08_;
	wire _09_;
	wire _10_;
	wire _11_;
	wire _12_;
	wire _13_;
	wire _14_;
	wire _15_;
	wire _16_;
	wire _17_;
	wire _18_;
	wire _19_;
	wire _20_;
	wire _21_;
	wire _22_;
	wire _23_;
	wire _24_;
	wire _25_;
	wire _26_;
	wire _27_;
	wire _28_;
	wire _29_;
	input wire [13:0] io_in;
	output wire [13:0] io_out;
	wire [5:0] \mchip.Shifted_A ;
	wire [5:0] \mchip.Shifted_B ;
	wire [3:0] \mchip.add.Out ;
	wire \mchip.clock ;
	reg [2:0] \mchip.curState ;
	wire \mchip.enRO ;
	wire \mchip.enRT ;
	wire [3:0] \mchip.inReg ;
	wire [11:0] \mchip.io_in ;
	wire [3:0] \mchip.io_out ;
	wire \mchip.mul.First ;
	wire \mchip.mul.Second ;
	wire [3:0] \mchip.mux.A ;
	wire [3:0] \mchip.mux.B ;
	wire [3:0] \mchip.oldSum ;
	wire [3:0] \mchip.registerOut.In ;
	reg [3:0] \mchip.registerOut.Out ;
	wire \mchip.registerOut.clk ;
	wire \mchip.registerOut.en ;
	wire [3:0] \mchip.registerTemp.In ;
	reg [3:0] \mchip.registerTemp.Out ;
	wire \mchip.registerTemp.clk ;
	wire \mchip.registerTemp.en ;
	wire \mchip.reset ;
	wire [5:0] \mchip.shiftA.In ;
	reg [5:0] \mchip.shiftA.Shifted ;
	wire \mchip.shiftA.clk ;
	wire [5:0] \mchip.shiftB.In ;
	reg [5:0] \mchip.shiftB.Shifted ;
	wire \mchip.shiftB.clk ;
	assign _12_ = ~(\mchip.curState [1] | \mchip.curState [0]);
	assign _13_ = _12_ & ~\mchip.curState [2];
	assign _14_ = ~\mchip.curState [2];
	assign _15_ = \mchip.curState [1] & \mchip.curState [0];
	assign _16_ = (\mchip.curState [2] ? _15_ : _12_);
	assign _01_ = _13_ | ~_16_;
	assign _17_ = ~_15_;
	assign _18_ = \mchip.curState [1] | ~\mchip.curState [0];
	assign \mchip.enRT  = (\mchip.curState [2] ? _17_ : _18_);
	assign \mchip.enRO  = _15_ & ~_14_;
	assign _07_ = (_13_ ? io_in[6] : \mchip.shiftB.Shifted [1]);
	assign _08_ = (_13_ ? io_in[7] : \mchip.shiftB.Shifted [2]);
	assign _09_ = (_13_ ? io_in[8] : \mchip.shiftB.Shifted [3]);
	assign _10_ = (_13_ ? io_in[9] : \mchip.shiftB.Shifted [4]);
	assign _11_ = (_13_ ? io_in[10] : \mchip.shiftB.Shifted [5]);
	assign _02_ = (_13_ ? io_in[0] : \mchip.shiftA.Shifted [1]);
	assign _03_ = (_13_ ? io_in[1] : \mchip.shiftA.Shifted [2]);
	assign _04_ = (_13_ ? io_in[2] : \mchip.shiftA.Shifted [3]);
	assign _05_ = (_13_ ? io_in[3] : \mchip.shiftA.Shifted [4]);
	assign _06_ = (_13_ ? io_in[4] : \mchip.shiftA.Shifted [5]);
	assign _19_ = ~\mchip.curState [0];
	assign _00_[0] = (\mchip.curState [2] ? _18_ : _19_);
	assign _20_ = ~_12_;
	assign _21_ = \mchip.curState [1] ^ \mchip.curState [0];
	assign _00_[1] = (\mchip.curState [2] ? _20_ : _21_);
	assign _00_[2] = _15_ | \mchip.curState [2];
	assign _22_ = \mchip.registerTemp.Out [0] & ~_16_;
	assign _23_ = ~(\mchip.shiftA.Shifted [0] & \mchip.shiftB.Shifted [0]);
	assign _24_ = _22_ & ~_23_;
	assign _25_ = _16_ | ~\mchip.registerTemp.Out [1];
	assign \mchip.registerTemp.In [1] = ~(_25_ ^ _24_);
	assign _26_ = _24_ & ~_25_;
	assign _27_ = _16_ | ~\mchip.registerTemp.Out [2];
	assign \mchip.registerTemp.In [2] = ~(_27_ ^ _26_);
	assign _28_ = _26_ & ~_27_;
	assign _29_ = \mchip.registerTemp.Out [3] & ~_16_;
	assign \mchip.registerTemp.In [3] = _29_ ^ _28_;
	assign \mchip.registerTemp.In [0] = ~(_23_ ^ _22_);
	always @(posedge io_in[12])
		if (_01_)
			if (!_13_)
				\mchip.shiftA.Shifted [5] <= 1'h0;
			else
				\mchip.shiftA.Shifted [5] <= io_in[5];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.curState [0] <= 1'h0;
		else
			\mchip.curState [0] <= _00_[0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.curState [1] <= 1'h0;
		else
			\mchip.curState [1] <= _00_[1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.curState [2] <= 1'h0;
		else
			\mchip.curState [2] <= _00_[2];
	always @(posedge io_in[12])
		if (_01_)
			\mchip.shiftA.Shifted [0] <= _02_;
	always @(posedge io_in[12])
		if (_01_)
			\mchip.shiftA.Shifted [1] <= _03_;
	always @(posedge io_in[12])
		if (_01_)
			\mchip.shiftA.Shifted [2] <= _04_;
	always @(posedge io_in[12])
		if (_01_)
			\mchip.shiftA.Shifted [3] <= _05_;
	always @(posedge io_in[12])
		if (_01_)
			\mchip.shiftA.Shifted [4] <= _06_;
	always @(posedge io_in[12])
		if (_01_)
			\mchip.shiftB.Shifted [0] <= _07_;
	always @(posedge io_in[12])
		if (_01_)
			\mchip.shiftB.Shifted [1] <= _08_;
	always @(posedge io_in[12])
		if (_01_)
			\mchip.shiftB.Shifted [2] <= _09_;
	always @(posedge io_in[12])
		if (_01_)
			\mchip.shiftB.Shifted [3] <= _10_;
	always @(posedge io_in[12])
		if (_01_)
			\mchip.shiftB.Shifted [4] <= _11_;
	always @(posedge io_in[12])
		if (\mchip.enRO )
			\mchip.registerOut.Out [0] <= \mchip.registerTemp.Out [0];
	always @(posedge io_in[12])
		if (\mchip.enRO )
			\mchip.registerOut.Out [1] <= \mchip.registerTemp.Out [1];
	always @(posedge io_in[12])
		if (\mchip.enRO )
			\mchip.registerOut.Out [2] <= \mchip.registerTemp.Out [2];
	always @(posedge io_in[12])
		if (\mchip.enRO )
			\mchip.registerOut.Out [3] <= \mchip.registerTemp.Out [3];
	always @(posedge io_in[12])
		if (_01_)
			if (!_13_)
				\mchip.shiftB.Shifted [5] <= 1'h0;
			else
				\mchip.shiftB.Shifted [5] <= io_in[11];
	always @(posedge io_in[12])
		if (\mchip.enRT )
			\mchip.registerTemp.Out [0] <= \mchip.registerTemp.In [0];
	always @(posedge io_in[12])
		if (\mchip.enRT )
			\mchip.registerTemp.Out [1] <= \mchip.registerTemp.In [1];
	always @(posedge io_in[12])
		if (\mchip.enRT )
			\mchip.registerTemp.Out [2] <= \mchip.registerTemp.In [2];
	always @(posedge io_in[12])
		if (\mchip.enRT )
			\mchip.registerTemp.Out [3] <= \mchip.registerTemp.In [3];
	assign io_out = {10'h000, \mchip.registerOut.Out };
	assign \mchip.Shifted_A  = \mchip.shiftA.Shifted ;
	assign \mchip.Shifted_B  = \mchip.shiftB.Shifted ;
	assign \mchip.add.Out  = \mchip.registerTemp.In ;
	assign \mchip.clock  = io_in[12];
	assign \mchip.inReg  = \mchip.registerTemp.In ;
	assign \mchip.io_in  = io_in[11:0];
	assign \mchip.io_out  = \mchip.registerOut.Out ;
	assign \mchip.mul.First  = \mchip.shiftA.Shifted [0];
	assign \mchip.mul.Second  = \mchip.shiftB.Shifted [0];
	assign \mchip.mux.A  = \mchip.registerTemp.Out ;
	assign \mchip.mux.B  = 4'h0;
	assign \mchip.oldSum  = \mchip.registerTemp.Out ;
	assign \mchip.registerOut.In  = \mchip.registerTemp.Out ;
	assign \mchip.registerOut.clk  = io_in[12];
	assign \mchip.registerOut.en  = \mchip.enRO ;
	assign \mchip.registerTemp.clk  = io_in[12];
	assign \mchip.registerTemp.en  = \mchip.enRT ;
	assign \mchip.reset  = io_in[13];
	assign \mchip.shiftA.In  = io_in[5:0];
	assign \mchip.shiftA.clk  = io_in[12];
	assign \mchip.shiftB.In  = io_in[11:6];
	assign \mchip.shiftB.clk  = io_in[12];
endmodule
module d23_zhiyingm_turing (
	io_in,
	io_out
);
	wire _0000_;
	wire _0001_;
	wire _0002_;
	wire _0003_;
	wire _0004_;
	wire _0005_;
	wire _0006_;
	wire _0007_;
	wire _0008_;
	wire _0009_;
	wire _0010_;
	wire _0011_;
	wire _0012_;
	wire _0013_;
	wire _0014_;
	wire _0015_;
	wire _0016_;
	wire _0017_;
	wire _0018_;
	wire _0019_;
	wire _0020_;
	wire _0021_;
	wire _0022_;
	wire _0023_;
	wire _0024_;
	wire _0025_;
	wire _0026_;
	wire _0027_;
	wire _0028_;
	wire _0029_;
	wire _0030_;
	wire _0031_;
	wire _0032_;
	wire _0033_;
	wire _0034_;
	wire _0035_;
	wire _0036_;
	wire _0037_;
	wire _0038_;
	wire _0039_;
	wire _0040_;
	wire _0041_;
	wire _0042_;
	wire _0043_;
	wire _0044_;
	wire _0045_;
	wire _0046_;
	wire _0047_;
	wire _0048_;
	wire _0049_;
	wire _0050_;
	wire _0051_;
	wire _0052_;
	wire _0053_;
	wire _0054_;
	wire _0055_;
	wire _0056_;
	wire _0057_;
	wire _0058_;
	wire _0059_;
	wire _0060_;
	wire _0061_;
	wire _0062_;
	wire _0063_;
	wire _0064_;
	wire _0065_;
	wire _0066_;
	wire _0067_;
	wire _0068_;
	wire _0069_;
	wire _0070_;
	wire _0071_;
	wire _0072_;
	wire _0073_;
	wire _0074_;
	wire _0075_;
	wire _0076_;
	wire _0077_;
	wire _0078_;
	wire _0079_;
	wire _0080_;
	wire _0081_;
	wire _0082_;
	wire _0083_;
	wire _0084_;
	wire _0085_;
	wire _0086_;
	wire _0087_;
	wire _0088_;
	wire _0089_;
	wire _0090_;
	wire _0091_;
	wire _0092_;
	wire _0093_;
	wire _0094_;
	wire _0095_;
	wire _0096_;
	wire _0097_;
	wire _0098_;
	wire _0099_;
	wire _0100_;
	wire _0101_;
	wire _0102_;
	wire _0103_;
	wire _0104_;
	wire _0105_;
	wire _0106_;
	wire _0107_;
	wire _0108_;
	wire _0109_;
	wire _0110_;
	wire _0111_;
	wire _0112_;
	wire _0113_;
	wire _0114_;
	wire _0115_;
	wire _0116_;
	wire _0117_;
	wire _0118_;
	wire _0119_;
	wire _0120_;
	wire _0121_;
	wire _0122_;
	wire _0123_;
	wire _0124_;
	wire _0125_;
	wire _0126_;
	wire _0127_;
	wire _0128_;
	wire _0129_;
	wire _0130_;
	wire _0131_;
	wire _0132_;
	wire _0133_;
	wire _0134_;
	wire _0135_;
	wire _0136_;
	wire _0137_;
	wire _0138_;
	wire _0139_;
	wire _0140_;
	wire _0141_;
	wire _0142_;
	wire _0143_;
	wire _0144_;
	wire _0145_;
	wire _0146_;
	wire _0147_;
	wire _0148_;
	wire _0149_;
	wire _0150_;
	wire _0151_;
	wire _0152_;
	wire _0153_;
	wire _0154_;
	wire _0155_;
	wire _0156_;
	wire _0157_;
	wire _0158_;
	wire _0159_;
	wire _0160_;
	wire _0161_;
	wire _0162_;
	wire _0163_;
	wire _0164_;
	wire _0165_;
	wire _0166_;
	wire _0167_;
	wire _0168_;
	wire _0169_;
	wire _0170_;
	wire _0171_;
	wire _0172_;
	wire _0173_;
	wire _0174_;
	wire _0175_;
	wire _0176_;
	wire _0177_;
	wire _0178_;
	wire _0179_;
	wire _0180_;
	wire _0181_;
	wire _0182_;
	wire _0183_;
	wire _0184_;
	wire _0185_;
	wire _0186_;
	wire _0187_;
	wire _0188_;
	wire _0189_;
	wire _0190_;
	wire _0191_;
	wire _0192_;
	wire _0193_;
	wire _0194_;
	wire _0195_;
	wire _0196_;
	wire _0197_;
	wire _0198_;
	wire _0199_;
	wire _0200_;
	wire _0201_;
	wire _0202_;
	wire _0203_;
	wire _0204_;
	wire _0205_;
	wire _0206_;
	wire _0207_;
	wire _0208_;
	wire _0209_;
	wire _0210_;
	wire _0211_;
	wire _0212_;
	wire _0213_;
	wire _0214_;
	wire _0215_;
	wire _0216_;
	wire _0217_;
	wire _0218_;
	wire _0219_;
	wire _0220_;
	wire _0221_;
	wire _0222_;
	wire _0223_;
	wire _0224_;
	wire _0225_;
	wire _0226_;
	wire _0227_;
	wire _0228_;
	wire _0229_;
	wire _0230_;
	wire _0231_;
	wire _0232_;
	wire _0233_;
	wire _0234_;
	wire _0235_;
	wire _0236_;
	wire _0237_;
	wire _0238_;
	wire _0239_;
	wire _0240_;
	wire _0241_;
	wire _0242_;
	wire _0243_;
	wire _0244_;
	wire _0245_;
	wire _0246_;
	wire _0247_;
	wire _0248_;
	wire _0249_;
	wire _0250_;
	wire _0251_;
	wire _0252_;
	wire _0253_;
	wire _0254_;
	wire _0255_;
	wire _0256_;
	wire _0257_;
	wire _0258_;
	wire _0259_;
	wire _0260_;
	wire _0261_;
	wire _0262_;
	wire _0263_;
	wire _0264_;
	wire _0265_;
	wire _0266_;
	wire _0267_;
	wire _0268_;
	wire _0269_;
	wire _0270_;
	wire _0271_;
	wire _0272_;
	wire _0273_;
	wire _0274_;
	wire _0275_;
	wire _0276_;
	wire _0277_;
	wire _0278_;
	wire _0279_;
	wire _0280_;
	wire _0281_;
	wire _0282_;
	wire _0283_;
	wire _0284_;
	wire _0285_;
	wire _0286_;
	wire _0287_;
	wire _0288_;
	wire _0289_;
	wire _0290_;
	wire _0291_;
	wire _0292_;
	wire _0293_;
	wire _0294_;
	wire _0295_;
	wire _0296_;
	wire _0297_;
	wire _0298_;
	wire _0299_;
	wire _0300_;
	wire _0301_;
	wire _0302_;
	wire _0303_;
	wire _0304_;
	wire _0305_;
	wire _0306_;
	wire _0307_;
	wire _0308_;
	wire _0309_;
	wire _0310_;
	wire _0311_;
	wire _0312_;
	wire _0313_;
	wire _0314_;
	wire _0315_;
	wire _0316_;
	wire _0317_;
	wire _0318_;
	wire _0319_;
	wire _0320_;
	wire _0321_;
	wire _0322_;
	wire _0323_;
	wire _0324_;
	wire _0325_;
	wire _0326_;
	wire _0327_;
	wire _0328_;
	wire _0329_;
	wire _0330_;
	wire _0331_;
	wire _0332_;
	wire _0333_;
	wire _0334_;
	wire _0335_;
	wire _0336_;
	wire _0337_;
	wire _0338_;
	wire _0339_;
	wire _0340_;
	wire _0341_;
	wire _0342_;
	wire _0343_;
	wire _0344_;
	wire _0345_;
	wire _0346_;
	wire _0347_;
	wire _0348_;
	wire _0349_;
	wire _0350_;
	wire _0351_;
	wire _0352_;
	wire _0353_;
	wire _0354_;
	wire _0355_;
	wire _0356_;
	wire _0357_;
	wire _0358_;
	wire _0359_;
	wire _0360_;
	wire _0361_;
	wire _0362_;
	wire _0363_;
	wire _0364_;
	wire _0365_;
	wire _0366_;
	wire _0367_;
	wire _0368_;
	wire _0369_;
	wire _0370_;
	wire _0371_;
	wire _0372_;
	wire _0373_;
	wire _0374_;
	wire _0375_;
	wire _0376_;
	wire _0377_;
	wire _0378_;
	wire _0379_;
	wire _0380_;
	wire _0381_;
	wire _0382_;
	wire _0383_;
	wire _0384_;
	wire _0385_;
	wire _0386_;
	wire _0387_;
	wire _0388_;
	wire _0389_;
	wire _0390_;
	wire _0391_;
	wire _0392_;
	wire _0393_;
	wire _0394_;
	wire _0395_;
	wire _0396_;
	wire _0397_;
	wire _0398_;
	wire _0399_;
	wire _0400_;
	wire _0401_;
	wire _0402_;
	wire _0403_;
	wire _0404_;
	wire _0405_;
	wire _0406_;
	wire _0407_;
	wire _0408_;
	wire _0409_;
	wire _0410_;
	wire _0411_;
	wire _0412_;
	wire _0413_;
	wire _0414_;
	wire _0415_;
	wire _0416_;
	wire _0417_;
	wire _0418_;
	wire _0419_;
	wire _0420_;
	wire _0421_;
	wire _0422_;
	wire _0423_;
	wire _0424_;
	wire _0425_;
	wire _0426_;
	wire _0427_;
	wire _0428_;
	wire _0429_;
	wire _0430_;
	wire _0431_;
	wire _0432_;
	wire _0433_;
	wire _0434_;
	wire _0435_;
	wire _0436_;
	wire _0437_;
	wire _0438_;
	wire _0439_;
	wire _0440_;
	wire _0441_;
	wire _0442_;
	wire _0443_;
	wire _0444_;
	wire _0445_;
	wire _0446_;
	wire _0447_;
	wire _0448_;
	wire _0449_;
	wire _0450_;
	wire _0451_;
	wire _0452_;
	wire _0453_;
	wire _0454_;
	wire _0455_;
	wire _0456_;
	wire _0457_;
	wire _0458_;
	wire _0459_;
	wire _0460_;
	wire _0461_;
	wire _0462_;
	wire _0463_;
	wire _0464_;
	wire _0465_;
	wire _0466_;
	wire _0467_;
	wire _0468_;
	wire _0469_;
	wire _0470_;
	wire _0471_;
	wire _0472_;
	wire _0473_;
	wire _0474_;
	wire _0475_;
	wire _0476_;
	wire _0477_;
	wire _0478_;
	wire _0479_;
	wire _0480_;
	wire _0481_;
	wire _0482_;
	wire _0483_;
	wire _0484_;
	wire _0485_;
	wire _0486_;
	wire _0487_;
	wire _0488_;
	wire _0489_;
	wire _0490_;
	wire _0491_;
	wire _0492_;
	wire _0493_;
	wire _0494_;
	wire _0495_;
	wire _0496_;
	wire _0497_;
	wire _0498_;
	wire _0499_;
	wire _0500_;
	wire _0501_;
	wire _0502_;
	wire _0503_;
	wire _0504_;
	wire _0505_;
	wire _0506_;
	wire _0507_;
	wire _0508_;
	wire _0509_;
	wire _0510_;
	wire _0511_;
	wire _0512_;
	wire _0513_;
	wire _0514_;
	wire _0515_;
	wire _0516_;
	wire _0517_;
	wire _0518_;
	wire _0519_;
	wire _0520_;
	wire _0521_;
	wire _0522_;
	wire _0523_;
	wire _0524_;
	wire _0525_;
	wire _0526_;
	wire _0527_;
	wire _0528_;
	wire _0529_;
	wire _0530_;
	wire _0531_;
	wire _0532_;
	wire _0533_;
	wire _0534_;
	wire _0535_;
	wire _0536_;
	wire _0537_;
	wire _0538_;
	wire _0539_;
	wire _0540_;
	wire _0541_;
	wire _0542_;
	wire _0543_;
	wire _0544_;
	wire _0545_;
	wire _0546_;
	wire _0547_;
	wire _0548_;
	wire _0549_;
	wire _0550_;
	wire _0551_;
	wire _0552_;
	wire _0553_;
	wire _0554_;
	wire _0555_;
	wire _0556_;
	wire _0557_;
	wire _0558_;
	wire _0559_;
	wire _0560_;
	wire _0561_;
	wire _0562_;
	wire _0563_;
	wire _0564_;
	wire _0565_;
	wire _0566_;
	wire _0567_;
	wire _0568_;
	wire _0569_;
	wire _0570_;
	wire _0571_;
	wire _0572_;
	wire _0573_;
	wire _0574_;
	wire _0575_;
	wire _0576_;
	wire _0577_;
	wire _0578_;
	wire _0579_;
	wire _0580_;
	wire _0581_;
	wire _0582_;
	wire _0583_;
	wire _0584_;
	wire _0585_;
	wire _0586_;
	wire _0587_;
	wire _0588_;
	wire _0589_;
	wire _0590_;
	wire _0591_;
	wire _0592_;
	wire _0593_;
	wire _0594_;
	wire _0595_;
	wire _0596_;
	wire _0597_;
	wire _0598_;
	wire _0599_;
	wire _0600_;
	wire _0601_;
	wire _0602_;
	wire _0603_;
	wire _0604_;
	wire _0605_;
	wire _0606_;
	wire _0607_;
	wire _0608_;
	wire _0609_;
	wire _0610_;
	wire _0611_;
	wire _0612_;
	wire _0613_;
	wire _0614_;
	wire _0615_;
	wire _0616_;
	wire _0617_;
	wire _0618_;
	wire _0619_;
	wire _0620_;
	wire _0621_;
	wire _0622_;
	wire _0623_;
	wire _0624_;
	wire _0625_;
	wire _0626_;
	wire _0627_;
	wire _0628_;
	wire _0629_;
	wire _0630_;
	wire _0631_;
	wire _0632_;
	wire _0633_;
	wire _0634_;
	wire _0635_;
	wire _0636_;
	wire _0637_;
	wire _0638_;
	wire _0639_;
	wire _0640_;
	wire _0641_;
	wire _0642_;
	wire _0643_;
	wire _0644_;
	wire _0645_;
	wire _0646_;
	wire _0647_;
	wire _0648_;
	wire _0649_;
	wire _0650_;
	wire _0651_;
	wire _0652_;
	wire _0653_;
	wire _0654_;
	wire _0655_;
	wire _0656_;
	wire _0657_;
	wire _0658_;
	wire _0659_;
	wire _0660_;
	wire _0661_;
	wire _0662_;
	wire _0663_;
	wire _0664_;
	wire _0665_;
	wire _0666_;
	wire _0667_;
	wire _0668_;
	wire _0669_;
	wire _0670_;
	wire _0671_;
	wire _0672_;
	wire _0673_;
	wire _0674_;
	wire _0675_;
	wire _0676_;
	wire _0677_;
	wire _0678_;
	wire _0679_;
	wire _0680_;
	wire _0681_;
	wire _0682_;
	wire _0683_;
	wire _0684_;
	wire _0685_;
	wire _0686_;
	wire _0687_;
	wire _0688_;
	wire _0689_;
	wire _0690_;
	wire _0691_;
	wire _0692_;
	wire _0693_;
	wire _0694_;
	wire _0695_;
	wire _0696_;
	wire _0697_;
	wire _0698_;
	wire _0699_;
	wire _0700_;
	wire _0701_;
	wire _0702_;
	wire _0703_;
	wire _0704_;
	wire _0705_;
	wire _0706_;
	wire _0707_;
	wire _0708_;
	wire _0709_;
	wire _0710_;
	wire _0711_;
	wire _0712_;
	wire _0713_;
	wire _0714_;
	wire _0715_;
	wire _0716_;
	wire _0717_;
	wire _0718_;
	wire _0719_;
	wire _0720_;
	wire _0721_;
	wire _0722_;
	wire _0723_;
	wire _0724_;
	wire _0725_;
	wire _0726_;
	wire _0727_;
	wire _0728_;
	wire _0729_;
	wire _0730_;
	wire _0731_;
	wire _0732_;
	wire _0733_;
	wire _0734_;
	wire _0735_;
	wire _0736_;
	wire _0737_;
	wire _0738_;
	wire _0739_;
	wire _0740_;
	wire _0741_;
	wire _0742_;
	wire _0743_;
	wire _0744_;
	wire _0745_;
	wire _0746_;
	wire _0747_;
	wire _0748_;
	wire _0749_;
	wire _0750_;
	wire _0751_;
	wire _0752_;
	wire _0753_;
	wire _0754_;
	wire _0755_;
	wire _0756_;
	wire _0757_;
	wire _0758_;
	wire _0759_;
	wire _0760_;
	wire _0761_;
	wire _0762_;
	wire _0763_;
	wire _0764_;
	wire _0765_;
	wire _0766_;
	wire _0767_;
	wire _0768_;
	wire _0769_;
	wire _0770_;
	wire _0771_;
	wire _0772_;
	wire _0773_;
	wire _0774_;
	wire _0775_;
	wire _0776_;
	wire _0777_;
	wire _0778_;
	wire _0779_;
	wire _0780_;
	wire _0781_;
	wire _0782_;
	wire _0783_;
	wire _0784_;
	wire _0785_;
	wire _0786_;
	wire _0787_;
	wire _0788_;
	wire _0789_;
	wire _0790_;
	wire _0791_;
	wire _0792_;
	wire _0793_;
	wire _0794_;
	wire _0795_;
	wire _0796_;
	wire _0797_;
	wire _0798_;
	wire _0799_;
	wire _0800_;
	wire _0801_;
	wire _0802_;
	wire _0803_;
	wire _0804_;
	wire _0805_;
	wire _0806_;
	wire _0807_;
	wire _0808_;
	wire _0809_;
	wire _0810_;
	wire _0811_;
	wire _0812_;
	wire _0813_;
	wire _0814_;
	wire _0815_;
	wire _0816_;
	wire _0817_;
	wire _0818_;
	wire _0819_;
	wire _0820_;
	wire _0821_;
	wire _0822_;
	wire _0823_;
	wire _0824_;
	wire _0825_;
	wire _0826_;
	wire _0827_;
	wire _0828_;
	wire _0829_;
	wire _0830_;
	wire _0831_;
	wire _0832_;
	wire _0833_;
	wire _0834_;
	wire _0835_;
	wire _0836_;
	wire _0837_;
	wire _0838_;
	wire _0839_;
	wire _0840_;
	wire _0841_;
	wire _0842_;
	wire _0843_;
	wire _0844_;
	wire _0845_;
	wire _0846_;
	wire _0847_;
	wire _0848_;
	wire _0849_;
	wire _0850_;
	wire _0851_;
	wire _0852_;
	wire _0853_;
	wire _0854_;
	wire _0855_;
	wire _0856_;
	wire _0857_;
	wire _0858_;
	wire _0859_;
	wire _0860_;
	wire _0861_;
	wire _0862_;
	wire _0863_;
	wire _0864_;
	wire _0865_;
	wire _0866_;
	wire _0867_;
	wire _0868_;
	wire _0869_;
	wire _0870_;
	wire _0871_;
	wire _0872_;
	wire _0873_;
	wire _0874_;
	wire _0875_;
	wire _0876_;
	wire _0877_;
	wire _0878_;
	wire _0879_;
	wire _0880_;
	wire _0881_;
	wire _0882_;
	wire _0883_;
	wire _0884_;
	wire _0885_;
	wire _0886_;
	wire _0887_;
	wire _0888_;
	wire _0889_;
	wire _0890_;
	wire _0891_;
	wire _0892_;
	wire _0893_;
	wire _0894_;
	wire _0895_;
	wire _0896_;
	wire _0897_;
	wire _0898_;
	wire _0899_;
	wire _0900_;
	wire _0901_;
	wire _0902_;
	wire _0903_;
	wire _0904_;
	wire _0905_;
	wire _0906_;
	wire _0907_;
	wire _0908_;
	wire _0909_;
	wire _0910_;
	wire _0911_;
	wire _0912_;
	wire _0913_;
	wire _0914_;
	wire _0915_;
	wire _0916_;
	wire _0917_;
	wire _0918_;
	wire _0919_;
	wire _0920_;
	wire _0921_;
	wire _0922_;
	wire _0923_;
	wire _0924_;
	wire _0925_;
	wire _0926_;
	wire _0927_;
	wire _0928_;
	wire _0929_;
	wire _0930_;
	wire _0931_;
	wire _0932_;
	wire _0933_;
	wire _0934_;
	wire _0935_;
	wire _0936_;
	wire _0937_;
	wire _0938_;
	wire _0939_;
	wire _0940_;
	wire _0941_;
	wire _0942_;
	wire _0943_;
	wire _0944_;
	wire _0945_;
	wire _0946_;
	wire _0947_;
	wire _0948_;
	wire _0949_;
	wire _0950_;
	wire _0951_;
	wire _0952_;
	wire _0953_;
	wire _0954_;
	wire _0955_;
	wire _0956_;
	wire _0957_;
	wire _0958_;
	wire _0959_;
	wire _0960_;
	wire _0961_;
	wire _0962_;
	wire _0963_;
	wire _0964_;
	wire _0965_;
	wire _0966_;
	wire _0967_;
	wire _0968_;
	wire _0969_;
	wire _0970_;
	wire _0971_;
	wire _0972_;
	wire _0973_;
	wire _0974_;
	wire _0975_;
	wire _0976_;
	wire _0977_;
	wire _0978_;
	wire _0979_;
	wire _0980_;
	wire _0981_;
	wire _0982_;
	wire _0983_;
	wire _0984_;
	wire _0985_;
	wire _0986_;
	wire _0987_;
	wire _0988_;
	wire _0989_;
	wire _0990_;
	wire _0991_;
	wire _0992_;
	wire _0993_;
	wire _0994_;
	wire _0995_;
	wire _0996_;
	wire _0997_;
	wire _0998_;
	wire _0999_;
	wire _1000_;
	wire _1001_;
	wire _1002_;
	wire _1003_;
	wire _1004_;
	wire _1005_;
	wire _1006_;
	wire _1007_;
	wire _1008_;
	wire _1009_;
	wire _1010_;
	wire _1011_;
	wire _1012_;
	wire _1013_;
	wire _1014_;
	wire _1015_;
	wire _1016_;
	wire _1017_;
	wire _1018_;
	wire _1019_;
	wire _1020_;
	wire _1021_;
	wire _1022_;
	wire _1023_;
	wire _1024_;
	wire _1025_;
	wire _1026_;
	wire _1027_;
	wire _1028_;
	wire _1029_;
	wire _1030_;
	wire _1031_;
	wire _1032_;
	wire _1033_;
	wire _1034_;
	wire _1035_;
	wire _1036_;
	wire _1037_;
	wire _1038_;
	wire _1039_;
	wire _1040_;
	wire _1041_;
	wire _1042_;
	wire _1043_;
	wire _1044_;
	wire _1045_;
	wire _1046_;
	wire _1047_;
	wire _1048_;
	wire _1049_;
	wire _1050_;
	wire _1051_;
	wire _1052_;
	wire _1053_;
	wire _1054_;
	wire _1055_;
	wire _1056_;
	wire _1057_;
	wire _1058_;
	wire _1059_;
	wire _1060_;
	wire _1061_;
	wire _1062_;
	wire _1063_;
	wire _1064_;
	wire _1065_;
	wire _1066_;
	wire _1067_;
	wire _1068_;
	wire _1069_;
	wire _1070_;
	wire _1071_;
	wire _1072_;
	wire _1073_;
	wire _1074_;
	wire _1075_;
	wire _1076_;
	wire _1077_;
	wire _1078_;
	wire _1079_;
	wire _1080_;
	wire _1081_;
	wire _1082_;
	wire _1083_;
	wire _1084_;
	wire _1085_;
	wire _1086_;
	wire _1087_;
	wire _1088_;
	wire _1089_;
	wire _1090_;
	wire _1091_;
	wire _1092_;
	wire _1093_;
	wire _1094_;
	wire _1095_;
	wire _1096_;
	wire _1097_;
	wire _1098_;
	wire _1099_;
	wire _1100_;
	wire _1101_;
	wire _1102_;
	wire _1103_;
	wire _1104_;
	wire _1105_;
	wire _1106_;
	wire _1107_;
	wire _1108_;
	wire _1109_;
	wire _1110_;
	wire _1111_;
	wire _1112_;
	wire _1113_;
	wire _1114_;
	wire _1115_;
	wire _1116_;
	wire _1117_;
	wire _1118_;
	wire _1119_;
	wire _1120_;
	wire _1121_;
	wire _1122_;
	wire _1123_;
	wire _1124_;
	wire _1125_;
	wire _1126_;
	wire _1127_;
	wire _1128_;
	wire _1129_;
	wire _1130_;
	wire _1131_;
	wire _1132_;
	wire _1133_;
	wire _1134_;
	wire _1135_;
	wire _1136_;
	wire _1137_;
	wire _1138_;
	wire _1139_;
	wire _1140_;
	wire _1141_;
	wire _1142_;
	wire _1143_;
	wire _1144_;
	wire _1145_;
	wire _1146_;
	wire _1147_;
	wire _1148_;
	wire _1149_;
	wire _1150_;
	wire _1151_;
	wire _1152_;
	wire _1153_;
	wire _1154_;
	wire _1155_;
	wire _1156_;
	wire _1157_;
	wire _1158_;
	wire _1159_;
	wire _1160_;
	wire _1161_;
	wire _1162_;
	wire _1163_;
	wire _1164_;
	wire _1165_;
	wire _1166_;
	wire _1167_;
	wire _1168_;
	wire _1169_;
	wire _1170_;
	wire _1171_;
	wire _1172_;
	wire _1173_;
	wire _1174_;
	wire _1175_;
	wire _1176_;
	wire _1177_;
	wire _1178_;
	wire _1179_;
	wire _1180_;
	wire _1181_;
	wire _1182_;
	wire _1183_;
	wire _1184_;
	wire _1185_;
	wire _1186_;
	wire _1187_;
	wire _1188_;
	wire _1189_;
	wire _1190_;
	wire _1191_;
	wire _1192_;
	wire _1193_;
	wire _1194_;
	wire _1195_;
	wire _1196_;
	wire _1197_;
	wire _1198_;
	wire _1199_;
	wire _1200_;
	wire _1201_;
	wire _1202_;
	wire _1203_;
	wire _1204_;
	wire _1205_;
	wire _1206_;
	wire _1207_;
	wire _1208_;
	wire _1209_;
	wire _1210_;
	wire _1211_;
	wire _1212_;
	wire _1213_;
	wire _1214_;
	wire _1215_;
	wire _1216_;
	wire _1217_;
	wire _1218_;
	wire _1219_;
	wire _1220_;
	wire _1221_;
	wire _1222_;
	wire _1223_;
	wire _1224_;
	wire _1225_;
	wire _1226_;
	wire _1227_;
	wire _1228_;
	wire _1229_;
	wire _1230_;
	wire _1231_;
	wire _1232_;
	wire _1233_;
	wire _1234_;
	wire _1235_;
	wire _1236_;
	wire _1237_;
	wire _1238_;
	wire _1239_;
	wire _1240_;
	wire _1241_;
	wire _1242_;
	wire _1243_;
	wire _1244_;
	wire _1245_;
	wire _1246_;
	wire _1247_;
	wire _1248_;
	wire _1249_;
	wire _1250_;
	wire _1251_;
	wire _1252_;
	wire _1253_;
	wire _1254_;
	wire _1255_;
	wire _1256_;
	wire _1257_;
	wire _1258_;
	wire _1259_;
	wire _1260_;
	wire _1261_;
	wire _1262_;
	wire _1263_;
	wire _1264_;
	wire _1265_;
	wire _1266_;
	wire _1267_;
	wire _1268_;
	wire _1269_;
	wire _1270_;
	wire _1271_;
	wire _1272_;
	wire _1273_;
	wire _1274_;
	wire _1275_;
	wire _1276_;
	wire _1277_;
	wire _1278_;
	wire _1279_;
	wire _1280_;
	wire _1281_;
	wire _1282_;
	wire _1283_;
	wire _1284_;
	wire _1285_;
	wire _1286_;
	wire _1287_;
	wire _1288_;
	wire _1289_;
	wire _1290_;
	wire _1291_;
	wire _1292_;
	wire _1293_;
	wire _1294_;
	wire _1295_;
	wire _1296_;
	wire _1297_;
	wire _1298_;
	wire _1299_;
	wire _1300_;
	wire _1301_;
	wire _1302_;
	wire _1303_;
	wire _1304_;
	wire _1305_;
	wire _1306_;
	wire _1307_;
	wire _1308_;
	wire _1309_;
	wire _1310_;
	wire _1311_;
	wire _1312_;
	wire _1313_;
	wire _1314_;
	wire _1315_;
	wire _1316_;
	wire _1317_;
	wire _1318_;
	wire _1319_;
	wire _1320_;
	wire _1321_;
	wire _1322_;
	wire _1323_;
	wire _1324_;
	wire _1325_;
	wire _1326_;
	wire _1327_;
	wire _1328_;
	wire _1329_;
	wire _1330_;
	wire _1331_;
	wire _1332_;
	wire _1333_;
	wire _1334_;
	wire _1335_;
	wire _1336_;
	wire _1337_;
	wire _1338_;
	wire _1339_;
	wire _1340_;
	wire _1341_;
	wire _1342_;
	wire _1343_;
	wire _1344_;
	wire _1345_;
	wire _1346_;
	wire _1347_;
	wire _1348_;
	wire _1349_;
	wire _1350_;
	wire _1351_;
	wire _1352_;
	wire _1353_;
	wire _1354_;
	wire _1355_;
	wire _1356_;
	wire _1357_;
	wire _1358_;
	wire _1359_;
	wire _1360_;
	wire _1361_;
	wire _1362_;
	wire _1363_;
	wire _1364_;
	wire _1365_;
	wire _1366_;
	wire _1367_;
	wire _1368_;
	wire _1369_;
	wire _1370_;
	wire _1371_;
	wire _1372_;
	wire _1373_;
	wire _1374_;
	wire _1375_;
	wire _1376_;
	wire _1377_;
	wire _1378_;
	wire _1379_;
	wire _1380_;
	wire _1381_;
	wire _1382_;
	wire _1383_;
	wire _1384_;
	wire _1385_;
	wire _1386_;
	wire _1387_;
	wire _1388_;
	wire _1389_;
	wire _1390_;
	wire _1391_;
	wire _1392_;
	wire _1393_;
	wire _1394_;
	wire _1395_;
	wire _1396_;
	wire _1397_;
	wire _1398_;
	wire _1399_;
	wire _1400_;
	wire _1401_;
	wire _1402_;
	wire _1403_;
	wire _1404_;
	wire _1405_;
	wire _1406_;
	wire _1407_;
	wire _1408_;
	wire _1409_;
	wire _1410_;
	wire _1411_;
	wire _1412_;
	wire _1413_;
	wire _1414_;
	wire _1415_;
	wire [6:0] _1416_;
	input wire [13:0] io_in;
	output wire [13:0] io_out;
	wire \mchip.Done ;
	wire \mchip.Next ;
	wire \mchip.clock ;
	wire \mchip.dut.Compute_done ;
	wire \mchip.dut.DataReg_en ;
	wire \mchip.dut.Done ;
	wire \mchip.dut.Halt ;
	wire \mchip.dut.Init ;
	wire \mchip.dut.InputAddr_en ;
	wire \mchip.dut.Left ;
	wire \mchip.dut.Next ;
	wire \mchip.dut.NextState_en ;
	wire \mchip.dut.Read_en ;
	wire \mchip.dut.StateAddr_ld ;
	wire \mchip.dut.TapeReg_en ;
	wire \mchip.dut.Tape_start ;
	wire \mchip.dut.clock ;
	reg \mchip.dut.data_reg.Q ;
	wire \mchip.dut.data_reg.clear ;
	wire \mchip.dut.data_reg.clock ;
	wire \mchip.dut.data_reg.en ;
	wire \mchip.dut.data_reg_out ;
	wire [4:0] \mchip.dut.demux.I ;
	wire [4:0] \mchip.dut.demux.Y0 ;
	wire [4:0] \mchip.dut.demux.Y1 ;
	wire [4:0] \mchip.dut.demux.Y2 ;
	wire [4:0] \mchip.dut.demux.Y3 ;
	wire [1:0] \mchip.dut.direction_in ;
	wire [1:0] \mchip.dut.direction_out ;
	wire [6:0] \mchip.dut.direction_reg.D ;
	wire [6:0] \mchip.dut.direction_reg.Q ;
	wire \mchip.dut.direction_reg.clear ;
	wire \mchip.dut.direction_reg.clock ;
	wire [10:0] \mchip.dut.display_out ;
	reg [10:0] \mchip.dut.display_reg.Q ;
	wire \mchip.dut.display_reg.clear ;
	wire \mchip.dut.display_reg.clock ;
	wire \mchip.dut.fsm.DataReg_en ;
	wire \mchip.dut.fsm.Done ;
	wire \mchip.dut.fsm.Halt ;
	wire \mchip.dut.fsm.Init ;
	wire \mchip.dut.fsm.InputAddr_en ;
	wire \mchip.dut.fsm.Left ;
	wire \mchip.dut.fsm.Next ;
	wire \mchip.dut.fsm.NextState_en ;
	wire \mchip.dut.fsm.Read_en ;
	wire \mchip.dut.fsm.StateAddr_ld ;
	wire \mchip.dut.fsm.TapeReg_en ;
	wire \mchip.dut.fsm.Tape_start ;
	wire \mchip.dut.fsm.clock ;
	wire [14:0] \mchip.dut.fsm.currState ;
	wire \mchip.dut.fsm.reset ;
	reg [6:0] \mchip.dut.input_addr.Q ;
	wire \mchip.dut.input_addr.clear ;
	wire \mchip.dut.input_addr.clock ;
	wire \mchip.dut.input_addr.en ;
	wire \mchip.dut.input_addr.load ;
	wire \mchip.dut.input_addr.up ;
	wire [6:0] \mchip.dut.input_addr_out ;
	wire [6:0] \mchip.dut.input_data ;
	reg [4:0] \mchip.dut.memory.M[0] ;
	reg [4:0] \mchip.dut.memory.M[100] ;
	reg [4:0] \mchip.dut.memory.M[101] ;
	reg [4:0] \mchip.dut.memory.M[102] ;
	reg [4:0] \mchip.dut.memory.M[103] ;
	reg [4:0] \mchip.dut.memory.M[104] ;
	reg [4:0] \mchip.dut.memory.M[105] ;
	reg [4:0] \mchip.dut.memory.M[106] ;
	reg [4:0] \mchip.dut.memory.M[107] ;
	reg [4:0] \mchip.dut.memory.M[108] ;
	reg [4:0] \mchip.dut.memory.M[109] ;
	reg [4:0] \mchip.dut.memory.M[10] ;
	reg [4:0] \mchip.dut.memory.M[110] ;
	reg [4:0] \mchip.dut.memory.M[111] ;
	reg [4:0] \mchip.dut.memory.M[112] ;
	reg [4:0] \mchip.dut.memory.M[113] ;
	reg [4:0] \mchip.dut.memory.M[114] ;
	reg [4:0] \mchip.dut.memory.M[115] ;
	reg [4:0] \mchip.dut.memory.M[116] ;
	reg [4:0] \mchip.dut.memory.M[117] ;
	reg [4:0] \mchip.dut.memory.M[118] ;
	reg [4:0] \mchip.dut.memory.M[119] ;
	reg [4:0] \mchip.dut.memory.M[11] ;
	reg [4:0] \mchip.dut.memory.M[120] ;
	reg [4:0] \mchip.dut.memory.M[121] ;
	reg [4:0] \mchip.dut.memory.M[122] ;
	reg [4:0] \mchip.dut.memory.M[123] ;
	reg [4:0] \mchip.dut.memory.M[124] ;
	reg [4:0] \mchip.dut.memory.M[125] ;
	reg [4:0] \mchip.dut.memory.M[126] ;
	reg [4:0] \mchip.dut.memory.M[127] ;
	reg [4:0] \mchip.dut.memory.M[12] ;
	reg [4:0] \mchip.dut.memory.M[13] ;
	reg [4:0] \mchip.dut.memory.M[14] ;
	reg [4:0] \mchip.dut.memory.M[15] ;
	reg [4:0] \mchip.dut.memory.M[16] ;
	reg [4:0] \mchip.dut.memory.M[17] ;
	reg [4:0] \mchip.dut.memory.M[18] ;
	reg [4:0] \mchip.dut.memory.M[19] ;
	reg [4:0] \mchip.dut.memory.M[1] ;
	reg [4:0] \mchip.dut.memory.M[20] ;
	reg [4:0] \mchip.dut.memory.M[21] ;
	reg [4:0] \mchip.dut.memory.M[22] ;
	reg [4:0] \mchip.dut.memory.M[23] ;
	reg [4:0] \mchip.dut.memory.M[24] ;
	reg [4:0] \mchip.dut.memory.M[25] ;
	reg [4:0] \mchip.dut.memory.M[26] ;
	reg [4:0] \mchip.dut.memory.M[27] ;
	reg [4:0] \mchip.dut.memory.M[28] ;
	reg [4:0] \mchip.dut.memory.M[29] ;
	reg [4:0] \mchip.dut.memory.M[2] ;
	reg [4:0] \mchip.dut.memory.M[30] ;
	reg [4:0] \mchip.dut.memory.M[31] ;
	reg [4:0] \mchip.dut.memory.M[32] ;
	reg [4:0] \mchip.dut.memory.M[33] ;
	reg [4:0] \mchip.dut.memory.M[34] ;
	reg [4:0] \mchip.dut.memory.M[35] ;
	reg [4:0] \mchip.dut.memory.M[36] ;
	reg [4:0] \mchip.dut.memory.M[37] ;
	reg [4:0] \mchip.dut.memory.M[38] ;
	reg [4:0] \mchip.dut.memory.M[39] ;
	reg [4:0] \mchip.dut.memory.M[3] ;
	reg [4:0] \mchip.dut.memory.M[40] ;
	reg [4:0] \mchip.dut.memory.M[41] ;
	reg [4:0] \mchip.dut.memory.M[42] ;
	reg [4:0] \mchip.dut.memory.M[43] ;
	reg [4:0] \mchip.dut.memory.M[44] ;
	reg [4:0] \mchip.dut.memory.M[45] ;
	reg [4:0] \mchip.dut.memory.M[46] ;
	reg [4:0] \mchip.dut.memory.M[47] ;
	reg [4:0] \mchip.dut.memory.M[48] ;
	reg [4:0] \mchip.dut.memory.M[49] ;
	reg [4:0] \mchip.dut.memory.M[4] ;
	reg [4:0] \mchip.dut.memory.M[50] ;
	reg [4:0] \mchip.dut.memory.M[51] ;
	reg [4:0] \mchip.dut.memory.M[52] ;
	reg [4:0] \mchip.dut.memory.M[53] ;
	reg [4:0] \mchip.dut.memory.M[54] ;
	reg [4:0] \mchip.dut.memory.M[55] ;
	reg [4:0] \mchip.dut.memory.M[56] ;
	reg [4:0] \mchip.dut.memory.M[57] ;
	reg [4:0] \mchip.dut.memory.M[58] ;
	reg [4:0] \mchip.dut.memory.M[59] ;
	reg [4:0] \mchip.dut.memory.M[5] ;
	reg [4:0] \mchip.dut.memory.M[60] ;
	reg [4:0] \mchip.dut.memory.M[61] ;
	reg [4:0] \mchip.dut.memory.M[62] ;
	reg [4:0] \mchip.dut.memory.M[63] ;
	reg [4:0] \mchip.dut.memory.M[64] ;
	reg [4:0] \mchip.dut.memory.M[65] ;
	reg [4:0] \mchip.dut.memory.M[66] ;
	reg [4:0] \mchip.dut.memory.M[67] ;
	reg [4:0] \mchip.dut.memory.M[68] ;
	reg [4:0] \mchip.dut.memory.M[69] ;
	reg [4:0] \mchip.dut.memory.M[6] ;
	reg [4:0] \mchip.dut.memory.M[70] ;
	reg [4:0] \mchip.dut.memory.M[71] ;
	reg [4:0] \mchip.dut.memory.M[72] ;
	reg [4:0] \mchip.dut.memory.M[73] ;
	reg [4:0] \mchip.dut.memory.M[74] ;
	reg [4:0] \mchip.dut.memory.M[75] ;
	reg [4:0] \mchip.dut.memory.M[76] ;
	reg [4:0] \mchip.dut.memory.M[77] ;
	reg [4:0] \mchip.dut.memory.M[78] ;
	reg [4:0] \mchip.dut.memory.M[79] ;
	reg [4:0] \mchip.dut.memory.M[7] ;
	reg [4:0] \mchip.dut.memory.M[80] ;
	reg [4:0] \mchip.dut.memory.M[81] ;
	reg [4:0] \mchip.dut.memory.M[82] ;
	reg [4:0] \mchip.dut.memory.M[83] ;
	reg [4:0] \mchip.dut.memory.M[84] ;
	reg [4:0] \mchip.dut.memory.M[85] ;
	reg [4:0] \mchip.dut.memory.M[86] ;
	reg [4:0] \mchip.dut.memory.M[87] ;
	reg [4:0] \mchip.dut.memory.M[88] ;
	reg [4:0] \mchip.dut.memory.M[89] ;
	reg [4:0] \mchip.dut.memory.M[8] ;
	reg [4:0] \mchip.dut.memory.M[90] ;
	reg [4:0] \mchip.dut.memory.M[91] ;
	reg [4:0] \mchip.dut.memory.M[92] ;
	reg [4:0] \mchip.dut.memory.M[93] ;
	reg [4:0] \mchip.dut.memory.M[94] ;
	reg [4:0] \mchip.dut.memory.M[95] ;
	reg [4:0] \mchip.dut.memory.M[96] ;
	reg [4:0] \mchip.dut.memory.M[97] ;
	reg [4:0] \mchip.dut.memory.M[98] ;
	reg [4:0] \mchip.dut.memory.M[99] ;
	reg [4:0] \mchip.dut.memory.M[9] ;
	wire \mchip.dut.memory.clock ;
	wire [4:0] \mchip.dut.memory.data_in ;
	wire [4:0] \mchip.dut.memory.data_out ;
	wire \mchip.dut.memory.re ;
	wire [6:0] \mchip.dut.mux_display.I0 ;
	wire [6:0] \mchip.dut.mux_display.I1 ;
	wire \mchip.dut.mux_display.S ;
	wire [6:0] \mchip.dut.mux_display.Y ;
	wire [4:0] \mchip.dut.mux_input_calculate.I0 ;
	wire [4:0] \mchip.dut.mux_input_calculate.I1 ;
	wire [4:0] \mchip.dut.mux_input_calculate.Y ;
	wire [6:0] \mchip.dut.mux_next_state.I0 ;
	wire [6:0] \mchip.dut.mux_next_state.I1 ;
	wire \mchip.dut.mux_next_state.S ;
	wire [6:0] \mchip.dut.mux_next_state.Y ;
	wire \mchip.dut.mux_prev_tape.I0 ;
	wire \mchip.dut.mux_prev_tape.I1 ;
	wire \mchip.dut.mux_prev_tape.Y ;
	wire [6:0] \mchip.dut.mux_state_tape_addr.I0 ;
	wire [6:0] \mchip.dut.mux_state_tape_addr.I1 ;
	wire [6:0] \mchip.dut.mux_state_tape_addr.I3 ;
	wire \mchip.dut.mux_tape_reg.I0 ;
	wire \mchip.dut.mux_tape_reg.I1 ;
	wire \mchip.dut.mux_tape_reg.S ;
	wire \mchip.dut.mux_tape_reg.Y ;
	wire [6:0] \mchip.dut.next_state.D ;
	wire [6:0] \mchip.dut.next_state.Q ;
	wire \mchip.dut.next_state.clear ;
	wire \mchip.dut.next_state.clock ;
	wire \mchip.dut.next_state.en ;
	wire [6:0] \mchip.dut.next_state_in ;
	wire [6:0] \mchip.dut.next_state_out ;
	wire [6:0] \mchip.dut.next_state_prep ;
	wire \mchip.dut.prev_tape_in ;
	wire \mchip.dut.prev_tape_out ;
	wire \mchip.dut.prev_tape_reg.D ;
	wire \mchip.dut.prev_tape_reg.Q ;
	wire \mchip.dut.prev_tape_reg.clear ;
	wire \mchip.dut.prev_tape_reg.clock ;
	wire [4:0] \mchip.dut.read_data ;
	wire \mchip.dut.reset ;
	wire [6:0] \mchip.dut.state_addr.D ;
	reg [6:0] \mchip.dut.state_addr.Q ;
	wire \mchip.dut.state_addr.clear ;
	wire \mchip.dut.state_addr.clock ;
	wire \mchip.dut.state_addr.load ;
	wire \mchip.dut.state_addr.up ;
	wire [6:0] \mchip.dut.state_addr_in ;
	wire [6:0] \mchip.dut.state_addr_out ;
	wire [6:0] \mchip.dut.tape_addr.D ;
	reg [6:0] \mchip.dut.tape_addr.Q ;
	wire \mchip.dut.tape_addr.clear ;
	wire \mchip.dut.tape_addr.clock ;
	wire [6:0] \mchip.dut.tape_addr_init.D ;
	wire [6:0] \mchip.dut.tape_addr_init.Q ;
	wire \mchip.dut.tape_addr_init.clear ;
	wire \mchip.dut.tape_addr_init.clock ;
	wire [6:0] \mchip.dut.tape_addr_min.D ;
	wire [6:0] \mchip.dut.tape_addr_min.Q ;
	wire \mchip.dut.tape_addr_min.clear ;
	wire \mchip.dut.tape_addr_min.clock ;
	wire \mchip.dut.tape_addr_min.en ;
	wire [6:0] \mchip.dut.tape_addr_out ;
	wire \mchip.dut.tape_in ;
	wire [6:0] \mchip.dut.tape_init_addr ;
	wire [6:0] \mchip.dut.tape_min_addr_in ;
	wire [6:0] \mchip.dut.tape_min_addr_out ;
	wire \mchip.dut.tape_reg.D ;
	reg \mchip.dut.tape_reg.Q ;
	wire \mchip.dut.tape_reg.clear ;
	wire \mchip.dut.tape_reg.clock ;
	wire \mchip.dut.tape_reg.en ;
	wire \mchip.dut.tape_reg_in ;
	wire \mchip.dut.tape_reg_out ;
	wire [4:0] \mchip.dut.write_data ;
	wire [6:0] \mchip.input_data ;
	wire [11:0] \mchip.io_in ;
	wire [11:0] \mchip.io_out ;
	wire \mchip.reset ;
	wire \mchip.sync1.async ;
	reg \mchip.sync1.async1 ;
	wire \mchip.sync1.clock ;
	reg \mchip.sync1.sync ;
	wire \mchip.sync2.async ;
	reg \mchip.sync2.async1 ;
	wire \mchip.sync2.clock ;
	reg \mchip.sync2.sync ;
	wire \mchip.sync3.async ;
	reg \mchip.sync3.async1 ;
	wire \mchip.sync3.clock ;
	reg \mchip.sync3.sync ;
	wire \mchip.sync4.async ;
	reg \mchip.sync4.async1 ;
	wire \mchip.sync4.clock ;
	reg \mchip.sync4.sync ;
	wire \mchip.sync5.async ;
	reg \mchip.sync5.async1 ;
	wire \mchip.sync5.clock ;
	reg \mchip.sync5.sync ;
	wire \mchip.sync6.async ;
	reg \mchip.sync6.async1 ;
	wire \mchip.sync6.clock ;
	reg \mchip.sync6.sync ;
	wire \mchip.sync7.async ;
	reg \mchip.sync7.async1 ;
	wire \mchip.sync7.clock ;
	reg \mchip.sync7.sync ;
	wire \mchip.sync8.async ;
	reg \mchip.sync8.async1 ;
	wire \mchip.sync8.clock ;
	reg \mchip.sync8.sync ;
	assign _1416_[0] = ~\mchip.dut.input_addr.Q [0];
	assign _0019_ = \mchip.dut.fsm.currState [9] | \mchip.dut.fsm.currState [0];
	assign _1339_ = ~\mchip.sync1.sync ;
	assign _1340_ = \mchip.dut.tape_reg.Q  ^ \mchip.dut.data_reg.Q ;
	assign _1341_ = _1340_ | _1339_;
	assign _1342_ = \mchip.dut.fsm.currState [5] & ~_1341_;
	assign _1343_ = _1342_ | \mchip.dut.fsm.currState [13];
	assign _1344_ = ~(\mchip.dut.fsm.currState [13] | \mchip.dut.fsm.currState [5]);
	assign _1345_ = _1343_ & ~_1344_;
	assign _0018_ = _1345_ | \mchip.dut.fsm.currState [0];
	assign _1346_ = \mchip.dut.fsm.currState [9] & ~\mchip.dut.direction_reg.Q [1];
	assign _1347_ = ~(_1340_ & \mchip.sync1.sync );
	assign _1348_ = \mchip.dut.fsm.currState [5] & ~_1347_;
	assign _0020_ = _1346_ & ~_1348_;
	assign _1349_ = ~\mchip.dut.fsm.currState [10];
	assign _1350_ = \mchip.sync1.sync  & ~io_in[13];
	assign _1351_ = _1350_ & ~_1349_;
	assign _1352_ = _1350_ & \mchip.dut.fsm.currState [2];
	assign _0006_ = _1352_ | _1351_;
	assign _1353_ = ~\mchip.dut.direction_reg.Q [0];
	assign _1354_ = \mchip.dut.direction_reg.Q [1] | ~\mchip.dut.fsm.currState [9];
	assign _1355_ = _1353_ & ~_1354_;
	assign _1356_ = \mchip.dut.direction_reg.Q [0] & ~_1354_;
	assign _1357_ = _1348_ | _1356_;
	assign _0017_ = _1357_ | _1355_;
	assign _1358_ = ~(\mchip.dut.tape_addr_min.Q [4] ^ \mchip.dut.tape_addr.Q [4]);
	assign _1359_ = \mchip.dut.tape_addr_min.Q [3] ^ \mchip.dut.tape_addr.Q [3];
	assign _1360_ = _1358_ & ~_1359_;
	assign _1361_ = \mchip.dut.tape_addr.Q [2] | ~\mchip.dut.tape_addr_min.Q [2];
	assign _1362_ = \mchip.dut.tape_addr_min.Q [1] | ~\mchip.dut.tape_addr.Q [1];
	assign _1363_ = \mchip.dut.tape_addr_min.Q [2] ^ \mchip.dut.tape_addr.Q [2];
	assign _1364_ = _1362_ & ~_1363_;
	assign _1365_ = _1361_ & ~_1364_;
	assign _1366_ = _1360_ & ~_1365_;
	assign _1367_ = \mchip.dut.tape_addr_min.Q [4] & ~\mchip.dut.tape_addr.Q [4];
	assign _1368_ = \mchip.dut.tape_addr.Q [3] | ~\mchip.dut.tape_addr_min.Q [3];
	assign _1369_ = _1358_ & ~_1368_;
	assign _1370_ = _1369_ | _1367_;
	assign _1371_ = _1370_ | _1366_;
	assign _1372_ = \mchip.dut.tape_addr_min.Q [5] ^ \mchip.dut.tape_addr.Q [5];
	assign _1373_ = \mchip.dut.tape_addr_min.Q [6] ^ \mchip.dut.tape_addr.Q [6];
	assign _1374_ = _1373_ | _1372_;
	assign _1375_ = _1371_ & ~_1374_;
	assign _1376_ = \mchip.dut.tape_addr_min.Q [5] & ~\mchip.dut.tape_addr.Q [5];
	assign _1377_ = _1376_ & ~_1373_;
	assign _1378_ = \mchip.dut.tape_addr_min.Q [6] & ~\mchip.dut.tape_addr.Q [6];
	assign _1379_ = _1378_ | _1377_;
	assign _1380_ = _1379_ | _1375_;
	assign _1381_ = \mchip.dut.tape_addr_min.Q [1] ^ \mchip.dut.tape_addr.Q [1];
	assign _1382_ = _1381_ | _1363_;
	assign _1383_ = _1360_ & ~_1382_;
	assign _1384_ = ~\mchip.dut.tape_addr.Q [0];
	assign _1385_ = _1374_ | _1384_;
	assign _1386_ = _1383_ & ~_1385_;
	assign _1387_ = _1380_ & ~_1386_;
	assign _1388_ = ~(\mchip.dut.tape_addr.Q [4] & \mchip.dut.tape_addr.Q [5]);
	assign _1389_ = \mchip.dut.tape_addr.Q [0] & \mchip.dut.tape_addr.Q [1];
	assign _1390_ = ~(\mchip.dut.tape_addr.Q [2] & \mchip.dut.tape_addr.Q [3]);
	assign _1391_ = _1389_ & ~_1390_;
	assign _1392_ = _1388_ | ~_1391_;
	assign _1393_ = \mchip.dut.tape_addr.Q [6] & ~_1392_;
	assign _1394_ = _1388_ | ~\mchip.dut.tape_addr.Q [6];
	assign _1395_ = _1391_ & ~_1394_;
	assign _1396_ = _1395_ | _1393_;
	assign _1397_ = _1396_ | _1387_;
	assign _1398_ = _1397_ | io_in[13];
	assign _1399_ = \mchip.dut.fsm.currState [11] & ~_1398_;
	assign _1400_ = ~\mchip.dut.input_addr.Q [6];
	assign _1401_ = ~(\mchip.dut.input_addr.Q [4] & \mchip.dut.input_addr.Q [5]);
	assign _1402_ = _1401_ | _1400_;
	assign _1403_ = \mchip.dut.input_addr.Q [1] & \mchip.dut.input_addr.Q [0];
	assign _1404_ = \mchip.dut.input_addr.Q [2] & \mchip.dut.input_addr.Q [3];
	assign _1405_ = ~(_1404_ & _1403_);
	assign _1406_ = _1405_ | _1402_;
	assign _1407_ = ~(_1405_ | _1401_);
	assign _1408_ = _1407_ & ~_1400_;
	assign _1409_ = _1406_ & ~_1408_;
	assign _1410_ = _1409_ | io_in[13];
	assign _1411_ = \mchip.dut.fsm.currState [1] & ~_1410_;
	assign _0013_ = _1411_ | _1399_;
	assign _1412_ = ~(io_in[13] | \mchip.sync1.sync );
	assign _1413_ = _1412_ & ~_1349_;
	assign _1414_ = _1412_ & \mchip.dut.fsm.currState [14];
	assign _1415_ = \mchip.sync2.sync  | io_in[13];
	assign _0177_ = _1415_ | \mchip.sync1.sync ;
	assign _0178_ = \mchip.dut.fsm.currState [6] & ~_0177_;
	assign _0179_ = _0178_ | _1414_;
	assign _0012_ = _0179_ | _1413_;
	assign _0180_ = io_in[13] | ~\mchip.sync2.sync ;
	assign _0181_ = _0180_ | \mchip.sync1.sync ;
	assign _0182_ = \mchip.dut.fsm.currState [4] & ~_0181_;
	assign _0183_ = _1412_ & \mchip.dut.fsm.currState [2];
	assign _0008_ = _0183_ | _0182_;
	assign _0184_ = ~(\mchip.dut.fsm.currState [11] | \mchip.dut.fsm.currState [1]);
	assign _0185_ = ~\mchip.dut.fsm.currState [1];
	assign _0186_ = _1409_ | _0185_;
	assign _0187_ = \mchip.dut.fsm.currState [11] & ~_1397_;
	assign _0188_ = _0186_ & ~_0187_;
	assign \mchip.dut.StateAddr_ld  = ~(_0188_ | _0184_);
	assign _0014_ = \mchip.dut.StateAddr_ld  | \mchip.dut.fsm.currState [0];
	assign _0189_ = io_in[13] | ~_1409_;
	assign _0190_ = \mchip.dut.fsm.currState [1] & ~_0189_;
	assign _0191_ = \mchip.dut.fsm.currState [6] & ~_0181_;
	assign _0007_ = _0191_ | _0190_;
	assign _0192_ = _0187_ | _1343_;
	assign _0193_ = _0186_ & ~_0192_;
	assign _0194_ = ~(\mchip.dut.fsm.currState [3] | \mchip.dut.fsm.currState [11]);
	assign _0195_ = ~(_0194_ & _1344_);
	assign _0196_ = _0185_ & ~_0195_;
	assign _0197_ = _0196_ | _0193_;
	assign _0198_ = \mchip.dut.fsm.currState [3] & ~\mchip.sync1.sync ;
	assign _0199_ = _0198_ | _0187_;
	assign _0200_ = _0186_ & ~_0199_;
	assign _0201_ = _0200_ | _0196_;
	assign _0202_ = _0201_ & _0197_;
	assign _0203_ = _0202_ | \mchip.dut.fsm.currState [0];
	assign _0023_ = _0203_ | ~_0197_;
	assign _0204_ = ~\mchip.dut.fsm.currState [5];
	assign _0205_ = _1412_ & ~_0204_;
	assign _0206_ = \mchip.dut.fsm.currState [9] & ~io_in[13];
	assign _0011_ = _0206_ | _0205_;
	assign _0207_ = \mchip.dut.fsm.currState [4] & ~_0177_;
	assign _0208_ = ~(\mchip.dut.fsm.currState [12] | \mchip.dut.fsm.currState [8]);
	assign _0209_ = _1412_ & ~_0208_;
	assign _0010_ = _0209_ | _0207_;
	assign _0210_ = ~(_0201_ | _0197_);
	assign _0211_ = _0210_ | ~_1345_;
	assign _0022_ = _0211_ | _0197_;
	assign _0212_ = \mchip.dut.fsm.currState [13] | \mchip.dut.fsm.currState [9];
	assign _0213_ = _0212_ | _1342_;
	assign _0214_ = _0204_ & ~_0212_;
	assign _0215_ = _0213_ & ~_0214_;
	assign _0016_ = _0215_ | \mchip.dut.StateAddr_ld ;
	assign _0216_ = ~\mchip.dut.fsm.currState [3];
	assign _0217_ = _1350_ & ~_0216_;
	assign _0218_ = \mchip.dut.fsm.currState [13] & ~io_in[13];
	assign _0219_ = _1340_ | io_in[13];
	assign _0220_ = _0219_ | _1339_;
	assign _0221_ = \mchip.dut.fsm.currState [5] & ~_0220_;
	assign _0222_ = _0221_ | _0218_;
	assign _0009_ = _0222_ | _0217_;
	assign _0223_ = \mchip.dut.direction_reg.Q [1] | \mchip.sync1.sync ;
	assign _0224_ = _0223_ | _0216_;
	assign _0225_ = _1353_ & ~_0224_;
	assign _0226_ = \mchip.dut.direction_reg.Q [0] & ~_0224_;
	assign _0227_ = \mchip.dut.fsm.currState [2] & \mchip.sync1.sync ;
	assign _0228_ = _0227_ | _0226_;
	assign _0015_ = _0228_ | _0225_;
	assign _0229_ = _0210_ | ~\mchip.dut.fsm.currState [9];
	assign _0230_ = _0201_ ^ _0197_;
	assign _0021_ = _0230_ | _0229_;
	assign _0231_ = _1412_ & \mchip.dut.fsm.currState [0];
	assign _0005_ = _0231_ | io_in[13];
	assign _0232_ = ~\mchip.dut.memory.M[127] [0];
	assign _0233_ = ~\mchip.dut.memory.M[126] [0];
	assign _0234_ = ~(\mchip.dut.fsm.currState [4] | \mchip.dut.fsm.currState [6]);
	assign _0235_ = \mchip.sync1.sync  & ~_0234_;
	assign _0236_ = _0235_ | \mchip.dut.fsm.currState [1];
	assign _0237_ = _1397_ | \mchip.dut.direction_reg.Q [0];
	assign _0238_ = \mchip.dut.fsm.currState [11] & ~_0237_;
	assign _0239_ = _0238_ | _1348_;
	assign _0240_ = _0239_ | _0236_;
	assign _0241_ = ~(_0234_ & _0185_);
	assign _0242_ = \mchip.dut.fsm.currState [11] | \mchip.dut.fsm.currState [5];
	assign _0243_ = _0242_ | _0241_;
	assign _0244_ = _1349_ & ~_0243_;
	assign _0245_ = _0240_ & ~_0244_;
	assign _0246_ = (_0245_ ? \mchip.dut.input_addr.Q [0] : _1384_);
	assign _0247_ = \mchip.dut.direction_reg.Q [0] & ~_1397_;
	assign _0248_ = ~(_0247_ & \mchip.dut.fsm.currState [11]);
	assign _0249_ = _1409_ & ~_0185_;
	assign _0250_ = _0249_ | _0235_;
	assign _0251_ = _0250_ | ~_0248_;
	assign _0252_ = _0251_ & ~_0244_;
	assign _0253_ = (_0245_ ? \mchip.dut.tape_addr.Q [0] : \mchip.dut.state_addr.Q [0]);
	assign _0254_ = (_0252_ ? _0246_ : _0253_);
	assign _0255_ = (_0254_ ? _0232_ : _0233_);
	assign _0256_ = \mchip.dut.tape_addr.Q [0] ^ \mchip.dut.tape_addr.Q [1];
	assign _0257_ = (_0245_ ? \mchip.dut.input_addr.Q [1] : _0256_);
	assign _0258_ = (_0245_ ? \mchip.dut.tape_addr.Q [1] : \mchip.dut.state_addr.Q [1]);
	assign _0259_ = (_0252_ ? _0257_ : _0258_);
	assign _0260_ = ~\mchip.dut.memory.M[125] [0];
	assign _0261_ = ~\mchip.dut.memory.M[124] [0];
	assign _0262_ = (_0254_ ? _0260_ : _0261_);
	assign _0263_ = (_0259_ ? _0255_ : _0262_);
	assign _0264_ = ~\mchip.dut.tape_addr.Q [2];
	assign _0265_ = _1389_ ^ _0264_;
	assign _0266_ = (_0245_ ? \mchip.dut.input_addr.Q [2] : _0265_);
	assign _0267_ = (_0245_ ? \mchip.dut.tape_addr.Q [2] : \mchip.dut.state_addr.Q [2]);
	assign _0268_ = (_0252_ ? _0266_ : _0267_);
	assign _0269_ = ~\mchip.dut.memory.M[123] [0];
	assign _0270_ = ~\mchip.dut.memory.M[122] [0];
	assign _0271_ = (_0254_ ? _0269_ : _0270_);
	assign _0272_ = ~\mchip.dut.memory.M[121] [0];
	assign _0273_ = ~\mchip.dut.memory.M[120] [0];
	assign _0274_ = (_0254_ ? _0272_ : _0273_);
	assign _0275_ = (_0259_ ? _0271_ : _0274_);
	assign _0276_ = (_0268_ ? _0263_ : _0275_);
	assign _0277_ = ~\mchip.dut.tape_addr.Q [3];
	assign _0278_ = _0264_ & ~_1389_;
	assign _0279_ = _0278_ ^ _0277_;
	assign _0280_ = (_0245_ ? \mchip.dut.input_addr.Q [3] : _0279_);
	assign _0281_ = (_0245_ ? \mchip.dut.tape_addr.Q [3] : \mchip.dut.state_addr.Q [3]);
	assign _0282_ = (_0252_ ? _0280_ : _0281_);
	assign _0283_ = ~\mchip.dut.memory.M[119] [0];
	assign _0284_ = ~\mchip.dut.memory.M[118] [0];
	assign _0285_ = (_0254_ ? _0283_ : _0284_);
	assign _0286_ = ~\mchip.dut.memory.M[117] [0];
	assign _0287_ = ~\mchip.dut.memory.M[116] [0];
	assign _0288_ = (_0254_ ? _0286_ : _0287_);
	assign _0289_ = (_0259_ ? _0285_ : _0288_);
	assign _0290_ = ~\mchip.dut.memory.M[115] [0];
	assign _0291_ = ~\mchip.dut.memory.M[114] [0];
	assign _0292_ = (_0254_ ? _0290_ : _0291_);
	assign _0293_ = ~\mchip.dut.memory.M[113] [0];
	assign _0294_ = ~\mchip.dut.memory.M[112] [0];
	assign _0295_ = (_0254_ ? _0293_ : _0294_);
	assign _0296_ = (_0259_ ? _0292_ : _0295_);
	assign _0297_ = (_0268_ ? _0289_ : _0296_);
	assign _0298_ = (_0282_ ? _0276_ : _0297_);
	assign _0299_ = \mchip.dut.tape_addr.Q [2] | ~\mchip.dut.tape_addr.Q [3];
	assign _0300_ = _1389_ & ~_0299_;
	assign _0301_ = _1390_ & ~_0300_;
	assign _0302_ = _0301_ ^ \mchip.dut.tape_addr.Q [4];
	assign _0303_ = (_0245_ ? \mchip.dut.input_addr.Q [4] : _0302_);
	assign _0304_ = (_0245_ ? \mchip.dut.tape_addr.Q [4] : \mchip.dut.state_addr.Q [4]);
	assign _0305_ = (_0252_ ? _0303_ : _0304_);
	assign _0306_ = ~\mchip.dut.memory.M[111] [0];
	assign _0307_ = ~\mchip.dut.memory.M[110] [0];
	assign _0308_ = (_0254_ ? _0306_ : _0307_);
	assign _0309_ = ~\mchip.dut.memory.M[109] [0];
	assign _0310_ = ~\mchip.dut.memory.M[108] [0];
	assign _0311_ = (_0254_ ? _0309_ : _0310_);
	assign _0312_ = (_0259_ ? _0308_ : _0311_);
	assign _0313_ = ~\mchip.dut.memory.M[107] [0];
	assign _0314_ = ~\mchip.dut.memory.M[106] [0];
	assign _0315_ = (_0254_ ? _0313_ : _0314_);
	assign _0316_ = ~\mchip.dut.memory.M[105] [0];
	assign _0317_ = ~\mchip.dut.memory.M[104] [0];
	assign _0318_ = (_0254_ ? _0316_ : _0317_);
	assign _0319_ = (_0259_ ? _0315_ : _0318_);
	assign _0320_ = (_0268_ ? _0312_ : _0319_);
	assign _0321_ = ~\mchip.dut.memory.M[103] [0];
	assign _0322_ = ~\mchip.dut.memory.M[102] [0];
	assign _0323_ = (_0254_ ? _0321_ : _0322_);
	assign _0324_ = ~\mchip.dut.memory.M[101] [0];
	assign _0325_ = ~\mchip.dut.memory.M[100] [0];
	assign _0326_ = (_0254_ ? _0324_ : _0325_);
	assign _0327_ = (_0259_ ? _0323_ : _0326_);
	assign _0328_ = ~\mchip.dut.memory.M[99] [0];
	assign _0329_ = ~\mchip.dut.memory.M[98] [0];
	assign _0330_ = (_0254_ ? _0328_ : _0329_);
	assign _0331_ = ~\mchip.dut.memory.M[97] [0];
	assign _0332_ = ~\mchip.dut.memory.M[96] [0];
	assign _0333_ = (_0254_ ? _0331_ : _0332_);
	assign _0334_ = (_0259_ ? _0330_ : _0333_);
	assign _0335_ = (_0268_ ? _0327_ : _0334_);
	assign _0336_ = (_0282_ ? _0320_ : _0335_);
	assign _0337_ = (_0305_ ? _0298_ : _0336_);
	assign _0338_ = _0301_ & ~\mchip.dut.tape_addr.Q [4];
	assign _0339_ = _0338_ ^ \mchip.dut.tape_addr.Q [5];
	assign _0340_ = (_0245_ ? \mchip.dut.input_addr.Q [5] : _0339_);
	assign _0341_ = (_0245_ ? \mchip.dut.tape_addr.Q [5] : \mchip.dut.state_addr.Q [5]);
	assign _0342_ = (_0252_ ? _0340_ : _0341_);
	assign _0343_ = ~\mchip.dut.memory.M[95] [0];
	assign _0344_ = ~\mchip.dut.memory.M[94] [0];
	assign _0345_ = (_0254_ ? _0343_ : _0344_);
	assign _0346_ = ~\mchip.dut.memory.M[93] [0];
	assign _0347_ = ~\mchip.dut.memory.M[92] [0];
	assign _0348_ = (_0254_ ? _0346_ : _0347_);
	assign _0349_ = (_0259_ ? _0345_ : _0348_);
	assign _0350_ = ~\mchip.dut.memory.M[91] [0];
	assign _0351_ = ~\mchip.dut.memory.M[90] [0];
	assign _0352_ = (_0254_ ? _0350_ : _0351_);
	assign _0353_ = ~\mchip.dut.memory.M[89] [0];
	assign _0354_ = ~\mchip.dut.memory.M[88] [0];
	assign _0355_ = (_0254_ ? _0353_ : _0354_);
	assign _0356_ = (_0259_ ? _0352_ : _0355_);
	assign _0357_ = (_0268_ ? _0349_ : _0356_);
	assign _0358_ = ~\mchip.dut.memory.M[87] [0];
	assign _0359_ = ~\mchip.dut.memory.M[86] [0];
	assign _0360_ = (_0254_ ? _0358_ : _0359_);
	assign _0361_ = ~\mchip.dut.memory.M[85] [0];
	assign _0362_ = ~\mchip.dut.memory.M[84] [0];
	assign _0363_ = (_0254_ ? _0361_ : _0362_);
	assign _0364_ = (_0259_ ? _0360_ : _0363_);
	assign _0365_ = ~\mchip.dut.memory.M[83] [0];
	assign _0366_ = ~\mchip.dut.memory.M[82] [0];
	assign _0367_ = (_0254_ ? _0365_ : _0366_);
	assign _0368_ = ~\mchip.dut.memory.M[81] [0];
	assign _0369_ = ~\mchip.dut.memory.M[80] [0];
	assign _0370_ = (_0254_ ? _0368_ : _0369_);
	assign _0371_ = (_0259_ ? _0367_ : _0370_);
	assign _0372_ = (_0268_ ? _0364_ : _0371_);
	assign _0373_ = (_0282_ ? _0357_ : _0372_);
	assign _0374_ = ~\mchip.dut.memory.M[79] [0];
	assign _0375_ = ~\mchip.dut.memory.M[78] [0];
	assign _0376_ = (_0254_ ? _0374_ : _0375_);
	assign _0377_ = ~\mchip.dut.memory.M[77] [0];
	assign _0378_ = ~\mchip.dut.memory.M[76] [0];
	assign _0379_ = (_0254_ ? _0377_ : _0378_);
	assign _0380_ = (_0259_ ? _0376_ : _0379_);
	assign _0381_ = ~\mchip.dut.memory.M[75] [0];
	assign _0382_ = ~\mchip.dut.memory.M[74] [0];
	assign _0383_ = (_0254_ ? _0381_ : _0382_);
	assign _0384_ = ~\mchip.dut.memory.M[73] [0];
	assign _0385_ = ~\mchip.dut.memory.M[72] [0];
	assign _0386_ = (_0254_ ? _0384_ : _0385_);
	assign _0387_ = (_0259_ ? _0383_ : _0386_);
	assign _0388_ = (_0268_ ? _0380_ : _0387_);
	assign _0389_ = ~\mchip.dut.memory.M[71] [0];
	assign _0390_ = ~\mchip.dut.memory.M[70] [0];
	assign _0391_ = (_0254_ ? _0389_ : _0390_);
	assign _0392_ = ~\mchip.dut.memory.M[69] [0];
	assign _0393_ = ~\mchip.dut.memory.M[68] [0];
	assign _0394_ = (_0254_ ? _0392_ : _0393_);
	assign _0395_ = (_0259_ ? _0391_ : _0394_);
	assign _0396_ = ~\mchip.dut.memory.M[67] [0];
	assign _0397_ = ~\mchip.dut.memory.M[66] [0];
	assign _0398_ = (_0254_ ? _0396_ : _0397_);
	assign _0399_ = ~\mchip.dut.memory.M[65] [0];
	assign _0400_ = ~\mchip.dut.memory.M[64] [0];
	assign _0401_ = (_0254_ ? _0399_ : _0400_);
	assign _0402_ = (_0259_ ? _0398_ : _0401_);
	assign _0403_ = (_0268_ ? _0395_ : _0402_);
	assign _0404_ = (_0282_ ? _0388_ : _0403_);
	assign _0405_ = (_0305_ ? _0373_ : _0404_);
	assign _0406_ = (_0342_ ? _0337_ : _0405_);
	assign _0407_ = \mchip.dut.tape_addr.Q [4] | \mchip.dut.tape_addr.Q [5];
	assign _0408_ = _0301_ & ~_0407_;
	assign _0409_ = _0408_ ^ \mchip.dut.tape_addr.Q [6];
	assign _0410_ = (_0245_ ? \mchip.dut.input_addr.Q [6] : _0409_);
	assign _0411_ = (_0245_ ? \mchip.dut.tape_addr.Q [6] : \mchip.dut.state_addr.Q [6]);
	assign _0412_ = (_0252_ ? _0410_ : _0411_);
	assign _0413_ = ~\mchip.dut.memory.M[63] [0];
	assign _0414_ = ~\mchip.dut.memory.M[62] [0];
	assign _0415_ = (_0254_ ? _0413_ : _0414_);
	assign _0416_ = ~\mchip.dut.memory.M[61] [0];
	assign _0417_ = ~\mchip.dut.memory.M[60] [0];
	assign _0418_ = (_0254_ ? _0416_ : _0417_);
	assign _0419_ = (_0259_ ? _0415_ : _0418_);
	assign _0420_ = ~\mchip.dut.memory.M[59] [0];
	assign _0421_ = ~\mchip.dut.memory.M[58] [0];
	assign _0422_ = (_0254_ ? _0420_ : _0421_);
	assign _0423_ = ~\mchip.dut.memory.M[57] [0];
	assign _0424_ = ~\mchip.dut.memory.M[56] [0];
	assign _0425_ = (_0254_ ? _0423_ : _0424_);
	assign _0426_ = (_0259_ ? _0422_ : _0425_);
	assign _0427_ = (_0268_ ? _0419_ : _0426_);
	assign _0428_ = ~\mchip.dut.memory.M[55] [0];
	assign _0429_ = ~\mchip.dut.memory.M[54] [0];
	assign _0430_ = (_0254_ ? _0428_ : _0429_);
	assign _0431_ = ~\mchip.dut.memory.M[53] [0];
	assign _0432_ = ~\mchip.dut.memory.M[52] [0];
	assign _0433_ = (_0254_ ? _0431_ : _0432_);
	assign _0434_ = (_0259_ ? _0430_ : _0433_);
	assign _0435_ = ~\mchip.dut.memory.M[51] [0];
	assign _0436_ = ~\mchip.dut.memory.M[50] [0];
	assign _0437_ = (_0254_ ? _0435_ : _0436_);
	assign _0438_ = ~\mchip.dut.memory.M[49] [0];
	assign _0439_ = ~\mchip.dut.memory.M[48] [0];
	assign _0440_ = (_0254_ ? _0438_ : _0439_);
	assign _0441_ = (_0259_ ? _0437_ : _0440_);
	assign _0442_ = (_0268_ ? _0434_ : _0441_);
	assign _0443_ = (_0282_ ? _0427_ : _0442_);
	assign _0444_ = ~\mchip.dut.memory.M[47] [0];
	assign _0445_ = ~\mchip.dut.memory.M[46] [0];
	assign _0446_ = (_0254_ ? _0444_ : _0445_);
	assign _0447_ = ~\mchip.dut.memory.M[45] [0];
	assign _0448_ = ~\mchip.dut.memory.M[44] [0];
	assign _0449_ = (_0254_ ? _0447_ : _0448_);
	assign _0450_ = (_0259_ ? _0446_ : _0449_);
	assign _0451_ = ~\mchip.dut.memory.M[43] [0];
	assign _0452_ = ~\mchip.dut.memory.M[42] [0];
	assign _0453_ = (_0254_ ? _0451_ : _0452_);
	assign _0454_ = ~\mchip.dut.memory.M[41] [0];
	assign _0455_ = ~\mchip.dut.memory.M[40] [0];
	assign _0456_ = (_0254_ ? _0454_ : _0455_);
	assign _0457_ = (_0259_ ? _0453_ : _0456_);
	assign _0458_ = (_0268_ ? _0450_ : _0457_);
	assign _0459_ = ~\mchip.dut.memory.M[39] [0];
	assign _0460_ = ~\mchip.dut.memory.M[38] [0];
	assign _0461_ = (_0254_ ? _0459_ : _0460_);
	assign _0462_ = ~\mchip.dut.memory.M[37] [0];
	assign _0463_ = ~\mchip.dut.memory.M[36] [0];
	assign _0464_ = (_0254_ ? _0462_ : _0463_);
	assign _0465_ = (_0259_ ? _0461_ : _0464_);
	assign _0466_ = ~\mchip.dut.memory.M[35] [0];
	assign _0467_ = ~\mchip.dut.memory.M[34] [0];
	assign _0468_ = (_0254_ ? _0466_ : _0467_);
	assign _0469_ = ~\mchip.dut.memory.M[33] [0];
	assign _0470_ = ~\mchip.dut.memory.M[32] [0];
	assign _0471_ = (_0254_ ? _0469_ : _0470_);
	assign _0472_ = (_0259_ ? _0468_ : _0471_);
	assign _0473_ = (_0268_ ? _0465_ : _0472_);
	assign _0474_ = (_0282_ ? _0458_ : _0473_);
	assign _0475_ = (_0305_ ? _0443_ : _0474_);
	assign _0476_ = ~\mchip.dut.memory.M[31] [0];
	assign _0477_ = ~\mchip.dut.memory.M[30] [0];
	assign _0478_ = (_0254_ ? _0476_ : _0477_);
	assign _0479_ = ~\mchip.dut.memory.M[29] [0];
	assign _0480_ = ~\mchip.dut.memory.M[28] [0];
	assign _0481_ = (_0254_ ? _0479_ : _0480_);
	assign _0482_ = (_0259_ ? _0478_ : _0481_);
	assign _0483_ = ~\mchip.dut.memory.M[27] [0];
	assign _0484_ = ~\mchip.dut.memory.M[26] [0];
	assign _0485_ = (_0254_ ? _0483_ : _0484_);
	assign _0486_ = ~\mchip.dut.memory.M[25] [0];
	assign _0487_ = ~\mchip.dut.memory.M[24] [0];
	assign _0488_ = (_0254_ ? _0486_ : _0487_);
	assign _0489_ = (_0259_ ? _0485_ : _0488_);
	assign _0490_ = (_0268_ ? _0482_ : _0489_);
	assign _0491_ = ~\mchip.dut.memory.M[23] [0];
	assign _0492_ = ~\mchip.dut.memory.M[22] [0];
	assign _0493_ = (_0254_ ? _0491_ : _0492_);
	assign _0494_ = ~\mchip.dut.memory.M[21] [0];
	assign _0495_ = ~\mchip.dut.memory.M[20] [0];
	assign _0496_ = (_0254_ ? _0494_ : _0495_);
	assign _0497_ = (_0259_ ? _0493_ : _0496_);
	assign _0498_ = ~\mchip.dut.memory.M[19] [0];
	assign _0499_ = ~\mchip.dut.memory.M[18] [0];
	assign _0500_ = (_0254_ ? _0498_ : _0499_);
	assign _0501_ = ~\mchip.dut.memory.M[17] [0];
	assign _0502_ = ~\mchip.dut.memory.M[16] [0];
	assign _0503_ = (_0254_ ? _0501_ : _0502_);
	assign _0504_ = (_0259_ ? _0500_ : _0503_);
	assign _0505_ = (_0268_ ? _0497_ : _0504_);
	assign _0506_ = (_0282_ ? _0490_ : _0505_);
	assign _0507_ = ~\mchip.dut.memory.M[15] [0];
	assign _0508_ = ~\mchip.dut.memory.M[14] [0];
	assign _0509_ = (_0254_ ? _0507_ : _0508_);
	assign _0510_ = ~\mchip.dut.memory.M[13] [0];
	assign _0511_ = ~\mchip.dut.memory.M[12] [0];
	assign _0512_ = (_0254_ ? _0510_ : _0511_);
	assign _0513_ = (_0259_ ? _0509_ : _0512_);
	assign _0514_ = ~\mchip.dut.memory.M[11] [0];
	assign _0515_ = ~\mchip.dut.memory.M[10] [0];
	assign _0516_ = (_0254_ ? _0514_ : _0515_);
	assign _0517_ = ~\mchip.dut.memory.M[9] [0];
	assign _0518_ = ~\mchip.dut.memory.M[8] [0];
	assign _0519_ = (_0254_ ? _0517_ : _0518_);
	assign _0520_ = (_0259_ ? _0516_ : _0519_);
	assign _0521_ = (_0268_ ? _0513_ : _0520_);
	assign _0522_ = ~\mchip.dut.memory.M[7] [0];
	assign _0523_ = ~\mchip.dut.memory.M[6] [0];
	assign _0524_ = (_0254_ ? _0522_ : _0523_);
	assign _0525_ = ~\mchip.dut.memory.M[5] [0];
	assign _0526_ = ~\mchip.dut.memory.M[4] [0];
	assign _0527_ = (_0254_ ? _0525_ : _0526_);
	assign _0528_ = (_0259_ ? _0524_ : _0527_);
	assign _0529_ = ~\mchip.dut.memory.M[3] [0];
	assign _0530_ = ~\mchip.dut.memory.M[2] [0];
	assign _0531_ = (_0254_ ? _0529_ : _0530_);
	assign _0532_ = ~\mchip.dut.memory.M[1] [0];
	assign _0533_ = ~\mchip.dut.memory.M[0] [0];
	assign _0534_ = (_0254_ ? _0532_ : _0533_);
	assign _0535_ = (_0259_ ? _0531_ : _0534_);
	assign _0536_ = (_0268_ ? _0528_ : _0535_);
	assign _0537_ = (_0282_ ? _0521_ : _0536_);
	assign _0538_ = (_0305_ ? _0506_ : _0537_);
	assign _0539_ = (_0342_ ? _0475_ : _0538_);
	assign _0540_ = (_0412_ ? _0406_ : _0539_);
	assign \mchip.dut.demux.I [0] = ~_0540_;
	assign _0541_ = (_0254_ ? \mchip.dut.memory.M[127] [1] : \mchip.dut.memory.M[126] [1]);
	assign _0542_ = (_0254_ ? \mchip.dut.memory.M[125] [1] : \mchip.dut.memory.M[124] [1]);
	assign _0543_ = (_0259_ ? _0541_ : _0542_);
	assign _0544_ = (_0254_ ? \mchip.dut.memory.M[123] [1] : \mchip.dut.memory.M[122] [1]);
	assign _0545_ = (_0254_ ? \mchip.dut.memory.M[121] [1] : \mchip.dut.memory.M[120] [1]);
	assign _0546_ = (_0259_ ? _0544_ : _0545_);
	assign _0547_ = (_0268_ ? _0543_ : _0546_);
	assign _0548_ = (_0254_ ? \mchip.dut.memory.M[119] [1] : \mchip.dut.memory.M[118] [1]);
	assign _0549_ = (_0254_ ? \mchip.dut.memory.M[117] [1] : \mchip.dut.memory.M[116] [1]);
	assign _0550_ = (_0259_ ? _0548_ : _0549_);
	assign _0551_ = (_0254_ ? \mchip.dut.memory.M[115] [1] : \mchip.dut.memory.M[114] [1]);
	assign _0552_ = (_0254_ ? \mchip.dut.memory.M[113] [1] : \mchip.dut.memory.M[112] [1]);
	assign _0553_ = (_0259_ ? _0551_ : _0552_);
	assign _0554_ = (_0268_ ? _0550_ : _0553_);
	assign _0555_ = (_0282_ ? _0547_ : _0554_);
	assign _0556_ = (_0254_ ? \mchip.dut.memory.M[111] [1] : \mchip.dut.memory.M[110] [1]);
	assign _0557_ = (_0254_ ? \mchip.dut.memory.M[109] [1] : \mchip.dut.memory.M[108] [1]);
	assign _0558_ = (_0259_ ? _0556_ : _0557_);
	assign _0559_ = (_0254_ ? \mchip.dut.memory.M[107] [1] : \mchip.dut.memory.M[106] [1]);
	assign _0560_ = (_0254_ ? \mchip.dut.memory.M[105] [1] : \mchip.dut.memory.M[104] [1]);
	assign _0561_ = (_0259_ ? _0559_ : _0560_);
	assign _0562_ = (_0268_ ? _0558_ : _0561_);
	assign _0563_ = (_0254_ ? \mchip.dut.memory.M[103] [1] : \mchip.dut.memory.M[102] [1]);
	assign _0564_ = (_0254_ ? \mchip.dut.memory.M[101] [1] : \mchip.dut.memory.M[100] [1]);
	assign _0565_ = (_0259_ ? _0563_ : _0564_);
	assign _0566_ = (_0254_ ? \mchip.dut.memory.M[99] [1] : \mchip.dut.memory.M[98] [1]);
	assign _0567_ = (_0254_ ? \mchip.dut.memory.M[97] [1] : \mchip.dut.memory.M[96] [1]);
	assign _0568_ = (_0259_ ? _0566_ : _0567_);
	assign _0569_ = (_0268_ ? _0565_ : _0568_);
	assign _0570_ = (_0282_ ? _0562_ : _0569_);
	assign _0571_ = (_0305_ ? _0555_ : _0570_);
	assign _0572_ = (_0254_ ? \mchip.dut.memory.M[95] [1] : \mchip.dut.memory.M[94] [1]);
	assign _0573_ = (_0254_ ? \mchip.dut.memory.M[93] [1] : \mchip.dut.memory.M[92] [1]);
	assign _0574_ = (_0259_ ? _0572_ : _0573_);
	assign _0575_ = (_0254_ ? \mchip.dut.memory.M[91] [1] : \mchip.dut.memory.M[90] [1]);
	assign _0576_ = (_0254_ ? \mchip.dut.memory.M[89] [1] : \mchip.dut.memory.M[88] [1]);
	assign _0577_ = (_0259_ ? _0575_ : _0576_);
	assign _0578_ = (_0268_ ? _0574_ : _0577_);
	assign _0579_ = (_0254_ ? \mchip.dut.memory.M[87] [1] : \mchip.dut.memory.M[86] [1]);
	assign _0580_ = (_0254_ ? \mchip.dut.memory.M[85] [1] : \mchip.dut.memory.M[84] [1]);
	assign _0581_ = (_0259_ ? _0579_ : _0580_);
	assign _0582_ = (_0254_ ? \mchip.dut.memory.M[83] [1] : \mchip.dut.memory.M[82] [1]);
	assign _0583_ = (_0254_ ? \mchip.dut.memory.M[81] [1] : \mchip.dut.memory.M[80] [1]);
	assign _0584_ = (_0259_ ? _0582_ : _0583_);
	assign _0585_ = (_0268_ ? _0581_ : _0584_);
	assign _0586_ = (_0282_ ? _0578_ : _0585_);
	assign _0587_ = (_0254_ ? \mchip.dut.memory.M[79] [1] : \mchip.dut.memory.M[78] [1]);
	assign _0588_ = (_0254_ ? \mchip.dut.memory.M[77] [1] : \mchip.dut.memory.M[76] [1]);
	assign _0589_ = (_0259_ ? _0587_ : _0588_);
	assign _0590_ = (_0254_ ? \mchip.dut.memory.M[75] [1] : \mchip.dut.memory.M[74] [1]);
	assign _0591_ = (_0254_ ? \mchip.dut.memory.M[73] [1] : \mchip.dut.memory.M[72] [1]);
	assign _0592_ = (_0259_ ? _0590_ : _0591_);
	assign _0593_ = (_0268_ ? _0589_ : _0592_);
	assign _0594_ = (_0254_ ? \mchip.dut.memory.M[71] [1] : \mchip.dut.memory.M[70] [1]);
	assign _0595_ = (_0254_ ? \mchip.dut.memory.M[69] [1] : \mchip.dut.memory.M[68] [1]);
	assign _0596_ = (_0259_ ? _0594_ : _0595_);
	assign _0597_ = (_0254_ ? \mchip.dut.memory.M[67] [1] : \mchip.dut.memory.M[66] [1]);
	assign _0598_ = (_0254_ ? \mchip.dut.memory.M[65] [1] : \mchip.dut.memory.M[64] [1]);
	assign _0599_ = (_0259_ ? _0597_ : _0598_);
	assign _0600_ = (_0268_ ? _0596_ : _0599_);
	assign _0601_ = (_0282_ ? _0593_ : _0600_);
	assign _0602_ = (_0305_ ? _0586_ : _0601_);
	assign _0603_ = (_0342_ ? _0571_ : _0602_);
	assign _0604_ = (_0254_ ? \mchip.dut.memory.M[63] [1] : \mchip.dut.memory.M[62] [1]);
	assign _0605_ = (_0254_ ? \mchip.dut.memory.M[61] [1] : \mchip.dut.memory.M[60] [1]);
	assign _0606_ = (_0259_ ? _0604_ : _0605_);
	assign _0607_ = (_0254_ ? \mchip.dut.memory.M[59] [1] : \mchip.dut.memory.M[58] [1]);
	assign _0608_ = (_0254_ ? \mchip.dut.memory.M[57] [1] : \mchip.dut.memory.M[56] [1]);
	assign _0609_ = (_0259_ ? _0607_ : _0608_);
	assign _0610_ = (_0268_ ? _0606_ : _0609_);
	assign _0611_ = (_0254_ ? \mchip.dut.memory.M[55] [1] : \mchip.dut.memory.M[54] [1]);
	assign _0612_ = (_0254_ ? \mchip.dut.memory.M[53] [1] : \mchip.dut.memory.M[52] [1]);
	assign _0613_ = (_0259_ ? _0611_ : _0612_);
	assign _0614_ = (_0254_ ? \mchip.dut.memory.M[51] [1] : \mchip.dut.memory.M[50] [1]);
	assign _0615_ = (_0254_ ? \mchip.dut.memory.M[49] [1] : \mchip.dut.memory.M[48] [1]);
	assign _0616_ = (_0259_ ? _0614_ : _0615_);
	assign _0617_ = (_0268_ ? _0613_ : _0616_);
	assign _0618_ = (_0282_ ? _0610_ : _0617_);
	assign _0619_ = (_0254_ ? \mchip.dut.memory.M[47] [1] : \mchip.dut.memory.M[46] [1]);
	assign _0620_ = (_0254_ ? \mchip.dut.memory.M[45] [1] : \mchip.dut.memory.M[44] [1]);
	assign _0621_ = (_0259_ ? _0619_ : _0620_);
	assign _0622_ = (_0254_ ? \mchip.dut.memory.M[43] [1] : \mchip.dut.memory.M[42] [1]);
	assign _0623_ = (_0254_ ? \mchip.dut.memory.M[41] [1] : \mchip.dut.memory.M[40] [1]);
	assign _0624_ = (_0259_ ? _0622_ : _0623_);
	assign _0625_ = (_0268_ ? _0621_ : _0624_);
	assign _0626_ = (_0254_ ? \mchip.dut.memory.M[39] [1] : \mchip.dut.memory.M[38] [1]);
	assign _0627_ = (_0254_ ? \mchip.dut.memory.M[37] [1] : \mchip.dut.memory.M[36] [1]);
	assign _0628_ = (_0259_ ? _0626_ : _0627_);
	assign _0629_ = (_0254_ ? \mchip.dut.memory.M[35] [1] : \mchip.dut.memory.M[34] [1]);
	assign _0630_ = (_0254_ ? \mchip.dut.memory.M[33] [1] : \mchip.dut.memory.M[32] [1]);
	assign _0631_ = (_0259_ ? _0629_ : _0630_);
	assign _0632_ = (_0268_ ? _0628_ : _0631_);
	assign _0633_ = (_0282_ ? _0625_ : _0632_);
	assign _0634_ = (_0305_ ? _0618_ : _0633_);
	assign _0635_ = (_0254_ ? \mchip.dut.memory.M[31] [1] : \mchip.dut.memory.M[30] [1]);
	assign _0636_ = (_0254_ ? \mchip.dut.memory.M[29] [1] : \mchip.dut.memory.M[28] [1]);
	assign _0637_ = (_0259_ ? _0635_ : _0636_);
	assign _0638_ = (_0254_ ? \mchip.dut.memory.M[27] [1] : \mchip.dut.memory.M[26] [1]);
	assign _0639_ = (_0254_ ? \mchip.dut.memory.M[25] [1] : \mchip.dut.memory.M[24] [1]);
	assign _0640_ = (_0259_ ? _0638_ : _0639_);
	assign _0641_ = (_0268_ ? _0637_ : _0640_);
	assign _0642_ = (_0254_ ? \mchip.dut.memory.M[23] [1] : \mchip.dut.memory.M[22] [1]);
	assign _0643_ = (_0254_ ? \mchip.dut.memory.M[21] [1] : \mchip.dut.memory.M[20] [1]);
	assign _0644_ = (_0259_ ? _0642_ : _0643_);
	assign _0645_ = (_0254_ ? \mchip.dut.memory.M[19] [1] : \mchip.dut.memory.M[18] [1]);
	assign _0646_ = (_0254_ ? \mchip.dut.memory.M[17] [1] : \mchip.dut.memory.M[16] [1]);
	assign _0647_ = (_0259_ ? _0645_ : _0646_);
	assign _0648_ = (_0268_ ? _0644_ : _0647_);
	assign _0649_ = (_0282_ ? _0641_ : _0648_);
	assign _0650_ = (_0254_ ? \mchip.dut.memory.M[15] [1] : \mchip.dut.memory.M[14] [1]);
	assign _0651_ = (_0254_ ? \mchip.dut.memory.M[13] [1] : \mchip.dut.memory.M[12] [1]);
	assign _0652_ = (_0259_ ? _0650_ : _0651_);
	assign _0653_ = (_0254_ ? \mchip.dut.memory.M[11] [1] : \mchip.dut.memory.M[10] [1]);
	assign _0654_ = (_0254_ ? \mchip.dut.memory.M[9] [1] : \mchip.dut.memory.M[8] [1]);
	assign _0655_ = (_0259_ ? _0653_ : _0654_);
	assign _0656_ = (_0268_ ? _0652_ : _0655_);
	assign _0657_ = (_0254_ ? \mchip.dut.memory.M[7] [1] : \mchip.dut.memory.M[6] [1]);
	assign _0658_ = (_0254_ ? \mchip.dut.memory.M[5] [1] : \mchip.dut.memory.M[4] [1]);
	assign _0659_ = (_0259_ ? _0657_ : _0658_);
	assign _0660_ = (_0254_ ? \mchip.dut.memory.M[3] [1] : \mchip.dut.memory.M[2] [1]);
	assign _0661_ = (_0254_ ? \mchip.dut.memory.M[1] [1] : \mchip.dut.memory.M[0] [1]);
	assign _0662_ = (_0259_ ? _0660_ : _0661_);
	assign _0663_ = (_0268_ ? _0659_ : _0662_);
	assign _0664_ = (_0282_ ? _0656_ : _0663_);
	assign _0665_ = (_0305_ ? _0649_ : _0664_);
	assign _0666_ = (_0342_ ? _0634_ : _0665_);
	assign \mchip.dut.demux.I [1] = (_0412_ ? _0603_ : _0666_);
	assign _0667_ = (_0254_ ? \mchip.dut.memory.M[127] [2] : \mchip.dut.memory.M[126] [2]);
	assign _0668_ = (_0254_ ? \mchip.dut.memory.M[125] [2] : \mchip.dut.memory.M[124] [2]);
	assign _0669_ = (_0259_ ? _0667_ : _0668_);
	assign _0670_ = (_0254_ ? \mchip.dut.memory.M[123] [2] : \mchip.dut.memory.M[122] [2]);
	assign _0671_ = (_0254_ ? \mchip.dut.memory.M[121] [2] : \mchip.dut.memory.M[120] [2]);
	assign _0672_ = (_0259_ ? _0670_ : _0671_);
	assign _0673_ = (_0268_ ? _0669_ : _0672_);
	assign _0674_ = (_0254_ ? \mchip.dut.memory.M[119] [2] : \mchip.dut.memory.M[118] [2]);
	assign _0675_ = (_0254_ ? \mchip.dut.memory.M[117] [2] : \mchip.dut.memory.M[116] [2]);
	assign _0676_ = (_0259_ ? _0674_ : _0675_);
	assign _0677_ = (_0254_ ? \mchip.dut.memory.M[115] [2] : \mchip.dut.memory.M[114] [2]);
	assign _0678_ = (_0254_ ? \mchip.dut.memory.M[113] [2] : \mchip.dut.memory.M[112] [2]);
	assign _0679_ = (_0259_ ? _0677_ : _0678_);
	assign _0680_ = (_0268_ ? _0676_ : _0679_);
	assign _0681_ = (_0282_ ? _0673_ : _0680_);
	assign _0682_ = (_0254_ ? \mchip.dut.memory.M[111] [2] : \mchip.dut.memory.M[110] [2]);
	assign _0683_ = (_0254_ ? \mchip.dut.memory.M[109] [2] : \mchip.dut.memory.M[108] [2]);
	assign _0684_ = (_0259_ ? _0682_ : _0683_);
	assign _0685_ = (_0254_ ? \mchip.dut.memory.M[107] [2] : \mchip.dut.memory.M[106] [2]);
	assign _0686_ = (_0254_ ? \mchip.dut.memory.M[105] [2] : \mchip.dut.memory.M[104] [2]);
	assign _0687_ = (_0259_ ? _0685_ : _0686_);
	assign _0688_ = (_0268_ ? _0684_ : _0687_);
	assign _0689_ = (_0254_ ? \mchip.dut.memory.M[103] [2] : \mchip.dut.memory.M[102] [2]);
	assign _0690_ = (_0254_ ? \mchip.dut.memory.M[101] [2] : \mchip.dut.memory.M[100] [2]);
	assign _0691_ = (_0259_ ? _0689_ : _0690_);
	assign _0692_ = (_0254_ ? \mchip.dut.memory.M[99] [2] : \mchip.dut.memory.M[98] [2]);
	assign _0693_ = (_0254_ ? \mchip.dut.memory.M[97] [2] : \mchip.dut.memory.M[96] [2]);
	assign _0694_ = (_0259_ ? _0692_ : _0693_);
	assign _0695_ = (_0268_ ? _0691_ : _0694_);
	assign _0696_ = (_0282_ ? _0688_ : _0695_);
	assign _0697_ = (_0305_ ? _0681_ : _0696_);
	assign _0698_ = (_0254_ ? \mchip.dut.memory.M[95] [2] : \mchip.dut.memory.M[94] [2]);
	assign _0699_ = (_0254_ ? \mchip.dut.memory.M[93] [2] : \mchip.dut.memory.M[92] [2]);
	assign _0700_ = (_0259_ ? _0698_ : _0699_);
	assign _0701_ = (_0254_ ? \mchip.dut.memory.M[91] [2] : \mchip.dut.memory.M[90] [2]);
	assign _0702_ = (_0254_ ? \mchip.dut.memory.M[89] [2] : \mchip.dut.memory.M[88] [2]);
	assign _0703_ = (_0259_ ? _0701_ : _0702_);
	assign _0704_ = (_0268_ ? _0700_ : _0703_);
	assign _0705_ = (_0254_ ? \mchip.dut.memory.M[87] [2] : \mchip.dut.memory.M[86] [2]);
	assign _0706_ = (_0254_ ? \mchip.dut.memory.M[85] [2] : \mchip.dut.memory.M[84] [2]);
	assign _0707_ = (_0259_ ? _0705_ : _0706_);
	assign _0708_ = (_0254_ ? \mchip.dut.memory.M[83] [2] : \mchip.dut.memory.M[82] [2]);
	assign _0709_ = (_0254_ ? \mchip.dut.memory.M[81] [2] : \mchip.dut.memory.M[80] [2]);
	assign _0710_ = (_0259_ ? _0708_ : _0709_);
	assign _0711_ = (_0268_ ? _0707_ : _0710_);
	assign _0712_ = (_0282_ ? _0704_ : _0711_);
	assign _0713_ = (_0254_ ? \mchip.dut.memory.M[79] [2] : \mchip.dut.memory.M[78] [2]);
	assign _0714_ = (_0254_ ? \mchip.dut.memory.M[77] [2] : \mchip.dut.memory.M[76] [2]);
	assign _0715_ = (_0259_ ? _0713_ : _0714_);
	assign _0716_ = (_0254_ ? \mchip.dut.memory.M[75] [2] : \mchip.dut.memory.M[74] [2]);
	assign _0717_ = (_0254_ ? \mchip.dut.memory.M[73] [2] : \mchip.dut.memory.M[72] [2]);
	assign _0718_ = (_0259_ ? _0716_ : _0717_);
	assign _0719_ = (_0268_ ? _0715_ : _0718_);
	assign _0720_ = (_0254_ ? \mchip.dut.memory.M[71] [2] : \mchip.dut.memory.M[70] [2]);
	assign _0721_ = (_0254_ ? \mchip.dut.memory.M[69] [2] : \mchip.dut.memory.M[68] [2]);
	assign _0722_ = (_0259_ ? _0720_ : _0721_);
	assign _0723_ = (_0254_ ? \mchip.dut.memory.M[67] [2] : \mchip.dut.memory.M[66] [2]);
	assign _0724_ = (_0254_ ? \mchip.dut.memory.M[65] [2] : \mchip.dut.memory.M[64] [2]);
	assign _0725_ = (_0259_ ? _0723_ : _0724_);
	assign _0726_ = (_0268_ ? _0722_ : _0725_);
	assign _0727_ = (_0282_ ? _0719_ : _0726_);
	assign _0728_ = (_0305_ ? _0712_ : _0727_);
	assign _0729_ = (_0342_ ? _0697_ : _0728_);
	assign _0730_ = (_0254_ ? \mchip.dut.memory.M[63] [2] : \mchip.dut.memory.M[62] [2]);
	assign _0731_ = (_0254_ ? \mchip.dut.memory.M[61] [2] : \mchip.dut.memory.M[60] [2]);
	assign _0732_ = (_0259_ ? _0730_ : _0731_);
	assign _0733_ = (_0254_ ? \mchip.dut.memory.M[59] [2] : \mchip.dut.memory.M[58] [2]);
	assign _0734_ = (_0254_ ? \mchip.dut.memory.M[57] [2] : \mchip.dut.memory.M[56] [2]);
	assign _0735_ = (_0259_ ? _0733_ : _0734_);
	assign _0736_ = (_0268_ ? _0732_ : _0735_);
	assign _0737_ = (_0254_ ? \mchip.dut.memory.M[55] [2] : \mchip.dut.memory.M[54] [2]);
	assign _0738_ = (_0254_ ? \mchip.dut.memory.M[53] [2] : \mchip.dut.memory.M[52] [2]);
	assign _0739_ = (_0259_ ? _0737_ : _0738_);
	assign _0740_ = (_0254_ ? \mchip.dut.memory.M[51] [2] : \mchip.dut.memory.M[50] [2]);
	assign _0741_ = (_0254_ ? \mchip.dut.memory.M[49] [2] : \mchip.dut.memory.M[48] [2]);
	assign _0742_ = (_0259_ ? _0740_ : _0741_);
	assign _0743_ = (_0268_ ? _0739_ : _0742_);
	assign _0744_ = (_0282_ ? _0736_ : _0743_);
	assign _0745_ = (_0254_ ? \mchip.dut.memory.M[47] [2] : \mchip.dut.memory.M[46] [2]);
	assign _0746_ = (_0254_ ? \mchip.dut.memory.M[45] [2] : \mchip.dut.memory.M[44] [2]);
	assign _0747_ = (_0259_ ? _0745_ : _0746_);
	assign _0748_ = (_0254_ ? \mchip.dut.memory.M[43] [2] : \mchip.dut.memory.M[42] [2]);
	assign _0749_ = (_0254_ ? \mchip.dut.memory.M[41] [2] : \mchip.dut.memory.M[40] [2]);
	assign _0750_ = (_0259_ ? _0748_ : _0749_);
	assign _0751_ = (_0268_ ? _0747_ : _0750_);
	assign _0752_ = (_0254_ ? \mchip.dut.memory.M[39] [2] : \mchip.dut.memory.M[38] [2]);
	assign _0753_ = (_0254_ ? \mchip.dut.memory.M[37] [2] : \mchip.dut.memory.M[36] [2]);
	assign _0754_ = (_0259_ ? _0752_ : _0753_);
	assign _0755_ = (_0254_ ? \mchip.dut.memory.M[35] [2] : \mchip.dut.memory.M[34] [2]);
	assign _0756_ = (_0254_ ? \mchip.dut.memory.M[33] [2] : \mchip.dut.memory.M[32] [2]);
	assign _0757_ = (_0259_ ? _0755_ : _0756_);
	assign _0758_ = (_0268_ ? _0754_ : _0757_);
	assign _0759_ = (_0282_ ? _0751_ : _0758_);
	assign _0760_ = (_0305_ ? _0744_ : _0759_);
	assign _0761_ = (_0254_ ? \mchip.dut.memory.M[31] [2] : \mchip.dut.memory.M[30] [2]);
	assign _0762_ = (_0254_ ? \mchip.dut.memory.M[29] [2] : \mchip.dut.memory.M[28] [2]);
	assign _0763_ = (_0259_ ? _0761_ : _0762_);
	assign _0764_ = (_0254_ ? \mchip.dut.memory.M[27] [2] : \mchip.dut.memory.M[26] [2]);
	assign _0765_ = (_0254_ ? \mchip.dut.memory.M[25] [2] : \mchip.dut.memory.M[24] [2]);
	assign _0766_ = (_0259_ ? _0764_ : _0765_);
	assign _0767_ = (_0268_ ? _0763_ : _0766_);
	assign _0768_ = (_0254_ ? \mchip.dut.memory.M[23] [2] : \mchip.dut.memory.M[22] [2]);
	assign _0769_ = (_0254_ ? \mchip.dut.memory.M[21] [2] : \mchip.dut.memory.M[20] [2]);
	assign _0770_ = (_0259_ ? _0768_ : _0769_);
	assign _0771_ = (_0254_ ? \mchip.dut.memory.M[19] [2] : \mchip.dut.memory.M[18] [2]);
	assign _0772_ = (_0254_ ? \mchip.dut.memory.M[17] [2] : \mchip.dut.memory.M[16] [2]);
	assign _0773_ = (_0259_ ? _0771_ : _0772_);
	assign _0774_ = (_0268_ ? _0770_ : _0773_);
	assign _0775_ = (_0282_ ? _0767_ : _0774_);
	assign _0776_ = (_0254_ ? \mchip.dut.memory.M[15] [2] : \mchip.dut.memory.M[14] [2]);
	assign _0777_ = (_0254_ ? \mchip.dut.memory.M[13] [2] : \mchip.dut.memory.M[12] [2]);
	assign _0778_ = (_0259_ ? _0776_ : _0777_);
	assign _0779_ = (_0254_ ? \mchip.dut.memory.M[11] [2] : \mchip.dut.memory.M[10] [2]);
	assign _0780_ = (_0254_ ? \mchip.dut.memory.M[9] [2] : \mchip.dut.memory.M[8] [2]);
	assign _0781_ = (_0259_ ? _0779_ : _0780_);
	assign _0782_ = (_0268_ ? _0778_ : _0781_);
	assign _0783_ = (_0254_ ? \mchip.dut.memory.M[7] [2] : \mchip.dut.memory.M[6] [2]);
	assign _0784_ = (_0254_ ? \mchip.dut.memory.M[5] [2] : \mchip.dut.memory.M[4] [2]);
	assign _0785_ = (_0259_ ? _0783_ : _0784_);
	assign _0786_ = (_0254_ ? \mchip.dut.memory.M[3] [2] : \mchip.dut.memory.M[2] [2]);
	assign _0787_ = (_0254_ ? \mchip.dut.memory.M[1] [2] : \mchip.dut.memory.M[0] [2]);
	assign _0788_ = (_0259_ ? _0786_ : _0787_);
	assign _0789_ = (_0268_ ? _0785_ : _0788_);
	assign _0790_ = (_0282_ ? _0782_ : _0789_);
	assign _0791_ = (_0305_ ? _0775_ : _0790_);
	assign _0792_ = (_0342_ ? _0760_ : _0791_);
	assign \mchip.dut.demux.I [2] = (_0412_ ? _0729_ : _0792_);
	assign _0793_ = (_0254_ ? \mchip.dut.memory.M[127] [3] : \mchip.dut.memory.M[126] [3]);
	assign _0794_ = (_0254_ ? \mchip.dut.memory.M[125] [3] : \mchip.dut.memory.M[124] [3]);
	assign _0795_ = (_0259_ ? _0793_ : _0794_);
	assign _0796_ = (_0254_ ? \mchip.dut.memory.M[123] [3] : \mchip.dut.memory.M[122] [3]);
	assign _0797_ = (_0254_ ? \mchip.dut.memory.M[121] [3] : \mchip.dut.memory.M[120] [3]);
	assign _0798_ = (_0259_ ? _0796_ : _0797_);
	assign _0799_ = (_0268_ ? _0795_ : _0798_);
	assign _0800_ = (_0254_ ? \mchip.dut.memory.M[119] [3] : \mchip.dut.memory.M[118] [3]);
	assign _0801_ = (_0254_ ? \mchip.dut.memory.M[117] [3] : \mchip.dut.memory.M[116] [3]);
	assign _0802_ = (_0259_ ? _0800_ : _0801_);
	assign _0803_ = (_0254_ ? \mchip.dut.memory.M[115] [3] : \mchip.dut.memory.M[114] [3]);
	assign _0804_ = (_0254_ ? \mchip.dut.memory.M[113] [3] : \mchip.dut.memory.M[112] [3]);
	assign _0805_ = (_0259_ ? _0803_ : _0804_);
	assign _0806_ = (_0268_ ? _0802_ : _0805_);
	assign _0807_ = (_0282_ ? _0799_ : _0806_);
	assign _0808_ = (_0254_ ? \mchip.dut.memory.M[111] [3] : \mchip.dut.memory.M[110] [3]);
	assign _0809_ = (_0254_ ? \mchip.dut.memory.M[109] [3] : \mchip.dut.memory.M[108] [3]);
	assign _0810_ = (_0259_ ? _0808_ : _0809_);
	assign _0811_ = (_0254_ ? \mchip.dut.memory.M[107] [3] : \mchip.dut.memory.M[106] [3]);
	assign _0812_ = (_0254_ ? \mchip.dut.memory.M[105] [3] : \mchip.dut.memory.M[104] [3]);
	assign _0813_ = (_0259_ ? _0811_ : _0812_);
	assign _0814_ = (_0268_ ? _0810_ : _0813_);
	assign _0815_ = (_0254_ ? \mchip.dut.memory.M[103] [3] : \mchip.dut.memory.M[102] [3]);
	assign _0816_ = (_0254_ ? \mchip.dut.memory.M[101] [3] : \mchip.dut.memory.M[100] [3]);
	assign _0817_ = (_0259_ ? _0815_ : _0816_);
	assign _0818_ = (_0254_ ? \mchip.dut.memory.M[99] [3] : \mchip.dut.memory.M[98] [3]);
	assign _0819_ = (_0254_ ? \mchip.dut.memory.M[97] [3] : \mchip.dut.memory.M[96] [3]);
	assign _0820_ = (_0259_ ? _0818_ : _0819_);
	assign _0821_ = (_0268_ ? _0817_ : _0820_);
	assign _0822_ = (_0282_ ? _0814_ : _0821_);
	assign _0823_ = (_0305_ ? _0807_ : _0822_);
	assign _0824_ = (_0254_ ? \mchip.dut.memory.M[95] [3] : \mchip.dut.memory.M[94] [3]);
	assign _0825_ = (_0254_ ? \mchip.dut.memory.M[93] [3] : \mchip.dut.memory.M[92] [3]);
	assign _0826_ = (_0259_ ? _0824_ : _0825_);
	assign _0827_ = (_0254_ ? \mchip.dut.memory.M[91] [3] : \mchip.dut.memory.M[90] [3]);
	assign _0828_ = (_0254_ ? \mchip.dut.memory.M[89] [3] : \mchip.dut.memory.M[88] [3]);
	assign _0829_ = (_0259_ ? _0827_ : _0828_);
	assign _0830_ = (_0268_ ? _0826_ : _0829_);
	assign _0831_ = (_0254_ ? \mchip.dut.memory.M[87] [3] : \mchip.dut.memory.M[86] [3]);
	assign _0832_ = (_0254_ ? \mchip.dut.memory.M[85] [3] : \mchip.dut.memory.M[84] [3]);
	assign _0833_ = (_0259_ ? _0831_ : _0832_);
	assign _0834_ = (_0254_ ? \mchip.dut.memory.M[83] [3] : \mchip.dut.memory.M[82] [3]);
	assign _0835_ = (_0254_ ? \mchip.dut.memory.M[81] [3] : \mchip.dut.memory.M[80] [3]);
	assign _0836_ = (_0259_ ? _0834_ : _0835_);
	assign _0837_ = (_0268_ ? _0833_ : _0836_);
	assign _0838_ = (_0282_ ? _0830_ : _0837_);
	assign _0839_ = (_0254_ ? \mchip.dut.memory.M[79] [3] : \mchip.dut.memory.M[78] [3]);
	assign _0840_ = (_0254_ ? \mchip.dut.memory.M[77] [3] : \mchip.dut.memory.M[76] [3]);
	assign _0841_ = (_0259_ ? _0839_ : _0840_);
	assign _0842_ = (_0254_ ? \mchip.dut.memory.M[75] [3] : \mchip.dut.memory.M[74] [3]);
	assign _0843_ = (_0254_ ? \mchip.dut.memory.M[73] [3] : \mchip.dut.memory.M[72] [3]);
	assign _0844_ = (_0259_ ? _0842_ : _0843_);
	assign _0845_ = (_0268_ ? _0841_ : _0844_);
	assign _0846_ = (_0254_ ? \mchip.dut.memory.M[71] [3] : \mchip.dut.memory.M[70] [3]);
	assign _0847_ = (_0254_ ? \mchip.dut.memory.M[69] [3] : \mchip.dut.memory.M[68] [3]);
	assign _0848_ = (_0259_ ? _0846_ : _0847_);
	assign _0849_ = (_0254_ ? \mchip.dut.memory.M[67] [3] : \mchip.dut.memory.M[66] [3]);
	assign _0850_ = (_0254_ ? \mchip.dut.memory.M[65] [3] : \mchip.dut.memory.M[64] [3]);
	assign _0851_ = (_0259_ ? _0849_ : _0850_);
	assign _0852_ = (_0268_ ? _0848_ : _0851_);
	assign _0853_ = (_0282_ ? _0845_ : _0852_);
	assign _0854_ = (_0305_ ? _0838_ : _0853_);
	assign _0855_ = (_0342_ ? _0823_ : _0854_);
	assign _0856_ = (_0254_ ? \mchip.dut.memory.M[63] [3] : \mchip.dut.memory.M[62] [3]);
	assign _0857_ = (_0254_ ? \mchip.dut.memory.M[61] [3] : \mchip.dut.memory.M[60] [3]);
	assign _0858_ = (_0259_ ? _0856_ : _0857_);
	assign _0859_ = (_0254_ ? \mchip.dut.memory.M[59] [3] : \mchip.dut.memory.M[58] [3]);
	assign _0860_ = (_0254_ ? \mchip.dut.memory.M[57] [3] : \mchip.dut.memory.M[56] [3]);
	assign _0861_ = (_0259_ ? _0859_ : _0860_);
	assign _0862_ = (_0268_ ? _0858_ : _0861_);
	assign _0863_ = (_0254_ ? \mchip.dut.memory.M[55] [3] : \mchip.dut.memory.M[54] [3]);
	assign _0864_ = (_0254_ ? \mchip.dut.memory.M[53] [3] : \mchip.dut.memory.M[52] [3]);
	assign _0865_ = (_0259_ ? _0863_ : _0864_);
	assign _0866_ = (_0254_ ? \mchip.dut.memory.M[51] [3] : \mchip.dut.memory.M[50] [3]);
	assign _0867_ = (_0254_ ? \mchip.dut.memory.M[49] [3] : \mchip.dut.memory.M[48] [3]);
	assign _0868_ = (_0259_ ? _0866_ : _0867_);
	assign _0869_ = (_0268_ ? _0865_ : _0868_);
	assign _0870_ = (_0282_ ? _0862_ : _0869_);
	assign _0871_ = (_0254_ ? \mchip.dut.memory.M[47] [3] : \mchip.dut.memory.M[46] [3]);
	assign _0872_ = (_0254_ ? \mchip.dut.memory.M[45] [3] : \mchip.dut.memory.M[44] [3]);
	assign _0873_ = (_0259_ ? _0871_ : _0872_);
	assign _0874_ = (_0254_ ? \mchip.dut.memory.M[43] [3] : \mchip.dut.memory.M[42] [3]);
	assign _0875_ = (_0254_ ? \mchip.dut.memory.M[41] [3] : \mchip.dut.memory.M[40] [3]);
	assign _0876_ = (_0259_ ? _0874_ : _0875_);
	assign _0877_ = (_0268_ ? _0873_ : _0876_);
	assign _0878_ = (_0254_ ? \mchip.dut.memory.M[39] [3] : \mchip.dut.memory.M[38] [3]);
	assign _0879_ = (_0254_ ? \mchip.dut.memory.M[37] [3] : \mchip.dut.memory.M[36] [3]);
	assign _0880_ = (_0259_ ? _0878_ : _0879_);
	assign _0881_ = (_0254_ ? \mchip.dut.memory.M[35] [3] : \mchip.dut.memory.M[34] [3]);
	assign _0882_ = (_0254_ ? \mchip.dut.memory.M[33] [3] : \mchip.dut.memory.M[32] [3]);
	assign _0883_ = (_0259_ ? _0881_ : _0882_);
	assign _0884_ = (_0268_ ? _0880_ : _0883_);
	assign _0885_ = (_0282_ ? _0877_ : _0884_);
	assign _0886_ = (_0305_ ? _0870_ : _0885_);
	assign _0887_ = (_0254_ ? \mchip.dut.memory.M[31] [3] : \mchip.dut.memory.M[30] [3]);
	assign _0888_ = (_0254_ ? \mchip.dut.memory.M[29] [3] : \mchip.dut.memory.M[28] [3]);
	assign _0889_ = (_0259_ ? _0887_ : _0888_);
	assign _0890_ = (_0254_ ? \mchip.dut.memory.M[27] [3] : \mchip.dut.memory.M[26] [3]);
	assign _0891_ = (_0254_ ? \mchip.dut.memory.M[25] [3] : \mchip.dut.memory.M[24] [3]);
	assign _0892_ = (_0259_ ? _0890_ : _0891_);
	assign _0893_ = (_0268_ ? _0889_ : _0892_);
	assign _0894_ = (_0254_ ? \mchip.dut.memory.M[23] [3] : \mchip.dut.memory.M[22] [3]);
	assign _0895_ = (_0254_ ? \mchip.dut.memory.M[21] [3] : \mchip.dut.memory.M[20] [3]);
	assign _0896_ = (_0259_ ? _0894_ : _0895_);
	assign _0897_ = (_0254_ ? \mchip.dut.memory.M[19] [3] : \mchip.dut.memory.M[18] [3]);
	assign _0898_ = (_0254_ ? \mchip.dut.memory.M[17] [3] : \mchip.dut.memory.M[16] [3]);
	assign _0899_ = (_0259_ ? _0897_ : _0898_);
	assign _0900_ = (_0268_ ? _0896_ : _0899_);
	assign _0901_ = (_0282_ ? _0893_ : _0900_);
	assign _0902_ = (_0254_ ? \mchip.dut.memory.M[15] [3] : \mchip.dut.memory.M[14] [3]);
	assign _0903_ = (_0254_ ? \mchip.dut.memory.M[13] [3] : \mchip.dut.memory.M[12] [3]);
	assign _0904_ = (_0259_ ? _0902_ : _0903_);
	assign _0905_ = (_0254_ ? \mchip.dut.memory.M[11] [3] : \mchip.dut.memory.M[10] [3]);
	assign _0906_ = (_0254_ ? \mchip.dut.memory.M[9] [3] : \mchip.dut.memory.M[8] [3]);
	assign _0907_ = (_0259_ ? _0905_ : _0906_);
	assign _0908_ = (_0268_ ? _0904_ : _0907_);
	assign _0909_ = (_0254_ ? \mchip.dut.memory.M[7] [3] : \mchip.dut.memory.M[6] [3]);
	assign _0910_ = (_0254_ ? \mchip.dut.memory.M[5] [3] : \mchip.dut.memory.M[4] [3]);
	assign _0911_ = (_0259_ ? _0909_ : _0910_);
	assign _0912_ = (_0254_ ? \mchip.dut.memory.M[3] [3] : \mchip.dut.memory.M[2] [3]);
	assign _0913_ = (_0254_ ? \mchip.dut.memory.M[1] [3] : \mchip.dut.memory.M[0] [3]);
	assign _0914_ = (_0259_ ? _0912_ : _0913_);
	assign _0915_ = (_0268_ ? _0911_ : _0914_);
	assign _0916_ = (_0282_ ? _0908_ : _0915_);
	assign _0917_ = (_0305_ ? _0901_ : _0916_);
	assign _0918_ = (_0342_ ? _0886_ : _0917_);
	assign \mchip.dut.demux.I [3] = (_0412_ ? _0855_ : _0918_);
	assign _0919_ = (_0254_ ? \mchip.dut.memory.M[127] [4] : \mchip.dut.memory.M[126] [4]);
	assign _0920_ = (_0254_ ? \mchip.dut.memory.M[125] [4] : \mchip.dut.memory.M[124] [4]);
	assign _0921_ = (_0259_ ? _0919_ : _0920_);
	assign _0922_ = (_0254_ ? \mchip.dut.memory.M[123] [4] : \mchip.dut.memory.M[122] [4]);
	assign _0923_ = (_0254_ ? \mchip.dut.memory.M[121] [4] : \mchip.dut.memory.M[120] [4]);
	assign _0924_ = (_0259_ ? _0922_ : _0923_);
	assign _0925_ = (_0268_ ? _0921_ : _0924_);
	assign _0926_ = (_0254_ ? \mchip.dut.memory.M[119] [4] : \mchip.dut.memory.M[118] [4]);
	assign _0927_ = (_0254_ ? \mchip.dut.memory.M[117] [4] : \mchip.dut.memory.M[116] [4]);
	assign _0928_ = (_0259_ ? _0926_ : _0927_);
	assign _0929_ = (_0254_ ? \mchip.dut.memory.M[115] [4] : \mchip.dut.memory.M[114] [4]);
	assign _0930_ = (_0254_ ? \mchip.dut.memory.M[113] [4] : \mchip.dut.memory.M[112] [4]);
	assign _0931_ = (_0259_ ? _0929_ : _0930_);
	assign _0932_ = (_0268_ ? _0928_ : _0931_);
	assign _0933_ = (_0282_ ? _0925_ : _0932_);
	assign _0934_ = (_0254_ ? \mchip.dut.memory.M[111] [4] : \mchip.dut.memory.M[110] [4]);
	assign _0935_ = (_0254_ ? \mchip.dut.memory.M[109] [4] : \mchip.dut.memory.M[108] [4]);
	assign _0936_ = (_0259_ ? _0934_ : _0935_);
	assign _0937_ = (_0254_ ? \mchip.dut.memory.M[107] [4] : \mchip.dut.memory.M[106] [4]);
	assign _0938_ = (_0254_ ? \mchip.dut.memory.M[105] [4] : \mchip.dut.memory.M[104] [4]);
	assign _0939_ = (_0259_ ? _0937_ : _0938_);
	assign _0940_ = (_0268_ ? _0936_ : _0939_);
	assign _0941_ = (_0254_ ? \mchip.dut.memory.M[103] [4] : \mchip.dut.memory.M[102] [4]);
	assign _0942_ = (_0254_ ? \mchip.dut.memory.M[101] [4] : \mchip.dut.memory.M[100] [4]);
	assign _0943_ = (_0259_ ? _0941_ : _0942_);
	assign _0944_ = (_0254_ ? \mchip.dut.memory.M[99] [4] : \mchip.dut.memory.M[98] [4]);
	assign _0945_ = (_0254_ ? \mchip.dut.memory.M[97] [4] : \mchip.dut.memory.M[96] [4]);
	assign _0946_ = (_0259_ ? _0944_ : _0945_);
	assign _0947_ = (_0268_ ? _0943_ : _0946_);
	assign _0948_ = (_0282_ ? _0940_ : _0947_);
	assign _0949_ = (_0305_ ? _0933_ : _0948_);
	assign _0950_ = (_0254_ ? \mchip.dut.memory.M[95] [4] : \mchip.dut.memory.M[94] [4]);
	assign _0951_ = (_0254_ ? \mchip.dut.memory.M[93] [4] : \mchip.dut.memory.M[92] [4]);
	assign _0952_ = (_0259_ ? _0950_ : _0951_);
	assign _0953_ = (_0254_ ? \mchip.dut.memory.M[91] [4] : \mchip.dut.memory.M[90] [4]);
	assign _0954_ = (_0254_ ? \mchip.dut.memory.M[89] [4] : \mchip.dut.memory.M[88] [4]);
	assign _0955_ = (_0259_ ? _0953_ : _0954_);
	assign _0956_ = (_0268_ ? _0952_ : _0955_);
	assign _0957_ = (_0254_ ? \mchip.dut.memory.M[87] [4] : \mchip.dut.memory.M[86] [4]);
	assign _0958_ = (_0254_ ? \mchip.dut.memory.M[85] [4] : \mchip.dut.memory.M[84] [4]);
	assign _0959_ = (_0259_ ? _0957_ : _0958_);
	assign _0960_ = (_0254_ ? \mchip.dut.memory.M[83] [4] : \mchip.dut.memory.M[82] [4]);
	assign _0961_ = (_0254_ ? \mchip.dut.memory.M[81] [4] : \mchip.dut.memory.M[80] [4]);
	assign _0962_ = (_0259_ ? _0960_ : _0961_);
	assign _0963_ = (_0268_ ? _0959_ : _0962_);
	assign _0964_ = (_0282_ ? _0956_ : _0963_);
	assign _0965_ = (_0254_ ? \mchip.dut.memory.M[79] [4] : \mchip.dut.memory.M[78] [4]);
	assign _0966_ = (_0254_ ? \mchip.dut.memory.M[77] [4] : \mchip.dut.memory.M[76] [4]);
	assign _0967_ = (_0259_ ? _0965_ : _0966_);
	assign _0968_ = (_0254_ ? \mchip.dut.memory.M[75] [4] : \mchip.dut.memory.M[74] [4]);
	assign _0969_ = (_0254_ ? \mchip.dut.memory.M[73] [4] : \mchip.dut.memory.M[72] [4]);
	assign _0970_ = (_0259_ ? _0968_ : _0969_);
	assign _0971_ = (_0268_ ? _0967_ : _0970_);
	assign _0972_ = (_0254_ ? \mchip.dut.memory.M[71] [4] : \mchip.dut.memory.M[70] [4]);
	assign _0973_ = (_0254_ ? \mchip.dut.memory.M[69] [4] : \mchip.dut.memory.M[68] [4]);
	assign _0974_ = (_0259_ ? _0972_ : _0973_);
	assign _0975_ = (_0254_ ? \mchip.dut.memory.M[67] [4] : \mchip.dut.memory.M[66] [4]);
	assign _0976_ = (_0254_ ? \mchip.dut.memory.M[65] [4] : \mchip.dut.memory.M[64] [4]);
	assign _0977_ = (_0259_ ? _0975_ : _0976_);
	assign _0978_ = (_0268_ ? _0974_ : _0977_);
	assign _0979_ = (_0282_ ? _0971_ : _0978_);
	assign _0980_ = (_0305_ ? _0964_ : _0979_);
	assign _0981_ = (_0342_ ? _0949_ : _0980_);
	assign _0982_ = (_0254_ ? \mchip.dut.memory.M[63] [4] : \mchip.dut.memory.M[62] [4]);
	assign _0983_ = (_0254_ ? \mchip.dut.memory.M[61] [4] : \mchip.dut.memory.M[60] [4]);
	assign _0984_ = (_0259_ ? _0982_ : _0983_);
	assign _0985_ = (_0254_ ? \mchip.dut.memory.M[59] [4] : \mchip.dut.memory.M[58] [4]);
	assign _0986_ = (_0254_ ? \mchip.dut.memory.M[57] [4] : \mchip.dut.memory.M[56] [4]);
	assign _0987_ = (_0259_ ? _0985_ : _0986_);
	assign _0988_ = (_0268_ ? _0984_ : _0987_);
	assign _0989_ = (_0254_ ? \mchip.dut.memory.M[55] [4] : \mchip.dut.memory.M[54] [4]);
	assign _0990_ = (_0254_ ? \mchip.dut.memory.M[53] [4] : \mchip.dut.memory.M[52] [4]);
	assign _0991_ = (_0259_ ? _0989_ : _0990_);
	assign _0992_ = (_0254_ ? \mchip.dut.memory.M[51] [4] : \mchip.dut.memory.M[50] [4]);
	assign _0993_ = (_0254_ ? \mchip.dut.memory.M[49] [4] : \mchip.dut.memory.M[48] [4]);
	assign _0994_ = (_0259_ ? _0992_ : _0993_);
	assign _0995_ = (_0268_ ? _0991_ : _0994_);
	assign _0996_ = (_0282_ ? _0988_ : _0995_);
	assign _0997_ = (_0254_ ? \mchip.dut.memory.M[47] [4] : \mchip.dut.memory.M[46] [4]);
	assign _0998_ = (_0254_ ? \mchip.dut.memory.M[45] [4] : \mchip.dut.memory.M[44] [4]);
	assign _0999_ = (_0259_ ? _0997_ : _0998_);
	assign _1000_ = (_0254_ ? \mchip.dut.memory.M[43] [4] : \mchip.dut.memory.M[42] [4]);
	assign _1001_ = (_0254_ ? \mchip.dut.memory.M[41] [4] : \mchip.dut.memory.M[40] [4]);
	assign _1002_ = (_0259_ ? _1000_ : _1001_);
	assign _1003_ = (_0268_ ? _0999_ : _1002_);
	assign _1004_ = (_0254_ ? \mchip.dut.memory.M[39] [4] : \mchip.dut.memory.M[38] [4]);
	assign _1005_ = (_0254_ ? \mchip.dut.memory.M[37] [4] : \mchip.dut.memory.M[36] [4]);
	assign _1006_ = (_0259_ ? _1004_ : _1005_);
	assign _1007_ = (_0254_ ? \mchip.dut.memory.M[35] [4] : \mchip.dut.memory.M[34] [4]);
	assign _1008_ = (_0254_ ? \mchip.dut.memory.M[33] [4] : \mchip.dut.memory.M[32] [4]);
	assign _1009_ = (_0259_ ? _1007_ : _1008_);
	assign _1010_ = (_0268_ ? _1006_ : _1009_);
	assign _1011_ = (_0282_ ? _1003_ : _1010_);
	assign _1012_ = (_0305_ ? _0996_ : _1011_);
	assign _1013_ = (_0254_ ? \mchip.dut.memory.M[31] [4] : \mchip.dut.memory.M[30] [4]);
	assign _1014_ = (_0254_ ? \mchip.dut.memory.M[29] [4] : \mchip.dut.memory.M[28] [4]);
	assign _1015_ = (_0259_ ? _1013_ : _1014_);
	assign _1016_ = (_0254_ ? \mchip.dut.memory.M[27] [4] : \mchip.dut.memory.M[26] [4]);
	assign _1017_ = (_0254_ ? \mchip.dut.memory.M[25] [4] : \mchip.dut.memory.M[24] [4]);
	assign _1018_ = (_0259_ ? _1016_ : _1017_);
	assign _1019_ = (_0268_ ? _1015_ : _1018_);
	assign _1020_ = (_0254_ ? \mchip.dut.memory.M[23] [4] : \mchip.dut.memory.M[22] [4]);
	assign _1021_ = (_0254_ ? \mchip.dut.memory.M[21] [4] : \mchip.dut.memory.M[20] [4]);
	assign _1022_ = (_0259_ ? _1020_ : _1021_);
	assign _1023_ = (_0254_ ? \mchip.dut.memory.M[19] [4] : \mchip.dut.memory.M[18] [4]);
	assign _1024_ = (_0254_ ? \mchip.dut.memory.M[17] [4] : \mchip.dut.memory.M[16] [4]);
	assign _1025_ = (_0259_ ? _1023_ : _1024_);
	assign _1026_ = (_0268_ ? _1022_ : _1025_);
	assign _1027_ = (_0282_ ? _1019_ : _1026_);
	assign _1028_ = (_0254_ ? \mchip.dut.memory.M[15] [4] : \mchip.dut.memory.M[14] [4]);
	assign _1029_ = (_0254_ ? \mchip.dut.memory.M[13] [4] : \mchip.dut.memory.M[12] [4]);
	assign _1030_ = (_0259_ ? _1028_ : _1029_);
	assign _1031_ = (_0254_ ? \mchip.dut.memory.M[11] [4] : \mchip.dut.memory.M[10] [4]);
	assign _1032_ = (_0254_ ? \mchip.dut.memory.M[9] [4] : \mchip.dut.memory.M[8] [4]);
	assign _1033_ = (_0259_ ? _1031_ : _1032_);
	assign _1034_ = (_0268_ ? _1030_ : _1033_);
	assign _1035_ = (_0254_ ? \mchip.dut.memory.M[7] [4] : \mchip.dut.memory.M[6] [4]);
	assign _1036_ = (_0254_ ? \mchip.dut.memory.M[5] [4] : \mchip.dut.memory.M[4] [4]);
	assign _1037_ = (_0259_ ? _1035_ : _1036_);
	assign _1038_ = (_0254_ ? \mchip.dut.memory.M[3] [4] : \mchip.dut.memory.M[2] [4]);
	assign _1039_ = (_0254_ ? \mchip.dut.memory.M[1] [4] : \mchip.dut.memory.M[0] [4]);
	assign _1040_ = (_0259_ ? _1038_ : _1039_);
	assign _1041_ = (_0268_ ? _1037_ : _1040_);
	assign _1042_ = (_0282_ ? _1034_ : _1041_);
	assign _1043_ = (_0305_ ? _1027_ : _1042_);
	assign _1044_ = (_0342_ ? _1012_ : _1043_);
	assign \mchip.dut.demux.I [4] = (_0412_ ? _0981_ : _1044_);
	assign _1045_ = _0210_ & ~_0540_;
	assign \mchip.dut.tape_reg.D  = (\mchip.dut.direction_reg.Q [0] ? \mchip.dut.display_reg.Q [1] : _1045_);
	assign _1046_ = ~\mchip.dut.state_addr.Q [0];
	assign _0035_ = (\mchip.dut.StateAddr_ld  ? _1045_ : _1046_);
	assign _1047_ = \mchip.dut.state_addr.Q [1] ^ \mchip.dut.state_addr.Q [0];
	assign _1048_ = ~(_1045_ ^ \mchip.dut.next_state.Q [0]);
	assign _0036_ = (\mchip.dut.StateAddr_ld  ? _1048_ : _1047_);
	assign _1049_ = \mchip.dut.state_addr.Q [1] & \mchip.dut.state_addr.Q [0];
	assign _1050_ = _1049_ ^ \mchip.dut.state_addr.Q [2];
	assign _1051_ = _1045_ & ~\mchip.dut.next_state.Q [0];
	assign _1052_ = \mchip.dut.next_state.Q [1] ^ \mchip.dut.next_state.Q [0];
	assign _1053_ = _1052_ ^ \mchip.dut.next_state.Q [0];
	assign _1054_ = _1053_ ^ _1051_;
	assign _0037_ = (\mchip.dut.StateAddr_ld  ? _1054_ : _1050_);
	assign _1055_ = _1049_ & \mchip.dut.state_addr.Q [2];
	assign _1056_ = _1055_ ^ \mchip.dut.state_addr.Q [3];
	assign _1057_ = _1053_ & _1051_;
	assign _1058_ = \mchip.dut.next_state.Q [0] & ~\mchip.dut.next_state.Q [1];
	assign _1059_ = \mchip.dut.next_state.Q [1] & \mchip.dut.next_state.Q [0];
	assign _1060_ = ~(\mchip.dut.next_state.Q [2] ^ \mchip.dut.next_state.Q [1]);
	assign _1061_ = _1060_ ^ _1059_;
	assign _1062_ = _1061_ ^ _1058_;
	assign _1063_ = _1062_ ^ _1057_;
	assign _0038_ = (\mchip.dut.StateAddr_ld  ? _1063_ : _1056_);
	assign _1064_ = ~(\mchip.dut.state_addr.Q [3] & \mchip.dut.state_addr.Q [2]);
	assign _1065_ = _1049_ & ~_1064_;
	assign _1066_ = _1065_ ^ \mchip.dut.state_addr.Q [4];
	assign _1067_ = ~(_1062_ & _1053_);
	assign _1068_ = _1051_ & ~_1067_;
	assign _1069_ = _1060_ & _1059_;
	assign _1070_ = _1061_ & _1058_;
	assign _1071_ = ~(_1070_ | _1069_);
	assign _1072_ = ~(\mchip.dut.next_state.Q [2] | \mchip.dut.next_state.Q [1]);
	assign _1073_ = ~(\mchip.dut.next_state.Q [3] ^ \mchip.dut.next_state.Q [2]);
	assign _1074_ = ~(_1073_ ^ _1072_);
	assign _1075_ = ~_1074_;
	assign _1076_ = _1075_ ^ _1071_;
	assign _1077_ = _1076_ ^ _1068_;
	assign _0039_ = (\mchip.dut.StateAddr_ld  ? _1077_ : _1066_);
	assign _1078_ = _1065_ & \mchip.dut.state_addr.Q [4];
	assign _1079_ = _1078_ ^ \mchip.dut.state_addr.Q [5];
	assign _1080_ = ~_1076_;
	assign _1081_ = _1068_ & ~_1080_;
	assign _1082_ = _1073_ & ~_1072_;
	assign _1083_ = _1074_ & _1069_;
	assign _1084_ = _1083_ | _1082_;
	assign _1085_ = ~(_1074_ & _1061_);
	assign _1086_ = _1058_ & ~_1085_;
	assign _1087_ = _1086_ | _1084_;
	assign _1088_ = ~(\mchip.dut.next_state.Q [3] | \mchip.dut.next_state.Q [2]);
	assign _1089_ = ~(\mchip.dut.next_state.Q [4] ^ \mchip.dut.next_state.Q [3]);
	assign _1090_ = ~(_1089_ ^ _1088_);
	assign _1091_ = _1090_ ^ _1087_;
	assign _1092_ = _1091_ ^ _1081_;
	assign _0040_ = (\mchip.dut.StateAddr_ld  ? _1092_ : _1079_);
	assign _1093_ = ~(\mchip.dut.state_addr.Q [5] & \mchip.dut.state_addr.Q [4]);
	assign _1094_ = _1065_ & ~_1093_;
	assign _1095_ = _1094_ ^ \mchip.dut.state_addr.Q [6];
	assign _1096_ = _1091_ & ~_1080_;
	assign _1097_ = ~(_1096_ & _1068_);
	assign _1098_ = \mchip.dut.next_state.Q [4] | ~\mchip.dut.next_state.Q [3];
	assign _1099_ = _1088_ | ~_1089_;
	assign _1100_ = _1090_ & _1087_;
	assign _1101_ = _1099_ & ~_1100_;
	assign _1102_ = _1101_ ^ _1098_;
	assign _1103_ = _1102_ ^ _1097_;
	assign _0041_ = (\mchip.dut.StateAddr_ld  ? _1103_ : _1095_);
	assign _0042_ = (_0227_ ? \mchip.sync3.sync  : _1384_);
	assign _1104_ = ~(_0225_ ^ \mchip.dut.tape_addr.Q [1]);
	assign _1105_ = _1104_ ^ \mchip.dut.tape_addr.Q [0];
	assign _0043_ = (_0227_ ? \mchip.sync4.sync  : _1105_);
	assign _1106_ = \mchip.dut.tape_addr.Q [1] & ~_0225_;
	assign _1107_ = _1104_ & ~_1384_;
	assign _1108_ = _1107_ | _1106_;
	assign _1109_ = _0225_ ^ _0264_;
	assign _1110_ = _1109_ ^ _1108_;
	assign _0044_ = (_0227_ ? \mchip.sync5.sync  : _1110_);
	assign _1111_ = \mchip.dut.tape_addr.Q [2] & ~_0225_;
	assign _1112_ = _1109_ & _1108_;
	assign _1113_ = _1112_ | _1111_;
	assign _1114_ = _0225_ ^ _0277_;
	assign _1115_ = _1114_ ^ _1113_;
	assign _0045_ = (_0227_ ? \mchip.sync6.sync  : _1115_);
	assign _1116_ = \mchip.dut.tape_addr.Q [3] & ~_0225_;
	assign _1117_ = _1114_ & _1111_;
	assign _1118_ = _1117_ | _1116_;
	assign _1119_ = ~(_1114_ & _1109_);
	assign _1120_ = _1108_ & ~_1119_;
	assign _1121_ = _1120_ | _1118_;
	assign _1122_ = ~(_0225_ ^ \mchip.dut.tape_addr.Q [4]);
	assign _1123_ = _1122_ ^ _1121_;
	assign _0046_ = (_0227_ ? \mchip.sync7.sync  : _1123_);
	assign _1124_ = \mchip.dut.tape_addr.Q [4] & ~_0225_;
	assign _1125_ = _1122_ & _1121_;
	assign _1126_ = _1125_ | _1124_;
	assign _1127_ = ~(_0225_ ^ \mchip.dut.tape_addr.Q [5]);
	assign _1128_ = _1127_ ^ _1126_;
	assign _0047_ = (_0227_ ? \mchip.sync8.sync  : _1128_);
	assign _1129_ = \mchip.dut.tape_addr.Q [5] & ~_0225_;
	assign _1130_ = _1127_ & _1124_;
	assign _1131_ = _1130_ | _1129_;
	assign _1132_ = ~(_1127_ & _1122_);
	assign _1133_ = _1121_ & ~_1132_;
	assign _1134_ = _1133_ | _1131_;
	assign _1135_ = _0225_ ^ \mchip.dut.tape_addr.Q [6];
	assign _1136_ = ~(_1135_ ^ _1134_);
	assign _0048_ = _1136_ & ~_0227_;
	assign _1137_ = _0197_ & ~_0201_;
	assign \mchip.dut.demux.Y2 [0] = _1137_ & ~_0540_;
	assign _1138_ = ~\mchip.dut.display_reg.Q [0];
	assign _1139_ = \mchip.dut.tape_reg.Q  & ~\mchip.dut.direction_reg.Q [0];
	assign _1140_ = (_1355_ ? _1139_ : \mchip.dut.display_reg.Q [1]);
	assign _0024_ = (_1348_ ? _1138_ : _1140_);
	assign _0026_ = (_1355_ ? \mchip.dut.display_reg.Q [0] : \mchip.dut.display_reg.Q [2]);
	assign _0027_ = (_1355_ ? \mchip.dut.display_reg.Q [1] : \mchip.dut.display_reg.Q [3]);
	assign _0028_ = (_1355_ ? \mchip.dut.display_reg.Q [2] : \mchip.dut.display_reg.Q [4]);
	assign _0029_ = (_1355_ ? \mchip.dut.display_reg.Q [3] : \mchip.dut.display_reg.Q [5]);
	assign _0030_ = (_1355_ ? \mchip.dut.display_reg.Q [4] : \mchip.dut.display_reg.Q [6]);
	assign _0031_ = (_1355_ ? \mchip.dut.display_reg.Q [5] : \mchip.dut.display_reg.Q [7]);
	assign _0032_ = (_1355_ ? \mchip.dut.display_reg.Q [6] : \mchip.dut.display_reg.Q [8]);
	assign _0033_ = (_1355_ ? \mchip.dut.display_reg.Q [7] : \mchip.dut.display_reg.Q [9]);
	assign _0034_ = (_1355_ ? \mchip.dut.display_reg.Q [8] : \mchip.dut.display_reg.Q [10]);
	assign _0025_ = (_1355_ ? \mchip.dut.display_reg.Q [9] : _1139_);
	assign \mchip.dut.memory.data_in [0] = (_0235_ ? \mchip.sync3.sync  : \mchip.dut.data_reg.Q );
	assign \mchip.dut.memory.data_in [1] = _0235_ & \mchip.sync4.sync ;
	assign \mchip.dut.memory.data_in [2] = _0235_ & \mchip.sync5.sync ;
	assign \mchip.dut.memory.data_in [3] = _0235_ & \mchip.sync6.sync ;
	assign \mchip.dut.memory.data_in [4] = _0235_ & \mchip.sync7.sync ;
	assign _1141_ = _0198_ | \mchip.dut.fsm.currState [0];
	assign _1142_ = ~(\mchip.dut.fsm.currState [3] | \mchip.dut.fsm.currState [0]);
	assign \mchip.dut.NextState_en  = _1141_ & ~_1142_;
	assign _1143_ = _1349_ & ~_0241_;
	assign \mchip.dut.InputAddr_en  = _0250_ & ~_1143_;
	assign _1144_ = _0249_ | _1348_;
	assign _1145_ = _1144_ | _0235_;
	assign _1146_ = ~(\mchip.dut.fsm.currState [1] | \mchip.dut.fsm.currState [5]);
	assign _1147_ = ~(_0234_ & _1349_);
	assign _1148_ = _1146_ & ~_1147_;
	assign _1149_ = _1145_ & ~_1148_;
	assign _1150_ = ~(_0412_ & _0342_);
	assign _1151_ = _0305_ | _0282_;
	assign _1152_ = _1151_ | _1150_;
	assign _1153_ = ~(_0268_ & _0259_);
	assign _1154_ = _1153_ | _0254_;
	assign _1155_ = _1154_ | _1152_;
	assign _0052_ = _1149_ & ~_1155_;
	assign _1156_ = ~_0254_;
	assign _1157_ = _0259_ | ~_0268_;
	assign _1158_ = _1157_ | _1156_;
	assign _1159_ = _1158_ | _1152_;
	assign _0051_ = _1149_ & ~_1159_;
	assign _1160_ = _1153_ | _1156_;
	assign _1161_ = _1160_ | _1152_;
	assign _0053_ = _1149_ & ~_1161_;
	assign _1162_ = _0412_ | _0342_;
	assign _1163_ = _1162_ | _1151_;
	assign _1164_ = _0268_ | _0259_;
	assign _1165_ = _1164_ | _0254_;
	assign _1166_ = _1165_ | _1163_;
	assign _0049_ = _1149_ & ~_1166_;
	assign _1167_ = _1164_ | _1156_;
	assign _1168_ = _1167_ | _1163_;
	assign _0088_ = _1149_ & ~_1168_;
	assign _1169_ = _0268_ | ~_0259_;
	assign _1170_ = _1169_ | _0254_;
	assign _1171_ = _1170_ | _1163_;
	assign _0099_ = _1149_ & ~_1171_;
	assign _1172_ = _1169_ | _1156_;
	assign _1173_ = _1172_ | _1163_;
	assign _0110_ = _1149_ & ~_1173_;
	assign _1174_ = _1157_ | _0254_;
	assign _1175_ = _1174_ | _1163_;
	assign _0121_ = _1149_ & ~_1175_;
	assign _1176_ = _1163_ | _1158_;
	assign _0132_ = _1149_ & ~_1176_;
	assign _1177_ = _1163_ | _1154_;
	assign _0143_ = _1149_ & ~_1177_;
	assign _1178_ = _1163_ | _1160_;
	assign _0154_ = _1149_ & ~_1178_;
	assign _1179_ = _0305_ | ~_0282_;
	assign _1180_ = _1179_ | _1162_;
	assign _1181_ = _1180_ | _1165_;
	assign _0165_ = _1149_ & ~_1181_;
	assign _1182_ = _1180_ | _1167_;
	assign _0176_ = _1149_ & ~_1182_;
	assign _1183_ = _1180_ | _1170_;
	assign _0060_ = _1149_ & ~_1183_;
	assign _1184_ = _1180_ | _1172_;
	assign _0071_ = _1149_ & ~_1184_;
	assign _1185_ = _1180_ | _1174_;
	assign _0080_ = _1149_ & ~_1185_;
	assign _1186_ = _1180_ | _1158_;
	assign _0081_ = _1149_ & ~_1186_;
	assign _1187_ = _1180_ | _1154_;
	assign _0082_ = _1149_ & ~_1187_;
	assign _1188_ = _1180_ | _1160_;
	assign _0083_ = _1149_ & ~_1188_;
	assign _1189_ = _0282_ | ~_0305_;
	assign _1190_ = _1189_ | _1162_;
	assign _1191_ = _1190_ | _1165_;
	assign _0084_ = _1149_ & ~_1191_;
	assign _1192_ = _1190_ | _1167_;
	assign _0085_ = _1149_ & ~_1192_;
	assign _1193_ = _1190_ | _1170_;
	assign _0086_ = _1149_ & ~_1193_;
	assign _1194_ = _1190_ | _1172_;
	assign _0087_ = _1149_ & ~_1194_;
	assign _1195_ = _1190_ | _1174_;
	assign _0089_ = _1149_ & ~_1195_;
	assign _1196_ = _1190_ | _1158_;
	assign _0090_ = _1149_ & ~_1196_;
	assign _1197_ = _1190_ | _1154_;
	assign _0091_ = _1149_ & ~_1197_;
	assign _1198_ = _1190_ | _1160_;
	assign _0092_ = _1149_ & ~_1198_;
	assign _1199_ = ~(_0305_ & _0282_);
	assign _1200_ = _1199_ | _1162_;
	assign _1201_ = _1200_ | _1165_;
	assign _0093_ = _1149_ & ~_1201_;
	assign _1202_ = _1200_ | _1167_;
	assign _0094_ = _1149_ & ~_1202_;
	assign _1203_ = _1200_ | _1170_;
	assign _0095_ = _1149_ & ~_1203_;
	assign _1204_ = _1200_ | _1172_;
	assign _0096_ = _1149_ & ~_1204_;
	assign _1205_ = _1200_ | _1174_;
	assign _0097_ = _1149_ & ~_1205_;
	assign _1206_ = _1200_ | _1158_;
	assign _0098_ = _1149_ & ~_1206_;
	assign _1207_ = _1200_ | _1154_;
	assign _0100_ = _1149_ & ~_1207_;
	assign _1208_ = _1200_ | _1160_;
	assign _0101_ = _1149_ & ~_1208_;
	assign _1209_ = _0412_ | ~_0342_;
	assign _1210_ = _1209_ | _1151_;
	assign _1211_ = _1210_ | _1165_;
	assign _0102_ = _1149_ & ~_1211_;
	assign _1212_ = _1210_ | _1167_;
	assign _0103_ = _1149_ & ~_1212_;
	assign _1213_ = _1210_ | _1170_;
	assign _0104_ = _1149_ & ~_1213_;
	assign _1214_ = _1210_ | _1172_;
	assign _0105_ = _1149_ & ~_1214_;
	assign _1215_ = _1210_ | _1174_;
	assign _0106_ = _1149_ & ~_1215_;
	assign _1216_ = _1210_ | _1158_;
	assign _0107_ = _1149_ & ~_1216_;
	assign _1217_ = _1210_ | _1154_;
	assign _0108_ = _1149_ & ~_1217_;
	assign _1218_ = _1210_ | _1160_;
	assign _0109_ = _1149_ & ~_1218_;
	assign _1219_ = _1209_ | _1179_;
	assign _1220_ = _1219_ | _1165_;
	assign _0111_ = _1149_ & ~_1220_;
	assign _1221_ = _1219_ | _1167_;
	assign _0112_ = _1149_ & ~_1221_;
	assign _1222_ = _1219_ | _1170_;
	assign _0113_ = _1149_ & ~_1222_;
	assign _1223_ = _1219_ | _1172_;
	assign _0114_ = _1149_ & ~_1223_;
	assign _1224_ = _1219_ | _1174_;
	assign _0115_ = _1149_ & ~_1224_;
	assign _1225_ = _1219_ | _1158_;
	assign _0116_ = _1149_ & ~_1225_;
	assign _1226_ = _1219_ | _1154_;
	assign _0117_ = _1149_ & ~_1226_;
	assign _1227_ = _1219_ | _1160_;
	assign _0118_ = _1149_ & ~_1227_;
	assign _1228_ = _1209_ | _1189_;
	assign _1229_ = _1228_ | _1165_;
	assign _0119_ = _1149_ & ~_1229_;
	assign _1230_ = _1228_ | _1167_;
	assign _0120_ = _1149_ & ~_1230_;
	assign _1231_ = _1228_ | _1170_;
	assign _0122_ = _1149_ & ~_1231_;
	assign _1232_ = _1228_ | _1172_;
	assign _0123_ = _1149_ & ~_1232_;
	assign _1233_ = _1228_ | _1174_;
	assign _0124_ = _1149_ & ~_1233_;
	assign _1234_ = _1228_ | _1158_;
	assign _0125_ = _1149_ & ~_1234_;
	assign _1235_ = _1228_ | _1154_;
	assign _0126_ = _1149_ & ~_1235_;
	assign _1236_ = _1228_ | _1160_;
	assign _0127_ = _1149_ & ~_1236_;
	assign _1237_ = _1209_ | _1199_;
	assign _1238_ = _1237_ | _1165_;
	assign _0128_ = _1149_ & ~_1238_;
	assign _1239_ = _1237_ | _1167_;
	assign _0129_ = _1149_ & ~_1239_;
	assign _1240_ = _1237_ | _1170_;
	assign _0130_ = _1149_ & ~_1240_;
	assign _1241_ = _1237_ | _1172_;
	assign _0131_ = _1149_ & ~_1241_;
	assign _1242_ = _1237_ | _1174_;
	assign _0133_ = _1149_ & ~_1242_;
	assign _1243_ = _1237_ | _1158_;
	assign _0134_ = _1149_ & ~_1243_;
	assign _1244_ = _1237_ | _1154_;
	assign _0135_ = _1149_ & ~_1244_;
	assign _1245_ = _1237_ | _1160_;
	assign _0136_ = _1149_ & ~_1245_;
	assign _1246_ = _0342_ | ~_0412_;
	assign _1247_ = _1246_ | _1151_;
	assign _1248_ = _1247_ | _1165_;
	assign _0137_ = _1149_ & ~_1248_;
	assign _1249_ = _1247_ | _1167_;
	assign _0138_ = _1149_ & ~_1249_;
	assign _1250_ = _1247_ | _1170_;
	assign _0139_ = _1149_ & ~_1250_;
	assign _1251_ = _1247_ | _1172_;
	assign _0140_ = _1149_ & ~_1251_;
	assign _1252_ = _1247_ | _1174_;
	assign _0141_ = _1149_ & ~_1252_;
	assign _1253_ = _1247_ | _1158_;
	assign _0142_ = _1149_ & ~_1253_;
	assign _1254_ = _1247_ | _1154_;
	assign _0144_ = _1149_ & ~_1254_;
	assign _1255_ = _1247_ | _1160_;
	assign _0145_ = _1149_ & ~_1255_;
	assign _1256_ = _1246_ | _1179_;
	assign _1257_ = _1256_ | _1165_;
	assign _0146_ = _1149_ & ~_1257_;
	assign _1258_ = _1256_ | _1167_;
	assign _0147_ = _1149_ & ~_1258_;
	assign _1259_ = _1256_ | _1170_;
	assign _0148_ = _1149_ & ~_1259_;
	assign _1260_ = _1256_ | _1172_;
	assign _0149_ = _1149_ & ~_1260_;
	assign _1261_ = _1256_ | _1174_;
	assign _0150_ = _1149_ & ~_1261_;
	assign _1262_ = _1256_ | _1158_;
	assign _0151_ = _1149_ & ~_1262_;
	assign _1263_ = _1256_ | _1154_;
	assign _0152_ = _1149_ & ~_1263_;
	assign _1264_ = _1256_ | _1160_;
	assign _0153_ = _1149_ & ~_1264_;
	assign _1265_ = _1246_ | _1189_;
	assign _1266_ = _1265_ | _1165_;
	assign _0155_ = _1149_ & ~_1266_;
	assign _1267_ = _1265_ | _1167_;
	assign _0156_ = _1149_ & ~_1267_;
	assign _1268_ = _1265_ | _1170_;
	assign _0157_ = _1149_ & ~_1268_;
	assign _1269_ = _1265_ | _1172_;
	assign _0158_ = _1149_ & ~_1269_;
	assign _1270_ = _1265_ | _1174_;
	assign _0159_ = _1149_ & ~_1270_;
	assign _1271_ = _1265_ | _1158_;
	assign _0160_ = _1149_ & ~_1271_;
	assign _1272_ = _1265_ | _1154_;
	assign _0161_ = _1149_ & ~_1272_;
	assign _1273_ = _1265_ | _1160_;
	assign _0162_ = _1149_ & ~_1273_;
	assign _1274_ = _1246_ | _1199_;
	assign _1275_ = _1274_ | _1165_;
	assign _0163_ = _1149_ & ~_1275_;
	assign _1276_ = _1274_ | _1167_;
	assign _0164_ = _1149_ & ~_1276_;
	assign _1277_ = _1274_ | _1170_;
	assign _0166_ = _1149_ & ~_1277_;
	assign _1278_ = _1274_ | _1172_;
	assign _0167_ = _1149_ & ~_1278_;
	assign _1279_ = _1274_ | _1174_;
	assign _0168_ = _1149_ & ~_1279_;
	assign _1280_ = _1274_ | _1158_;
	assign _0169_ = _1149_ & ~_1280_;
	assign _1281_ = _1274_ | _1154_;
	assign _0170_ = _1149_ & ~_1281_;
	assign _1282_ = _1274_ | _1160_;
	assign _0171_ = _1149_ & ~_1282_;
	assign _1283_ = _1165_ | _1152_;
	assign _0172_ = _1149_ & ~_1283_;
	assign _1284_ = _1167_ | _1152_;
	assign _0173_ = _1149_ & ~_1284_;
	assign _1285_ = _1170_ | _1152_;
	assign _0174_ = _1149_ & ~_1285_;
	assign _1286_ = _1172_ | _1152_;
	assign _0175_ = _1149_ & ~_1286_;
	assign _1287_ = _1174_ | _1152_;
	assign _0050_ = _1149_ & ~_1287_;
	assign _1288_ = _1179_ | _1150_;
	assign _1289_ = _1288_ | _1165_;
	assign _0054_ = _1149_ & ~_1289_;
	assign _1290_ = _1288_ | _1167_;
	assign _0055_ = _1149_ & ~_1290_;
	assign _1291_ = _1288_ | _1170_;
	assign _0056_ = _1149_ & ~_1291_;
	assign _1292_ = _1288_ | _1172_;
	assign _0057_ = _1149_ & ~_1292_;
	assign _1293_ = _1288_ | _1174_;
	assign _0058_ = _1149_ & ~_1293_;
	assign _1294_ = _1288_ | _1158_;
	assign _0059_ = _1149_ & ~_1294_;
	assign _1295_ = _1288_ | _1154_;
	assign _0061_ = _1149_ & ~_1295_;
	assign _1296_ = _1288_ | _1160_;
	assign _0062_ = _1149_ & ~_1296_;
	assign _1297_ = _1189_ | _1150_;
	assign _1298_ = _1297_ | _1165_;
	assign _0063_ = _1149_ & ~_1298_;
	assign _1299_ = _1297_ | _1167_;
	assign _0064_ = _1149_ & ~_1299_;
	assign _1300_ = _1297_ | _1170_;
	assign _0065_ = _1149_ & ~_1300_;
	assign _1301_ = _1297_ | _1172_;
	assign _0066_ = _1149_ & ~_1301_;
	assign _1302_ = _1297_ | _1174_;
	assign _0067_ = _1149_ & ~_1302_;
	assign _1303_ = _1297_ | _1158_;
	assign _0068_ = _1149_ & ~_1303_;
	assign _1304_ = _1297_ | _1154_;
	assign _0069_ = _1149_ & ~_1304_;
	assign _1305_ = _1297_ | _1160_;
	assign _0070_ = _1149_ & ~_1305_;
	assign _1306_ = _1199_ | _1150_;
	assign _1307_ = _1306_ | _1165_;
	assign _0072_ = _1149_ & ~_1307_;
	assign _1308_ = _1306_ | _1167_;
	assign _0073_ = _1149_ & ~_1308_;
	assign _1309_ = _1306_ | _1170_;
	assign _0074_ = _1149_ & ~_1309_;
	assign _1310_ = _1306_ | _1172_;
	assign _0075_ = _1149_ & ~_1310_;
	assign _1311_ = _1306_ | _1174_;
	assign _0076_ = _1149_ & ~_1311_;
	assign _1312_ = _1306_ | _1158_;
	assign _0077_ = _1149_ & ~_1312_;
	assign _1313_ = _1306_ | _1154_;
	assign _0078_ = _1149_ & ~_1313_;
	assign _1314_ = _1306_ | _1160_;
	assign _0079_ = _1149_ & ~_1314_;
	assign _1315_ = ~(\mchip.dut.fsm.currState [14] | \mchip.dut.fsm.currState [6]);
	assign _0004_ = _1350_ & ~_1315_;
	assign _1316_ = io_in[13] | ~_1340_;
	assign _1317_ = _1316_ | _1339_;
	assign _0003_ = \mchip.dut.fsm.currState [5] & ~_1317_;
	assign _1318_ = ~(\mchip.dut.fsm.currState [12] | \mchip.dut.fsm.currState [4]);
	assign _0002_ = _1350_ & ~_1318_;
	assign _0001_ = _1412_ & ~_0216_;
	assign _1319_ = ~(\mchip.dut.fsm.currState [8] | \mchip.dut.fsm.currState [0]);
	assign _0000_ = _1350_ & ~_1319_;
	assign \mchip.dut.Compute_done  = _1397_ | \mchip.dut.direction_reg.Q [1];
	assign _1320_ = _1403_ & \mchip.dut.input_addr.Q [2];
	assign _1416_[3] = _1320_ ^ \mchip.dut.input_addr.Q [3];
	assign _1416_[4] = ~(_1405_ ^ \mchip.dut.input_addr.Q [4]);
	assign _1321_ = \mchip.dut.input_addr.Q [4] & ~_1405_;
	assign _1416_[5] = _1321_ ^ \mchip.dut.input_addr.Q [5];
	assign _1416_[6] = _1407_ ^ \mchip.dut.input_addr.Q [6];
	assign _1416_[1] = \mchip.dut.input_addr.Q [1] ^ \mchip.dut.input_addr.Q [0];
	assign _1416_[2] = _1403_ ^ \mchip.dut.input_addr.Q [2];
	assign _1322_ = \mchip.sync4.sync  & \mchip.sync3.sync ;
	assign _1323_ = \mchip.sync5.sync  ^ \mchip.sync4.sync ;
	assign \mchip.dut.tape_addr_min.D [3] = _1323_ ^ _1322_;
	assign _1324_ = \mchip.sync5.sync  & \mchip.sync4.sync ;
	assign _1325_ = _1323_ & _1322_;
	assign _1326_ = _1325_ | _1324_;
	assign _1327_ = \mchip.sync6.sync  ^ \mchip.sync5.sync ;
	assign \mchip.dut.tape_addr_min.D [4] = _1327_ ^ _1326_;
	assign _1328_ = \mchip.sync6.sync  & \mchip.sync5.sync ;
	assign _1329_ = _1327_ & _1324_;
	assign _1330_ = _1329_ | _1328_;
	assign _1331_ = ~(_1327_ & _1323_);
	assign _1332_ = _1322_ & ~_1331_;
	assign _1333_ = _1332_ | _1330_;
	assign _1334_ = \mchip.sync7.sync  ^ \mchip.sync6.sync ;
	assign \mchip.dut.tape_addr_min.D [5] = _1334_ ^ _1333_;
	assign _1335_ = \mchip.sync7.sync  & \mchip.sync6.sync ;
	assign _1336_ = _1334_ & _1333_;
	assign _1337_ = _1336_ | _1335_;
	assign _1338_ = \mchip.sync8.sync  ^ \mchip.sync7.sync ;
	assign \mchip.dut.tape_addr_min.D [6] = _1338_ ^ _1337_;
	assign \mchip.dut.tape_addr_min.D [2] = \mchip.sync4.sync  ^ \mchip.sync3.sync ;
	reg \mchip.dut.tape_addr_min.Q_reg[1] ;
	always @(posedge io_in[12])
		if (\mchip.dut.fsm.currState [0])
			\mchip.dut.tape_addr_min.Q_reg[1]  <= \mchip.sync3.sync ;
	assign \mchip.dut.tape_addr_min.Q [1] = \mchip.dut.tape_addr_min.Q_reg[1] ;
	reg \mchip.dut.tape_addr_min.Q_reg[2] ;
	always @(posedge io_in[12])
		if (\mchip.dut.fsm.currState [0])
			\mchip.dut.tape_addr_min.Q_reg[2]  <= \mchip.dut.tape_addr_min.D [2];
	assign \mchip.dut.tape_addr_min.Q [2] = \mchip.dut.tape_addr_min.Q_reg[2] ;
	reg \mchip.dut.tape_addr_min.Q_reg[3] ;
	always @(posedge io_in[12])
		if (\mchip.dut.fsm.currState [0])
			\mchip.dut.tape_addr_min.Q_reg[3]  <= \mchip.dut.tape_addr_min.D [3];
	assign \mchip.dut.tape_addr_min.Q [3] = \mchip.dut.tape_addr_min.Q_reg[3] ;
	reg \mchip.dut.tape_addr_min.Q_reg[4] ;
	always @(posedge io_in[12])
		if (\mchip.dut.fsm.currState [0])
			\mchip.dut.tape_addr_min.Q_reg[4]  <= \mchip.dut.tape_addr_min.D [4];
	assign \mchip.dut.tape_addr_min.Q [4] = \mchip.dut.tape_addr_min.Q_reg[4] ;
	reg \mchip.dut.tape_addr_min.Q_reg[5] ;
	always @(posedge io_in[12])
		if (\mchip.dut.fsm.currState [0])
			\mchip.dut.tape_addr_min.Q_reg[5]  <= \mchip.dut.tape_addr_min.D [5];
	assign \mchip.dut.tape_addr_min.Q [5] = \mchip.dut.tape_addr_min.Q_reg[5] ;
	reg \mchip.dut.tape_addr_min.Q_reg[6] ;
	always @(posedge io_in[12])
		if (\mchip.dut.fsm.currState [0])
			\mchip.dut.tape_addr_min.Q_reg[6]  <= \mchip.dut.tape_addr_min.D [6];
	assign \mchip.dut.tape_addr_min.Q [6] = \mchip.dut.tape_addr_min.Q_reg[6] ;
	always @(posedge io_in[12])
		if (_0082_)
			\mchip.dut.memory.M[14] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0082_)
			\mchip.dut.memory.M[14] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0082_)
			\mchip.dut.memory.M[14] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0082_)
			\mchip.dut.memory.M[14] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0082_)
			\mchip.dut.memory.M[14] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0081_)
			\mchip.dut.memory.M[13] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0081_)
			\mchip.dut.memory.M[13] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0081_)
			\mchip.dut.memory.M[13] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0081_)
			\mchip.dut.memory.M[13] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0081_)
			\mchip.dut.memory.M[13] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0118_)
			\mchip.dut.memory.M[47] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0118_)
			\mchip.dut.memory.M[47] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0118_)
			\mchip.dut.memory.M[47] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0118_)
			\mchip.dut.memory.M[47] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0118_)
			\mchip.dut.memory.M[47] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0117_)
			\mchip.dut.memory.M[46] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0117_)
			\mchip.dut.memory.M[46] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0117_)
			\mchip.dut.memory.M[46] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0117_)
			\mchip.dut.memory.M[46] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0117_)
			\mchip.dut.memory.M[46] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0116_)
			\mchip.dut.memory.M[45] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0116_)
			\mchip.dut.memory.M[45] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0116_)
			\mchip.dut.memory.M[45] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0116_)
			\mchip.dut.memory.M[45] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0116_)
			\mchip.dut.memory.M[45] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0115_)
			\mchip.dut.memory.M[44] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0115_)
			\mchip.dut.memory.M[44] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0115_)
			\mchip.dut.memory.M[44] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0115_)
			\mchip.dut.memory.M[44] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0115_)
			\mchip.dut.memory.M[44] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0114_)
			\mchip.dut.memory.M[43] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0114_)
			\mchip.dut.memory.M[43] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0114_)
			\mchip.dut.memory.M[43] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0114_)
			\mchip.dut.memory.M[43] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0114_)
			\mchip.dut.memory.M[43] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0113_)
			\mchip.dut.memory.M[42] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0113_)
			\mchip.dut.memory.M[42] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0113_)
			\mchip.dut.memory.M[42] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0113_)
			\mchip.dut.memory.M[42] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0113_)
			\mchip.dut.memory.M[42] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0112_)
			\mchip.dut.memory.M[41] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0112_)
			\mchip.dut.memory.M[41] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0112_)
			\mchip.dut.memory.M[41] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0112_)
			\mchip.dut.memory.M[41] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0112_)
			\mchip.dut.memory.M[41] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0111_)
			\mchip.dut.memory.M[40] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0111_)
			\mchip.dut.memory.M[40] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0111_)
			\mchip.dut.memory.M[40] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0111_)
			\mchip.dut.memory.M[40] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0111_)
			\mchip.dut.memory.M[40] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0110_)
			\mchip.dut.memory.M[3] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0110_)
			\mchip.dut.memory.M[3] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0110_)
			\mchip.dut.memory.M[3] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0110_)
			\mchip.dut.memory.M[3] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0110_)
			\mchip.dut.memory.M[3] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0108_)
			\mchip.dut.memory.M[38] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0108_)
			\mchip.dut.memory.M[38] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0108_)
			\mchip.dut.memory.M[38] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0108_)
			\mchip.dut.memory.M[38] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0108_)
			\mchip.dut.memory.M[38] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0107_)
			\mchip.dut.memory.M[37] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0107_)
			\mchip.dut.memory.M[37] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0107_)
			\mchip.dut.memory.M[37] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0107_)
			\mchip.dut.memory.M[37] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0107_)
			\mchip.dut.memory.M[37] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0106_)
			\mchip.dut.memory.M[36] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0106_)
			\mchip.dut.memory.M[36] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0106_)
			\mchip.dut.memory.M[36] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0106_)
			\mchip.dut.memory.M[36] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0106_)
			\mchip.dut.memory.M[36] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0105_)
			\mchip.dut.memory.M[35] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0105_)
			\mchip.dut.memory.M[35] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0105_)
			\mchip.dut.memory.M[35] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0105_)
			\mchip.dut.memory.M[35] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0105_)
			\mchip.dut.memory.M[35] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0104_)
			\mchip.dut.memory.M[34] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0104_)
			\mchip.dut.memory.M[34] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0104_)
			\mchip.dut.memory.M[34] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0104_)
			\mchip.dut.memory.M[34] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0104_)
			\mchip.dut.memory.M[34] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0103_)
			\mchip.dut.memory.M[33] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0103_)
			\mchip.dut.memory.M[33] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0103_)
			\mchip.dut.memory.M[33] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0103_)
			\mchip.dut.memory.M[33] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0103_)
			\mchip.dut.memory.M[33] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0102_)
			\mchip.dut.memory.M[32] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0102_)
			\mchip.dut.memory.M[32] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0102_)
			\mchip.dut.memory.M[32] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0102_)
			\mchip.dut.memory.M[32] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0102_)
			\mchip.dut.memory.M[32] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0101_)
			\mchip.dut.memory.M[31] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0101_)
			\mchip.dut.memory.M[31] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0101_)
			\mchip.dut.memory.M[31] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0101_)
			\mchip.dut.memory.M[31] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0101_)
			\mchip.dut.memory.M[31] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0100_)
			\mchip.dut.memory.M[30] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0100_)
			\mchip.dut.memory.M[30] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0100_)
			\mchip.dut.memory.M[30] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0100_)
			\mchip.dut.memory.M[30] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0100_)
			\mchip.dut.memory.M[30] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0099_)
			\mchip.dut.memory.M[2] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0099_)
			\mchip.dut.memory.M[2] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0099_)
			\mchip.dut.memory.M[2] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0099_)
			\mchip.dut.memory.M[2] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0099_)
			\mchip.dut.memory.M[2] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0097_)
			\mchip.dut.memory.M[28] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0097_)
			\mchip.dut.memory.M[28] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0097_)
			\mchip.dut.memory.M[28] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0097_)
			\mchip.dut.memory.M[28] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0097_)
			\mchip.dut.memory.M[28] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0096_)
			\mchip.dut.memory.M[27] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0096_)
			\mchip.dut.memory.M[27] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0096_)
			\mchip.dut.memory.M[27] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0096_)
			\mchip.dut.memory.M[27] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0096_)
			\mchip.dut.memory.M[27] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0095_)
			\mchip.dut.memory.M[26] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0095_)
			\mchip.dut.memory.M[26] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0095_)
			\mchip.dut.memory.M[26] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0095_)
			\mchip.dut.memory.M[26] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0095_)
			\mchip.dut.memory.M[26] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0094_)
			\mchip.dut.memory.M[25] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0094_)
			\mchip.dut.memory.M[25] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0094_)
			\mchip.dut.memory.M[25] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0094_)
			\mchip.dut.memory.M[25] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0094_)
			\mchip.dut.memory.M[25] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0093_)
			\mchip.dut.memory.M[24] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0093_)
			\mchip.dut.memory.M[24] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0093_)
			\mchip.dut.memory.M[24] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0093_)
			\mchip.dut.memory.M[24] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0093_)
			\mchip.dut.memory.M[24] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0092_)
			\mchip.dut.memory.M[23] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0092_)
			\mchip.dut.memory.M[23] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0092_)
			\mchip.dut.memory.M[23] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0092_)
			\mchip.dut.memory.M[23] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0092_)
			\mchip.dut.memory.M[23] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0091_)
			\mchip.dut.memory.M[22] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0091_)
			\mchip.dut.memory.M[22] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0091_)
			\mchip.dut.memory.M[22] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0091_)
			\mchip.dut.memory.M[22] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0091_)
			\mchip.dut.memory.M[22] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0090_)
			\mchip.dut.memory.M[21] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0090_)
			\mchip.dut.memory.M[21] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0090_)
			\mchip.dut.memory.M[21] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0090_)
			\mchip.dut.memory.M[21] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0090_)
			\mchip.dut.memory.M[21] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0089_)
			\mchip.dut.memory.M[20] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0089_)
			\mchip.dut.memory.M[20] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0089_)
			\mchip.dut.memory.M[20] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0089_)
			\mchip.dut.memory.M[20] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0089_)
			\mchip.dut.memory.M[20] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0088_)
			\mchip.dut.memory.M[1] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0088_)
			\mchip.dut.memory.M[1] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0088_)
			\mchip.dut.memory.M[1] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0088_)
			\mchip.dut.memory.M[1] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0088_)
			\mchip.dut.memory.M[1] [4] <= \mchip.dut.memory.data_in [4];
	reg \mchip.dut.next_state.Q_reg[1] ;
	always @(posedge io_in[12])
		if (\mchip.dut.NextState_en )
			if (_0023_)
				\mchip.dut.next_state.Q_reg[1]  <= 1'h0;
			else
				\mchip.dut.next_state.Q_reg[1]  <= \mchip.dut.demux.I [1];
	assign \mchip.dut.next_state.Q [1] = \mchip.dut.next_state.Q_reg[1] ;
	reg \mchip.dut.next_state.Q_reg[2] ;
	always @(posedge io_in[12])
		if (\mchip.dut.NextState_en )
			if (_0023_)
				\mchip.dut.next_state.Q_reg[2]  <= 1'h0;
			else
				\mchip.dut.next_state.Q_reg[2]  <= \mchip.dut.demux.I [2];
	assign \mchip.dut.next_state.Q [2] = \mchip.dut.next_state.Q_reg[2] ;
	reg \mchip.dut.next_state.Q_reg[3] ;
	always @(posedge io_in[12])
		if (\mchip.dut.NextState_en )
			if (_0023_)
				\mchip.dut.next_state.Q_reg[3]  <= 1'h0;
			else
				\mchip.dut.next_state.Q_reg[3]  <= \mchip.dut.demux.I [3];
	assign \mchip.dut.next_state.Q [3] = \mchip.dut.next_state.Q_reg[3] ;
	reg \mchip.dut.next_state.Q_reg[4] ;
	always @(posedge io_in[12])
		if (\mchip.dut.NextState_en )
			if (_0023_)
				\mchip.dut.next_state.Q_reg[4]  <= 1'h0;
			else
				\mchip.dut.next_state.Q_reg[4]  <= \mchip.dut.demux.I [4];
	assign \mchip.dut.next_state.Q [4] = \mchip.dut.next_state.Q_reg[4] ;
	always @(posedge io_in[12])
		if (\mchip.dut.fsm.currState [0])
			\mchip.dut.display_reg.Q [1] <= 1'h0;
		else if (_0020_)
			\mchip.dut.display_reg.Q [1] <= _0026_;
	always @(posedge io_in[12])
		if (\mchip.dut.fsm.currState [0])
			\mchip.dut.display_reg.Q [2] <= 1'h0;
		else if (_0020_)
			\mchip.dut.display_reg.Q [2] <= _0027_;
	always @(posedge io_in[12])
		if (\mchip.dut.fsm.currState [0])
			\mchip.dut.display_reg.Q [3] <= 1'h0;
		else if (_0020_)
			\mchip.dut.display_reg.Q [3] <= _0028_;
	always @(posedge io_in[12])
		if (\mchip.dut.fsm.currState [0])
			\mchip.dut.display_reg.Q [4] <= 1'h0;
		else if (_0020_)
			\mchip.dut.display_reg.Q [4] <= _0029_;
	always @(posedge io_in[12])
		if (\mchip.dut.fsm.currState [0])
			\mchip.dut.display_reg.Q [5] <= 1'h0;
		else if (_0020_)
			\mchip.dut.display_reg.Q [5] <= _0030_;
	always @(posedge io_in[12])
		if (\mchip.dut.fsm.currState [0])
			\mchip.dut.display_reg.Q [6] <= 1'h0;
		else if (_0020_)
			\mchip.dut.display_reg.Q [6] <= _0031_;
	always @(posedge io_in[12])
		if (\mchip.dut.fsm.currState [0])
			\mchip.dut.display_reg.Q [7] <= 1'h0;
		else if (_0020_)
			\mchip.dut.display_reg.Q [7] <= _0032_;
	always @(posedge io_in[12])
		if (\mchip.dut.fsm.currState [0])
			\mchip.dut.display_reg.Q [8] <= 1'h0;
		else if (_0020_)
			\mchip.dut.display_reg.Q [8] <= _0033_;
	always @(posedge io_in[12])
		if (\mchip.dut.fsm.currState [0])
			\mchip.dut.display_reg.Q [9] <= 1'h0;
		else if (_0020_)
			\mchip.dut.display_reg.Q [9] <= _0034_;
	always @(posedge io_in[12])
		if (\mchip.dut.fsm.currState [0])
			\mchip.dut.display_reg.Q [10] <= 1'h0;
		else if (_0020_)
			\mchip.dut.display_reg.Q [10] <= _0025_;
	always @(posedge io_in[12])
		if (_0083_)
			\mchip.dut.memory.M[15] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0083_)
			\mchip.dut.memory.M[15] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0083_)
			\mchip.dut.memory.M[15] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0083_)
			\mchip.dut.memory.M[15] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0083_)
			\mchip.dut.memory.M[15] [4] <= \mchip.dut.memory.data_in [4];
	reg \mchip.dut.fsm.currState_reg[0] ;
	always @(posedge io_in[12]) \mchip.dut.fsm.currState_reg[0]  <= _0005_;
	assign \mchip.dut.fsm.currState [0] = \mchip.dut.fsm.currState_reg[0] ;
	reg \mchip.dut.fsm.currState_reg[1] ;
	always @(posedge io_in[12]) \mchip.dut.fsm.currState_reg[1]  <= _0007_;
	assign \mchip.dut.fsm.currState [1] = \mchip.dut.fsm.currState_reg[1] ;
	reg \mchip.dut.fsm.currState_reg[2] ;
	always @(posedge io_in[12]) \mchip.dut.fsm.currState_reg[2]  <= _0008_;
	assign \mchip.dut.fsm.currState [2] = \mchip.dut.fsm.currState_reg[2] ;
	reg \mchip.dut.fsm.currState_reg[3] ;
	always @(posedge io_in[12]) \mchip.dut.fsm.currState_reg[3]  <= _0009_;
	assign \mchip.dut.fsm.currState [3] = \mchip.dut.fsm.currState_reg[3] ;
	reg \mchip.dut.fsm.currState_reg[4] ;
	always @(posedge io_in[12]) \mchip.dut.fsm.currState_reg[4]  <= _0010_;
	assign \mchip.dut.fsm.currState [4] = \mchip.dut.fsm.currState_reg[4] ;
	reg \mchip.dut.fsm.currState_reg[5] ;
	always @(posedge io_in[12]) \mchip.dut.fsm.currState_reg[5]  <= _0011_;
	assign \mchip.dut.fsm.currState [5] = \mchip.dut.fsm.currState_reg[5] ;
	reg \mchip.dut.fsm.currState_reg[6] ;
	always @(posedge io_in[12]) \mchip.dut.fsm.currState_reg[6]  <= _0012_;
	assign \mchip.dut.fsm.currState [6] = \mchip.dut.fsm.currState_reg[6] ;
	reg \mchip.dut.fsm.currState_reg[8] ;
	always @(posedge io_in[12]) \mchip.dut.fsm.currState_reg[8]  <= _0000_;
	assign \mchip.dut.fsm.currState [8] = \mchip.dut.fsm.currState_reg[8] ;
	reg \mchip.dut.fsm.currState_reg[9] ;
	always @(posedge io_in[12]) \mchip.dut.fsm.currState_reg[9]  <= _0013_;
	assign \mchip.dut.fsm.currState [9] = \mchip.dut.fsm.currState_reg[9] ;
	reg \mchip.dut.fsm.currState_reg[10] ;
	always @(posedge io_in[12]) \mchip.dut.fsm.currState_reg[10]  <= _0006_;
	assign \mchip.dut.fsm.currState [10] = \mchip.dut.fsm.currState_reg[10] ;
	reg \mchip.dut.fsm.currState_reg[11] ;
	always @(posedge io_in[12]) \mchip.dut.fsm.currState_reg[11]  <= _0001_;
	assign \mchip.dut.fsm.currState [11] = \mchip.dut.fsm.currState_reg[11] ;
	reg \mchip.dut.fsm.currState_reg[12] ;
	always @(posedge io_in[12]) \mchip.dut.fsm.currState_reg[12]  <= _0002_;
	assign \mchip.dut.fsm.currState [12] = \mchip.dut.fsm.currState_reg[12] ;
	reg \mchip.dut.fsm.currState_reg[13] ;
	always @(posedge io_in[12]) \mchip.dut.fsm.currState_reg[13]  <= _0003_;
	assign \mchip.dut.fsm.currState [13] = \mchip.dut.fsm.currState_reg[13] ;
	reg \mchip.dut.fsm.currState_reg[14] ;
	always @(posedge io_in[12]) \mchip.dut.fsm.currState_reg[14]  <= _0004_;
	assign \mchip.dut.fsm.currState [14] = \mchip.dut.fsm.currState_reg[14] ;
	always @(posedge io_in[12])
		if (_0120_)
			\mchip.dut.memory.M[49] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0120_)
			\mchip.dut.memory.M[49] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0120_)
			\mchip.dut.memory.M[49] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0120_)
			\mchip.dut.memory.M[49] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0120_)
			\mchip.dut.memory.M[49] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0078_)
			\mchip.dut.memory.M[126] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0078_)
			\mchip.dut.memory.M[126] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0078_)
			\mchip.dut.memory.M[126] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0078_)
			\mchip.dut.memory.M[126] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0078_)
			\mchip.dut.memory.M[126] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0077_)
			\mchip.dut.memory.M[125] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0077_)
			\mchip.dut.memory.M[125] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0077_)
			\mchip.dut.memory.M[125] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0077_)
			\mchip.dut.memory.M[125] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0077_)
			\mchip.dut.memory.M[125] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0131_)
			\mchip.dut.memory.M[59] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0131_)
			\mchip.dut.memory.M[59] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0131_)
			\mchip.dut.memory.M[59] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0131_)
			\mchip.dut.memory.M[59] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0131_)
			\mchip.dut.memory.M[59] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0076_)
			\mchip.dut.memory.M[124] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0076_)
			\mchip.dut.memory.M[124] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0076_)
			\mchip.dut.memory.M[124] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0076_)
			\mchip.dut.memory.M[124] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0076_)
			\mchip.dut.memory.M[124] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0075_)
			\mchip.dut.memory.M[123] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0075_)
			\mchip.dut.memory.M[123] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0075_)
			\mchip.dut.memory.M[123] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0075_)
			\mchip.dut.memory.M[123] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0075_)
			\mchip.dut.memory.M[123] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0074_)
			\mchip.dut.memory.M[122] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0074_)
			\mchip.dut.memory.M[122] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0074_)
			\mchip.dut.memory.M[122] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0074_)
			\mchip.dut.memory.M[122] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0074_)
			\mchip.dut.memory.M[122] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0073_)
			\mchip.dut.memory.M[121] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0073_)
			\mchip.dut.memory.M[121] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0073_)
			\mchip.dut.memory.M[121] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0073_)
			\mchip.dut.memory.M[121] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0073_)
			\mchip.dut.memory.M[121] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0072_)
			\mchip.dut.memory.M[120] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0072_)
			\mchip.dut.memory.M[120] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0072_)
			\mchip.dut.memory.M[120] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0072_)
			\mchip.dut.memory.M[120] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0072_)
			\mchip.dut.memory.M[120] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0071_)
			\mchip.dut.memory.M[11] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0071_)
			\mchip.dut.memory.M[11] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0071_)
			\mchip.dut.memory.M[11] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0071_)
			\mchip.dut.memory.M[11] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0071_)
			\mchip.dut.memory.M[11] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0153_)
			\mchip.dut.memory.M[79] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0153_)
			\mchip.dut.memory.M[79] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0153_)
			\mchip.dut.memory.M[79] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0153_)
			\mchip.dut.memory.M[79] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0153_)
			\mchip.dut.memory.M[79] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0069_)
			\mchip.dut.memory.M[118] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0069_)
			\mchip.dut.memory.M[118] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0069_)
			\mchip.dut.memory.M[118] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0069_)
			\mchip.dut.memory.M[118] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0069_)
			\mchip.dut.memory.M[118] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0068_)
			\mchip.dut.memory.M[117] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0068_)
			\mchip.dut.memory.M[117] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0068_)
			\mchip.dut.memory.M[117] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0068_)
			\mchip.dut.memory.M[117] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0068_)
			\mchip.dut.memory.M[117] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0142_)
			\mchip.dut.memory.M[69] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0142_)
			\mchip.dut.memory.M[69] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0142_)
			\mchip.dut.memory.M[69] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0142_)
			\mchip.dut.memory.M[69] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0142_)
			\mchip.dut.memory.M[69] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0067_)
			\mchip.dut.memory.M[116] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0067_)
			\mchip.dut.memory.M[116] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0067_)
			\mchip.dut.memory.M[116] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0067_)
			\mchip.dut.memory.M[116] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0067_)
			\mchip.dut.memory.M[116] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0080_)
			\mchip.dut.memory.M[12] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0080_)
			\mchip.dut.memory.M[12] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0080_)
			\mchip.dut.memory.M[12] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0080_)
			\mchip.dut.memory.M[12] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0080_)
			\mchip.dut.memory.M[12] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0066_)
			\mchip.dut.memory.M[115] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0066_)
			\mchip.dut.memory.M[115] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0066_)
			\mchip.dut.memory.M[115] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0066_)
			\mchip.dut.memory.M[115] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0066_)
			\mchip.dut.memory.M[115] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0065_)
			\mchip.dut.memory.M[114] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0065_)
			\mchip.dut.memory.M[114] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0065_)
			\mchip.dut.memory.M[114] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0065_)
			\mchip.dut.memory.M[114] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0065_)
			\mchip.dut.memory.M[114] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0109_)
			\mchip.dut.memory.M[39] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0109_)
			\mchip.dut.memory.M[39] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0109_)
			\mchip.dut.memory.M[39] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0109_)
			\mchip.dut.memory.M[39] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0109_)
			\mchip.dut.memory.M[39] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0064_)
			\mchip.dut.memory.M[113] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0064_)
			\mchip.dut.memory.M[113] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0064_)
			\mchip.dut.memory.M[113] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0064_)
			\mchip.dut.memory.M[113] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0064_)
			\mchip.dut.memory.M[113] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0063_)
			\mchip.dut.memory.M[112] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0063_)
			\mchip.dut.memory.M[112] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0063_)
			\mchip.dut.memory.M[112] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0063_)
			\mchip.dut.memory.M[112] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0063_)
			\mchip.dut.memory.M[112] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0062_)
			\mchip.dut.memory.M[111] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0062_)
			\mchip.dut.memory.M[111] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0062_)
			\mchip.dut.memory.M[111] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0062_)
			\mchip.dut.memory.M[111] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0062_)
			\mchip.dut.memory.M[111] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0061_)
			\mchip.dut.memory.M[110] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0061_)
			\mchip.dut.memory.M[110] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0061_)
			\mchip.dut.memory.M[110] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0061_)
			\mchip.dut.memory.M[110] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0061_)
			\mchip.dut.memory.M[110] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0060_)
			\mchip.dut.memory.M[10] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0060_)
			\mchip.dut.memory.M[10] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0060_)
			\mchip.dut.memory.M[10] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0060_)
			\mchip.dut.memory.M[10] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0060_)
			\mchip.dut.memory.M[10] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0058_)
			\mchip.dut.memory.M[108] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0058_)
			\mchip.dut.memory.M[108] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0058_)
			\mchip.dut.memory.M[108] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0058_)
			\mchip.dut.memory.M[108] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0058_)
			\mchip.dut.memory.M[108] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0085_)
			\mchip.dut.memory.M[17] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0085_)
			\mchip.dut.memory.M[17] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0085_)
			\mchip.dut.memory.M[17] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0085_)
			\mchip.dut.memory.M[17] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0085_)
			\mchip.dut.memory.M[17] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0084_)
			\mchip.dut.memory.M[16] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0084_)
			\mchip.dut.memory.M[16] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0084_)
			\mchip.dut.memory.M[16] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0084_)
			\mchip.dut.memory.M[16] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0084_)
			\mchip.dut.memory.M[16] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0079_)
			\mchip.dut.memory.M[127] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0079_)
			\mchip.dut.memory.M[127] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0079_)
			\mchip.dut.memory.M[127] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0079_)
			\mchip.dut.memory.M[127] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0079_)
			\mchip.dut.memory.M[127] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0098_)
			\mchip.dut.memory.M[29] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0098_)
			\mchip.dut.memory.M[29] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0098_)
			\mchip.dut.memory.M[29] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0098_)
			\mchip.dut.memory.M[29] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0098_)
			\mchip.dut.memory.M[29] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0057_)
			\mchip.dut.memory.M[107] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0057_)
			\mchip.dut.memory.M[107] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0057_)
			\mchip.dut.memory.M[107] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0057_)
			\mchip.dut.memory.M[107] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0057_)
			\mchip.dut.memory.M[107] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (\mchip.dut.fsm.currState [0])
			\mchip.dut.input_addr.Q [0] <= 1'h0;
		else if (\mchip.dut.InputAddr_en )
			\mchip.dut.input_addr.Q [0] <= _1416_[0];
	always @(posedge io_in[12])
		if (\mchip.dut.fsm.currState [0])
			\mchip.dut.input_addr.Q [1] <= 1'h0;
		else if (\mchip.dut.InputAddr_en )
			\mchip.dut.input_addr.Q [1] <= _1416_[1];
	always @(posedge io_in[12])
		if (\mchip.dut.fsm.currState [0])
			\mchip.dut.input_addr.Q [2] <= 1'h0;
		else if (\mchip.dut.InputAddr_en )
			\mchip.dut.input_addr.Q [2] <= _1416_[2];
	always @(posedge io_in[12])
		if (\mchip.dut.fsm.currState [0])
			\mchip.dut.input_addr.Q [3] <= 1'h0;
		else if (\mchip.dut.InputAddr_en )
			\mchip.dut.input_addr.Q [3] <= _1416_[3];
	always @(posedge io_in[12])
		if (\mchip.dut.fsm.currState [0])
			\mchip.dut.input_addr.Q [4] <= 1'h0;
		else if (\mchip.dut.InputAddr_en )
			\mchip.dut.input_addr.Q [4] <= _1416_[4];
	always @(posedge io_in[12])
		if (\mchip.dut.fsm.currState [0])
			\mchip.dut.input_addr.Q [5] <= 1'h0;
		else if (\mchip.dut.InputAddr_en )
			\mchip.dut.input_addr.Q [5] <= _1416_[5];
	always @(posedge io_in[12])
		if (\mchip.dut.fsm.currState [0])
			\mchip.dut.input_addr.Q [6] <= 1'h0;
		else if (\mchip.dut.InputAddr_en )
			\mchip.dut.input_addr.Q [6] <= _1416_[6];
	always @(posedge io_in[12])
		if (_0146_)
			\mchip.dut.memory.M[72] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0146_)
			\mchip.dut.memory.M[72] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0146_)
			\mchip.dut.memory.M[72] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0146_)
			\mchip.dut.memory.M[72] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0146_)
			\mchip.dut.memory.M[72] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0147_)
			\mchip.dut.memory.M[73] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0147_)
			\mchip.dut.memory.M[73] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0147_)
			\mchip.dut.memory.M[73] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0147_)
			\mchip.dut.memory.M[73] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0147_)
			\mchip.dut.memory.M[73] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0148_)
			\mchip.dut.memory.M[74] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0148_)
			\mchip.dut.memory.M[74] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0148_)
			\mchip.dut.memory.M[74] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0148_)
			\mchip.dut.memory.M[74] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0148_)
			\mchip.dut.memory.M[74] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0149_)
			\mchip.dut.memory.M[75] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0149_)
			\mchip.dut.memory.M[75] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0149_)
			\mchip.dut.memory.M[75] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0149_)
			\mchip.dut.memory.M[75] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0149_)
			\mchip.dut.memory.M[75] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0150_)
			\mchip.dut.memory.M[76] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0150_)
			\mchip.dut.memory.M[76] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0150_)
			\mchip.dut.memory.M[76] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0150_)
			\mchip.dut.memory.M[76] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0150_)
			\mchip.dut.memory.M[76] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0119_)
			\mchip.dut.memory.M[48] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0119_)
			\mchip.dut.memory.M[48] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0119_)
			\mchip.dut.memory.M[48] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0119_)
			\mchip.dut.memory.M[48] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0119_)
			\mchip.dut.memory.M[48] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0151_)
			\mchip.dut.memory.M[77] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0151_)
			\mchip.dut.memory.M[77] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0151_)
			\mchip.dut.memory.M[77] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0151_)
			\mchip.dut.memory.M[77] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0151_)
			\mchip.dut.memory.M[77] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0152_)
			\mchip.dut.memory.M[78] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0152_)
			\mchip.dut.memory.M[78] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0152_)
			\mchip.dut.memory.M[78] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0152_)
			\mchip.dut.memory.M[78] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0152_)
			\mchip.dut.memory.M[78] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0154_)
			\mchip.dut.memory.M[7] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0154_)
			\mchip.dut.memory.M[7] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0154_)
			\mchip.dut.memory.M[7] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0154_)
			\mchip.dut.memory.M[7] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0154_)
			\mchip.dut.memory.M[7] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0155_)
			\mchip.dut.memory.M[80] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0155_)
			\mchip.dut.memory.M[80] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0155_)
			\mchip.dut.memory.M[80] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0155_)
			\mchip.dut.memory.M[80] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0155_)
			\mchip.dut.memory.M[80] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0156_)
			\mchip.dut.memory.M[81] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0156_)
			\mchip.dut.memory.M[81] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0156_)
			\mchip.dut.memory.M[81] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0156_)
			\mchip.dut.memory.M[81] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0156_)
			\mchip.dut.memory.M[81] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0157_)
			\mchip.dut.memory.M[82] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0157_)
			\mchip.dut.memory.M[82] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0157_)
			\mchip.dut.memory.M[82] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0157_)
			\mchip.dut.memory.M[82] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0157_)
			\mchip.dut.memory.M[82] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0158_)
			\mchip.dut.memory.M[83] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0158_)
			\mchip.dut.memory.M[83] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0158_)
			\mchip.dut.memory.M[83] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0158_)
			\mchip.dut.memory.M[83] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0158_)
			\mchip.dut.memory.M[83] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0159_)
			\mchip.dut.memory.M[84] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0159_)
			\mchip.dut.memory.M[84] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0159_)
			\mchip.dut.memory.M[84] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0159_)
			\mchip.dut.memory.M[84] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0159_)
			\mchip.dut.memory.M[84] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0160_)
			\mchip.dut.memory.M[85] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0160_)
			\mchip.dut.memory.M[85] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0160_)
			\mchip.dut.memory.M[85] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0160_)
			\mchip.dut.memory.M[85] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0160_)
			\mchip.dut.memory.M[85] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0161_)
			\mchip.dut.memory.M[86] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0161_)
			\mchip.dut.memory.M[86] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0161_)
			\mchip.dut.memory.M[86] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0161_)
			\mchip.dut.memory.M[86] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0161_)
			\mchip.dut.memory.M[86] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0162_)
			\mchip.dut.memory.M[87] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0162_)
			\mchip.dut.memory.M[87] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0162_)
			\mchip.dut.memory.M[87] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0162_)
			\mchip.dut.memory.M[87] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0162_)
			\mchip.dut.memory.M[87] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0163_)
			\mchip.dut.memory.M[88] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0163_)
			\mchip.dut.memory.M[88] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0163_)
			\mchip.dut.memory.M[88] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0163_)
			\mchip.dut.memory.M[88] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0163_)
			\mchip.dut.memory.M[88] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0070_)
			\mchip.dut.memory.M[119] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0070_)
			\mchip.dut.memory.M[119] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0070_)
			\mchip.dut.memory.M[119] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0070_)
			\mchip.dut.memory.M[119] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0070_)
			\mchip.dut.memory.M[119] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0130_)
			\mchip.dut.memory.M[58] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0130_)
			\mchip.dut.memory.M[58] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0130_)
			\mchip.dut.memory.M[58] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0130_)
			\mchip.dut.memory.M[58] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0130_)
			\mchip.dut.memory.M[58] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0165_)
			\mchip.dut.memory.M[8] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0165_)
			\mchip.dut.memory.M[8] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0165_)
			\mchip.dut.memory.M[8] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0165_)
			\mchip.dut.memory.M[8] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0165_)
			\mchip.dut.memory.M[8] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0122_)
			\mchip.dut.memory.M[50] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0122_)
			\mchip.dut.memory.M[50] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0122_)
			\mchip.dut.memory.M[50] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0122_)
			\mchip.dut.memory.M[50] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0122_)
			\mchip.dut.memory.M[50] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0132_)
			\mchip.dut.memory.M[5] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0132_)
			\mchip.dut.memory.M[5] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0132_)
			\mchip.dut.memory.M[5] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0132_)
			\mchip.dut.memory.M[5] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0132_)
			\mchip.dut.memory.M[5] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0123_)
			\mchip.dut.memory.M[51] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0123_)
			\mchip.dut.memory.M[51] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0123_)
			\mchip.dut.memory.M[51] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0123_)
			\mchip.dut.memory.M[51] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0123_)
			\mchip.dut.memory.M[51] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0166_)
			\mchip.dut.memory.M[90] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0166_)
			\mchip.dut.memory.M[90] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0166_)
			\mchip.dut.memory.M[90] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0166_)
			\mchip.dut.memory.M[90] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0166_)
			\mchip.dut.memory.M[90] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0133_)
			\mchip.dut.memory.M[60] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0133_)
			\mchip.dut.memory.M[60] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0133_)
			\mchip.dut.memory.M[60] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0133_)
			\mchip.dut.memory.M[60] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0133_)
			\mchip.dut.memory.M[60] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0176_)
			\mchip.dut.memory.M[9] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0176_)
			\mchip.dut.memory.M[9] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0176_)
			\mchip.dut.memory.M[9] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0176_)
			\mchip.dut.memory.M[9] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0176_)
			\mchip.dut.memory.M[9] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0124_)
			\mchip.dut.memory.M[52] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0124_)
			\mchip.dut.memory.M[52] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0124_)
			\mchip.dut.memory.M[52] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0124_)
			\mchip.dut.memory.M[52] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0124_)
			\mchip.dut.memory.M[52] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.dut.memory.M[61] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.dut.memory.M[61] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.dut.memory.M[61] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.dut.memory.M[61] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0134_)
			\mchip.dut.memory.M[61] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0167_)
			\mchip.dut.memory.M[91] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0167_)
			\mchip.dut.memory.M[91] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0167_)
			\mchip.dut.memory.M[91] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0167_)
			\mchip.dut.memory.M[91] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0167_)
			\mchip.dut.memory.M[91] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.dut.memory.M[62] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.dut.memory.M[62] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.dut.memory.M[62] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.dut.memory.M[62] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0135_)
			\mchip.dut.memory.M[62] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0125_)
			\mchip.dut.memory.M[53] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0125_)
			\mchip.dut.memory.M[53] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0125_)
			\mchip.dut.memory.M[53] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0125_)
			\mchip.dut.memory.M[53] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0125_)
			\mchip.dut.memory.M[53] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0168_)
			\mchip.dut.memory.M[92] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0168_)
			\mchip.dut.memory.M[92] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0168_)
			\mchip.dut.memory.M[92] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0168_)
			\mchip.dut.memory.M[92] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0168_)
			\mchip.dut.memory.M[92] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0136_)
			\mchip.dut.memory.M[63] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0136_)
			\mchip.dut.memory.M[63] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0136_)
			\mchip.dut.memory.M[63] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0136_)
			\mchip.dut.memory.M[63] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0136_)
			\mchip.dut.memory.M[63] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0169_)
			\mchip.dut.memory.M[93] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0169_)
			\mchip.dut.memory.M[93] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0169_)
			\mchip.dut.memory.M[93] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0169_)
			\mchip.dut.memory.M[93] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0169_)
			\mchip.dut.memory.M[93] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0137_)
			\mchip.dut.memory.M[64] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0137_)
			\mchip.dut.memory.M[64] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0137_)
			\mchip.dut.memory.M[64] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0137_)
			\mchip.dut.memory.M[64] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0137_)
			\mchip.dut.memory.M[64] [4] <= \mchip.dut.memory.data_in [4];
	reg \mchip.dut.next_state.Q_reg[0] ;
	always @(posedge io_in[12])
		if (\mchip.dut.NextState_en )
			if (\mchip.dut.fsm.currState [0])
				\mchip.dut.next_state.Q_reg[0]  <= 1'h1;
			else
				\mchip.dut.next_state.Q_reg[0]  <= \mchip.dut.demux.Y2 [0];
	assign \mchip.dut.next_state.Q [0] = \mchip.dut.next_state.Q_reg[0] ;
	always @(posedge io_in[12])
		if (_0170_)
			\mchip.dut.memory.M[94] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0170_)
			\mchip.dut.memory.M[94] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0170_)
			\mchip.dut.memory.M[94] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0170_)
			\mchip.dut.memory.M[94] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0170_)
			\mchip.dut.memory.M[94] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0138_)
			\mchip.dut.memory.M[65] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0138_)
			\mchip.dut.memory.M[65] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0138_)
			\mchip.dut.memory.M[65] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0138_)
			\mchip.dut.memory.M[65] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0138_)
			\mchip.dut.memory.M[65] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0171_)
			\mchip.dut.memory.M[95] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0171_)
			\mchip.dut.memory.M[95] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0171_)
			\mchip.dut.memory.M[95] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0171_)
			\mchip.dut.memory.M[95] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0171_)
			\mchip.dut.memory.M[95] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0139_)
			\mchip.dut.memory.M[66] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0139_)
			\mchip.dut.memory.M[66] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0139_)
			\mchip.dut.memory.M[66] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0139_)
			\mchip.dut.memory.M[66] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0139_)
			\mchip.dut.memory.M[66] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0172_)
			\mchip.dut.memory.M[96] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0172_)
			\mchip.dut.memory.M[96] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0172_)
			\mchip.dut.memory.M[96] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0172_)
			\mchip.dut.memory.M[96] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0172_)
			\mchip.dut.memory.M[96] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0140_)
			\mchip.dut.memory.M[67] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0140_)
			\mchip.dut.memory.M[67] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0140_)
			\mchip.dut.memory.M[67] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0140_)
			\mchip.dut.memory.M[67] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0140_)
			\mchip.dut.memory.M[67] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0121_)
			\mchip.dut.memory.M[4] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0121_)
			\mchip.dut.memory.M[4] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0121_)
			\mchip.dut.memory.M[4] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0121_)
			\mchip.dut.memory.M[4] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0121_)
			\mchip.dut.memory.M[4] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0141_)
			\mchip.dut.memory.M[68] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0141_)
			\mchip.dut.memory.M[68] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0141_)
			\mchip.dut.memory.M[68] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0141_)
			\mchip.dut.memory.M[68] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0141_)
			\mchip.dut.memory.M[68] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0173_)
			\mchip.dut.memory.M[97] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0173_)
			\mchip.dut.memory.M[97] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0173_)
			\mchip.dut.memory.M[97] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0173_)
			\mchip.dut.memory.M[97] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0173_)
			\mchip.dut.memory.M[97] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0143_)
			\mchip.dut.memory.M[6] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0143_)
			\mchip.dut.memory.M[6] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0143_)
			\mchip.dut.memory.M[6] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0143_)
			\mchip.dut.memory.M[6] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0143_)
			\mchip.dut.memory.M[6] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0086_)
			\mchip.dut.memory.M[18] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0086_)
			\mchip.dut.memory.M[18] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0086_)
			\mchip.dut.memory.M[18] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0086_)
			\mchip.dut.memory.M[18] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0086_)
			\mchip.dut.memory.M[18] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0144_)
			\mchip.dut.memory.M[70] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0144_)
			\mchip.dut.memory.M[70] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0144_)
			\mchip.dut.memory.M[70] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0144_)
			\mchip.dut.memory.M[70] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0144_)
			\mchip.dut.memory.M[70] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0145_)
			\mchip.dut.memory.M[71] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0145_)
			\mchip.dut.memory.M[71] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0145_)
			\mchip.dut.memory.M[71] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0145_)
			\mchip.dut.memory.M[71] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0145_)
			\mchip.dut.memory.M[71] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0174_)
			\mchip.dut.memory.M[98] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0174_)
			\mchip.dut.memory.M[98] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0174_)
			\mchip.dut.memory.M[98] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0174_)
			\mchip.dut.memory.M[98] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0174_)
			\mchip.dut.memory.M[98] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0019_)
			if (_0021_)
				\mchip.dut.data_reg.Q  <= 1'h0;
			else
				\mchip.dut.data_reg.Q  <= \mchip.dut.demux.I [0];
	always @(posedge io_in[12])
		if (_0087_)
			\mchip.dut.memory.M[19] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0087_)
			\mchip.dut.memory.M[19] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0087_)
			\mchip.dut.memory.M[19] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0087_)
			\mchip.dut.memory.M[19] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0087_)
			\mchip.dut.memory.M[19] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0049_)
			\mchip.dut.memory.M[0] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0049_)
			\mchip.dut.memory.M[0] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0049_)
			\mchip.dut.memory.M[0] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0049_)
			\mchip.dut.memory.M[0] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0049_)
			\mchip.dut.memory.M[0] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0050_)
			\mchip.dut.memory.M[100] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0050_)
			\mchip.dut.memory.M[100] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0050_)
			\mchip.dut.memory.M[100] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0050_)
			\mchip.dut.memory.M[100] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0050_)
			\mchip.dut.memory.M[100] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0126_)
			\mchip.dut.memory.M[54] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0126_)
			\mchip.dut.memory.M[54] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0126_)
			\mchip.dut.memory.M[54] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0126_)
			\mchip.dut.memory.M[54] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0126_)
			\mchip.dut.memory.M[54] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0051_)
			\mchip.dut.memory.M[101] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0051_)
			\mchip.dut.memory.M[101] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0051_)
			\mchip.dut.memory.M[101] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0051_)
			\mchip.dut.memory.M[101] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0051_)
			\mchip.dut.memory.M[101] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0127_)
			\mchip.dut.memory.M[55] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0127_)
			\mchip.dut.memory.M[55] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0127_)
			\mchip.dut.memory.M[55] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0127_)
			\mchip.dut.memory.M[55] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0127_)
			\mchip.dut.memory.M[55] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0128_)
			\mchip.dut.memory.M[56] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0128_)
			\mchip.dut.memory.M[56] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0128_)
			\mchip.dut.memory.M[56] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0128_)
			\mchip.dut.memory.M[56] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0128_)
			\mchip.dut.memory.M[56] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0052_)
			\mchip.dut.memory.M[102] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0052_)
			\mchip.dut.memory.M[102] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0052_)
			\mchip.dut.memory.M[102] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0052_)
			\mchip.dut.memory.M[102] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0052_)
			\mchip.dut.memory.M[102] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0129_)
			\mchip.dut.memory.M[57] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0129_)
			\mchip.dut.memory.M[57] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0129_)
			\mchip.dut.memory.M[57] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0129_)
			\mchip.dut.memory.M[57] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0129_)
			\mchip.dut.memory.M[57] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0014_)
			if (!\mchip.dut.StateAddr_ld )
				\mchip.dut.tape_reg.Q  <= 1'h0;
			else
				\mchip.dut.tape_reg.Q  <= \mchip.dut.tape_reg.D ;
	always @(posedge io_in[12])
		if (_0016_)
			\mchip.dut.state_addr.Q [0] <= _0035_;
	always @(posedge io_in[12])
		if (_0016_)
			\mchip.dut.state_addr.Q [1] <= _0036_;
	always @(posedge io_in[12])
		if (_0016_)
			\mchip.dut.state_addr.Q [2] <= _0037_;
	always @(posedge io_in[12])
		if (_0016_)
			\mchip.dut.state_addr.Q [3] <= _0038_;
	always @(posedge io_in[12])
		if (_0016_)
			\mchip.dut.state_addr.Q [4] <= _0039_;
	always @(posedge io_in[12])
		if (_0016_)
			\mchip.dut.state_addr.Q [5] <= _0040_;
	always @(posedge io_in[12])
		if (_0016_)
			\mchip.dut.state_addr.Q [6] <= _0041_;
	always @(posedge io_in[12])
		if (_0059_)
			\mchip.dut.memory.M[109] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0059_)
			\mchip.dut.memory.M[109] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0059_)
			\mchip.dut.memory.M[109] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0059_)
			\mchip.dut.memory.M[109] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0059_)
			\mchip.dut.memory.M[109] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.dut.tape_addr.Q [0] <= _0042_;
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.dut.tape_addr.Q [1] <= _0043_;
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.dut.tape_addr.Q [2] <= _0044_;
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.dut.tape_addr.Q [3] <= _0045_;
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.dut.tape_addr.Q [4] <= _0046_;
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.dut.tape_addr.Q [5] <= _0047_;
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.dut.tape_addr.Q [6] <= _0048_;
	always @(posedge io_in[12])
		if (_0053_)
			\mchip.dut.memory.M[103] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0053_)
			\mchip.dut.memory.M[103] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0053_)
			\mchip.dut.memory.M[103] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0053_)
			\mchip.dut.memory.M[103] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0053_)
			\mchip.dut.memory.M[103] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0054_)
			\mchip.dut.memory.M[104] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0054_)
			\mchip.dut.memory.M[104] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0054_)
			\mchip.dut.memory.M[104] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0054_)
			\mchip.dut.memory.M[104] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0054_)
			\mchip.dut.memory.M[104] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0055_)
			\mchip.dut.memory.M[105] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0055_)
			\mchip.dut.memory.M[105] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0055_)
			\mchip.dut.memory.M[105] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0055_)
			\mchip.dut.memory.M[105] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0055_)
			\mchip.dut.memory.M[105] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0056_)
			\mchip.dut.memory.M[106] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0056_)
			\mchip.dut.memory.M[106] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0056_)
			\mchip.dut.memory.M[106] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0056_)
			\mchip.dut.memory.M[106] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0056_)
			\mchip.dut.memory.M[106] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12])
		if (_0175_)
			\mchip.dut.memory.M[99] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0175_)
			\mchip.dut.memory.M[99] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0175_)
			\mchip.dut.memory.M[99] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0175_)
			\mchip.dut.memory.M[99] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0175_)
			\mchip.dut.memory.M[99] [4] <= \mchip.dut.memory.data_in [4];
	reg \mchip.dut.direction_reg.Q_reg[0] ;
	always @(posedge io_in[12])
		if (_0018_)
			if (_0022_)
				\mchip.dut.direction_reg.Q_reg[0]  <= 1'h0;
			else
				\mchip.dut.direction_reg.Q_reg[0]  <= \mchip.dut.demux.I [0];
	assign \mchip.dut.direction_reg.Q [0] = \mchip.dut.direction_reg.Q_reg[0] ;
	reg \mchip.dut.direction_reg.Q_reg[1] ;
	always @(posedge io_in[12])
		if (_0018_)
			if (_0022_)
				\mchip.dut.direction_reg.Q_reg[1]  <= 1'h0;
			else
				\mchip.dut.direction_reg.Q_reg[1]  <= \mchip.dut.demux.I [1];
	assign \mchip.dut.direction_reg.Q [1] = \mchip.dut.direction_reg.Q_reg[1] ;
	always @(posedge io_in[12])
		if (\mchip.dut.fsm.currState [0])
			\mchip.dut.display_reg.Q [0] <= 1'h0;
		else if (_0017_)
			\mchip.dut.display_reg.Q [0] <= _0024_;
	always @(posedge io_in[12])
		if (_0164_)
			\mchip.dut.memory.M[89] [0] <= \mchip.dut.memory.data_in [0];
	always @(posedge io_in[12])
		if (_0164_)
			\mchip.dut.memory.M[89] [1] <= \mchip.dut.memory.data_in [1];
	always @(posedge io_in[12])
		if (_0164_)
			\mchip.dut.memory.M[89] [2] <= \mchip.dut.memory.data_in [2];
	always @(posedge io_in[12])
		if (_0164_)
			\mchip.dut.memory.M[89] [3] <= \mchip.dut.memory.data_in [3];
	always @(posedge io_in[12])
		if (_0164_)
			\mchip.dut.memory.M[89] [4] <= \mchip.dut.memory.data_in [4];
	always @(posedge io_in[12]) \mchip.sync8.async1  <= io_in[7];
	always @(posedge io_in[12]) \mchip.sync7.async1  <= io_in[6];
	always @(posedge io_in[12]) \mchip.sync6.async1  <= io_in[5];
	always @(posedge io_in[12]) \mchip.sync5.async1  <= io_in[4];
	always @(posedge io_in[12]) \mchip.sync4.async1  <= io_in[3];
	always @(posedge io_in[12]) \mchip.sync3.async1  <= io_in[2];
	always @(posedge io_in[12]) \mchip.sync2.async1  <= io_in[0];
	always @(posedge io_in[12]) \mchip.sync1.async1  <= io_in[1];
	always @(posedge io_in[12]) \mchip.sync8.sync  <= \mchip.sync8.async1 ;
	always @(posedge io_in[12]) \mchip.sync7.sync  <= \mchip.sync7.async1 ;
	always @(posedge io_in[12]) \mchip.sync6.sync  <= \mchip.sync6.async1 ;
	always @(posedge io_in[12]) \mchip.sync5.sync  <= \mchip.sync5.async1 ;
	always @(posedge io_in[12]) \mchip.sync4.sync  <= \mchip.sync4.async1 ;
	always @(posedge io_in[12]) \mchip.sync3.sync  <= \mchip.sync3.async1 ;
	always @(posedge io_in[12]) \mchip.sync2.sync  <= \mchip.sync2.async1 ;
	always @(posedge io_in[12]) \mchip.sync1.sync  <= \mchip.sync1.async1 ;
	assign io_out = {2'h0, \mchip.dut.display_reg.Q , \mchip.dut.Compute_done };
	assign \mchip.Done  = \mchip.sync2.sync ;
	assign \mchip.Next  = \mchip.sync1.sync ;
	assign \mchip.clock  = io_in[12];
	assign \mchip.dut.DataReg_en  = \mchip.dut.fsm.currState [9];
	assign \mchip.dut.Done  = \mchip.sync2.sync ;
	assign \mchip.dut.Halt  = \mchip.dut.direction_reg.Q [1];
	assign \mchip.dut.Init  = \mchip.dut.fsm.currState [0];
	assign \mchip.dut.Left  = \mchip.dut.direction_reg.Q [0];
	assign \mchip.dut.Next  = \mchip.sync1.sync ;
	assign \mchip.dut.Read_en  = 1'h1;
	assign \mchip.dut.TapeReg_en  = \mchip.dut.StateAddr_ld ;
	assign \mchip.dut.Tape_start  = 1'h1;
	assign \mchip.dut.clock  = io_in[12];
	assign \mchip.dut.data_reg.clear  = \mchip.dut.fsm.currState [0];
	assign \mchip.dut.data_reg.clock  = io_in[12];
	assign \mchip.dut.data_reg.en  = \mchip.dut.fsm.currState [9];
	assign \mchip.dut.data_reg_out  = \mchip.dut.data_reg.Q ;
	assign \mchip.dut.demux.Y0  = 5'h00;
	assign \mchip.dut.demux.Y1  = 5'h00;
	assign \mchip.dut.demux.Y2 [4:1] = 4'h0;
	assign \mchip.dut.demux.Y3  = 5'h00;
	assign \mchip.dut.direction_in  = 2'h0;
	assign \mchip.dut.direction_out  = \mchip.dut.direction_reg.Q [1:0];
	assign \mchip.dut.direction_reg.D  = 7'h00;
	assign \mchip.dut.direction_reg.Q [6:2] = 5'h00;
	assign \mchip.dut.direction_reg.clear  = \mchip.dut.fsm.currState [0];
	assign \mchip.dut.direction_reg.clock  = io_in[12];
	assign \mchip.dut.display_out  = \mchip.dut.display_reg.Q ;
	assign \mchip.dut.display_reg.clear  = \mchip.dut.fsm.currState [0];
	assign \mchip.dut.display_reg.clock  = io_in[12];
	assign \mchip.dut.fsm.DataReg_en  = \mchip.dut.fsm.currState [9];
	assign \mchip.dut.fsm.Done  = \mchip.sync2.sync ;
	assign \mchip.dut.fsm.Halt  = \mchip.dut.direction_reg.Q [1];
	assign \mchip.dut.fsm.Init  = \mchip.dut.fsm.currState [0];
	assign \mchip.dut.fsm.InputAddr_en  = \mchip.dut.InputAddr_en ;
	assign \mchip.dut.fsm.Left  = \mchip.dut.direction_reg.Q [0];
	assign \mchip.dut.fsm.Next  = \mchip.sync1.sync ;
	assign \mchip.dut.fsm.NextState_en  = \mchip.dut.NextState_en ;
	assign \mchip.dut.fsm.Read_en  = 1'h1;
	assign \mchip.dut.fsm.StateAddr_ld  = \mchip.dut.StateAddr_ld ;
	assign \mchip.dut.fsm.TapeReg_en  = \mchip.dut.StateAddr_ld ;
	assign \mchip.dut.fsm.Tape_start  = 1'h1;
	assign \mchip.dut.fsm.clock  = io_in[12];
	assign \mchip.dut.fsm.currState [7] = 1'h0;
	assign \mchip.dut.fsm.reset  = io_in[13];
	assign \mchip.dut.input_addr.clear  = \mchip.dut.fsm.currState [0];
	assign \mchip.dut.input_addr.clock  = io_in[12];
	assign \mchip.dut.input_addr.en  = \mchip.dut.InputAddr_en ;
	assign \mchip.dut.input_addr.load  = 1'h0;
	assign \mchip.dut.input_addr.up  = 1'h1;
	assign \mchip.dut.input_addr_out  = \mchip.dut.input_addr.Q ;
	assign \mchip.dut.input_data  = {1'h0, \mchip.sync8.sync , \mchip.sync7.sync , \mchip.sync6.sync , \mchip.sync5.sync , \mchip.sync4.sync , \mchip.sync3.sync };
	assign \mchip.dut.memory.clock  = io_in[12];
	assign \mchip.dut.memory.data_out  = \mchip.dut.demux.I ;
	assign \mchip.dut.memory.re  = 1'h1;
	assign \mchip.dut.mux_display.I0  = {6'h00, \mchip.dut.tape_reg.Q };
	assign \mchip.dut.mux_display.I1  = 7'h00;
	assign \mchip.dut.mux_display.S  = \mchip.dut.direction_reg.Q [0];
	assign \mchip.dut.mux_display.Y  = 7'h00;
	assign \mchip.dut.mux_input_calculate.I0  = {4'h0, \mchip.dut.data_reg.Q };
	assign \mchip.dut.mux_input_calculate.I1  = {\mchip.sync7.sync , \mchip.sync6.sync , \mchip.sync5.sync , \mchip.sync4.sync , \mchip.sync3.sync };
	assign \mchip.dut.mux_input_calculate.Y  = \mchip.dut.memory.data_in ;
	assign \mchip.dut.mux_next_state.I0  = {6'h00, \mchip.dut.demux.Y2 [0]};
	assign \mchip.dut.mux_next_state.I1  = 7'h01;
	assign \mchip.dut.mux_next_state.S  = \mchip.dut.fsm.currState [0];
	assign \mchip.dut.mux_next_state.Y  = 7'h00;
	assign \mchip.dut.mux_prev_tape.I0  = 1'h0;
	assign \mchip.dut.mux_prev_tape.I1  = 1'h0;
	assign \mchip.dut.mux_prev_tape.Y  = 1'h0;
	assign \mchip.dut.mux_state_tape_addr.I0  = \mchip.dut.state_addr.Q ;
	assign \mchip.dut.mux_state_tape_addr.I1  = \mchip.dut.tape_addr.Q ;
	assign \mchip.dut.mux_state_tape_addr.I3  = \mchip.dut.input_addr.Q ;
	assign \mchip.dut.mux_tape_reg.I0  = 1'h0;
	assign \mchip.dut.mux_tape_reg.I1  = \mchip.dut.display_reg.Q [1];
	assign \mchip.dut.mux_tape_reg.S  = \mchip.dut.direction_reg.Q [0];
	assign \mchip.dut.mux_tape_reg.Y  = \mchip.dut.tape_reg.D ;
	assign \mchip.dut.next_state.D  = 7'h00;
	assign \mchip.dut.next_state.Q [6:5] = 2'h0;
	assign \mchip.dut.next_state.clear  = 1'h0;
	assign \mchip.dut.next_state.clock  = io_in[12];
	assign \mchip.dut.next_state.en  = \mchip.dut.NextState_en ;
	assign \mchip.dut.next_state_in  = 7'h00;
	assign \mchip.dut.next_state_out  = {2'h0, \mchip.dut.next_state.Q [4:0]};
	assign \mchip.dut.next_state_prep  = {6'h00, \mchip.dut.demux.Y2 [0]};
	assign \mchip.dut.prev_tape_in  = 1'h0;
	assign \mchip.dut.prev_tape_out  = 1'h0;
	assign \mchip.dut.prev_tape_reg.D  = 1'h0;
	assign \mchip.dut.prev_tape_reg.Q  = 1'h0;
	assign \mchip.dut.prev_tape_reg.clear  = \mchip.dut.fsm.currState [0];
	assign \mchip.dut.prev_tape_reg.clock  = io_in[12];
	assign \mchip.dut.read_data  = \mchip.dut.demux.I ;
	assign \mchip.dut.reset  = io_in[13];
	assign \mchip.dut.state_addr.D  = 7'h00;
	assign \mchip.dut.state_addr.clear  = 1'h0;
	assign \mchip.dut.state_addr.clock  = io_in[12];
	assign \mchip.dut.state_addr.load  = \mchip.dut.StateAddr_ld ;
	assign \mchip.dut.state_addr.up  = 1'h1;
	assign \mchip.dut.state_addr_in  = 7'h00;
	assign \mchip.dut.state_addr_out  = \mchip.dut.state_addr.Q ;
	assign \mchip.dut.tape_addr.D  = {1'h0, \mchip.sync8.sync , \mchip.sync7.sync , \mchip.sync6.sync , \mchip.sync5.sync , \mchip.sync4.sync , \mchip.sync3.sync };
	assign \mchip.dut.tape_addr.clear  = 1'h0;
	assign \mchip.dut.tape_addr.clock  = io_in[12];
	assign \mchip.dut.tape_addr_init.D  = {1'h0, \mchip.sync8.sync , \mchip.sync7.sync , \mchip.sync6.sync , \mchip.sync5.sync , \mchip.sync4.sync , \mchip.sync3.sync };
	assign \mchip.dut.tape_addr_init.Q  = 7'h00;
	assign \mchip.dut.tape_addr_init.clear  = 1'h0;
	assign \mchip.dut.tape_addr_init.clock  = io_in[12];
	assign \mchip.dut.tape_addr_min.D [1:0] = {\mchip.sync3.sync , 1'h1};
	assign \mchip.dut.tape_addr_min.Q [0] = 1'h1;
	assign \mchip.dut.tape_addr_min.clear  = 1'h0;
	assign \mchip.dut.tape_addr_min.clock  = io_in[12];
	assign \mchip.dut.tape_addr_min.en  = \mchip.dut.fsm.currState [0];
	assign \mchip.dut.tape_addr_out  = \mchip.dut.tape_addr.Q ;
	assign \mchip.dut.tape_in  = 1'h0;
	assign \mchip.dut.tape_init_addr  = 7'h00;
	assign \mchip.dut.tape_min_addr_in  = {\mchip.dut.tape_addr_min.D [6:2], \mchip.sync3.sync , 1'h1};
	assign \mchip.dut.tape_min_addr_out  = {\mchip.dut.tape_addr_min.Q [6:1], 1'h1};
	assign \mchip.dut.tape_reg.clear  = \mchip.dut.fsm.currState [0];
	assign \mchip.dut.tape_reg.clock  = io_in[12];
	assign \mchip.dut.tape_reg.en  = \mchip.dut.StateAddr_ld ;
	assign \mchip.dut.tape_reg_in  = \mchip.dut.tape_reg.D ;
	assign \mchip.dut.tape_reg_out  = \mchip.dut.tape_reg.Q ;
	assign \mchip.dut.write_data  = \mchip.dut.memory.data_in ;
	assign \mchip.input_data  = {1'h0, \mchip.sync8.sync , \mchip.sync7.sync , \mchip.sync6.sync , \mchip.sync5.sync , \mchip.sync4.sync , \mchip.sync3.sync };
	assign \mchip.io_in  = io_in[11:0];
	assign \mchip.io_out  = {\mchip.dut.display_reg.Q , \mchip.dut.Compute_done };
	assign \mchip.reset  = io_in[13];
	assign \mchip.sync1.async  = io_in[1];
	assign \mchip.sync1.clock  = io_in[12];
	assign \mchip.sync2.async  = io_in[0];
	assign \mchip.sync2.clock  = io_in[12];
	assign \mchip.sync3.async  = io_in[2];
	assign \mchip.sync3.clock  = io_in[12];
	assign \mchip.sync4.async  = io_in[3];
	assign \mchip.sync4.clock  = io_in[12];
	assign \mchip.sync5.async  = io_in[4];
	assign \mchip.sync5.clock  = io_in[12];
	assign \mchip.sync6.async  = io_in[5];
	assign \mchip.sync6.clock  = io_in[12];
	assign \mchip.sync7.async  = io_in[6];
	assign \mchip.sync7.clock  = io_in[12];
	assign \mchip.sync8.async  = io_in[7];
	assign \mchip.sync8.clock  = io_in[12];
endmodule
module d24_mnguyen2_tpu (
	io_in,
	io_out
);
	wire _000_;
	wire _001_;
	wire _002_;
	wire _003_;
	wire _004_;
	wire _005_;
	wire _006_;
	wire _007_;
	wire _008_;
	wire _009_;
	wire _010_;
	wire _011_;
	wire _012_;
	wire _013_;
	wire _014_;
	wire _015_;
	wire _016_;
	wire _017_;
	wire _018_;
	wire _019_;
	wire _020_;
	wire _021_;
	wire _022_;
	wire _023_;
	wire _024_;
	wire _025_;
	wire _026_;
	wire _027_;
	wire _028_;
	wire _029_;
	wire _030_;
	wire _031_;
	wire _032_;
	wire _033_;
	wire _034_;
	wire _035_;
	wire _036_;
	wire _037_;
	wire _038_;
	wire _039_;
	wire _040_;
	wire _041_;
	wire _042_;
	wire _043_;
	wire _044_;
	wire _045_;
	wire _046_;
	wire _047_;
	wire _048_;
	wire _049_;
	wire _050_;
	wire _051_;
	wire _052_;
	wire _053_;
	wire _054_;
	wire _055_;
	wire _056_;
	wire _057_;
	wire _058_;
	wire _059_;
	wire _060_;
	wire _061_;
	wire _062_;
	wire _063_;
	wire _064_;
	wire _065_;
	wire _066_;
	wire _067_;
	wire _068_;
	wire _069_;
	wire _070_;
	wire _071_;
	wire _072_;
	wire _073_;
	wire _074_;
	wire _075_;
	wire _076_;
	wire _077_;
	wire _078_;
	wire _079_;
	wire _080_;
	wire _081_;
	wire _082_;
	wire _083_;
	wire _084_;
	wire _085_;
	wire _086_;
	wire _087_;
	wire _088_;
	wire _089_;
	wire _090_;
	wire _091_;
	wire _092_;
	wire _093_;
	wire _094_;
	wire _095_;
	wire _096_;
	wire _097_;
	wire _098_;
	wire _099_;
	wire _100_;
	wire _101_;
	wire _102_;
	wire _103_;
	wire _104_;
	wire _105_;
	wire _106_;
	wire _107_;
	wire _108_;
	wire _109_;
	wire _110_;
	wire _111_;
	wire _112_;
	wire _113_;
	wire _114_;
	wire _115_;
	wire _116_;
	wire _117_;
	wire _118_;
	wire _119_;
	wire _120_;
	wire _121_;
	wire _122_;
	wire _123_;
	wire _124_;
	wire _125_;
	wire _126_;
	wire _127_;
	wire _128_;
	wire _129_;
	wire _130_;
	wire _131_;
	wire _132_;
	wire _133_;
	wire _134_;
	wire _135_;
	wire _136_;
	wire _137_;
	wire _138_;
	wire _139_;
	wire _140_;
	wire _141_;
	wire _142_;
	wire _143_;
	wire _144_;
	wire _145_;
	wire _146_;
	wire _147_;
	wire _148_;
	wire _149_;
	wire _150_;
	wire _151_;
	wire _152_;
	wire _153_;
	wire _154_;
	wire _155_;
	wire _156_;
	wire _157_;
	wire _158_;
	wire _159_;
	wire _160_;
	wire _161_;
	wire _162_;
	wire _163_;
	wire _164_;
	wire _165_;
	wire _166_;
	wire _167_;
	wire _168_;
	wire _169_;
	wire _170_;
	wire _171_;
	wire _172_;
	wire _173_;
	wire _174_;
	wire _175_;
	wire _176_;
	wire _177_;
	wire _178_;
	wire _179_;
	wire _180_;
	wire _181_;
	wire _182_;
	wire _183_;
	wire _184_;
	wire _185_;
	wire _186_;
	wire _187_;
	wire _188_;
	wire _189_;
	wire _190_;
	wire _191_;
	wire _192_;
	wire _193_;
	wire _194_;
	wire _195_;
	wire _196_;
	wire _197_;
	wire _198_;
	wire _199_;
	wire _200_;
	wire _201_;
	wire _202_;
	wire _203_;
	wire _204_;
	wire _205_;
	wire _206_;
	wire _207_;
	wire _208_;
	wire _209_;
	wire _210_;
	wire _211_;
	wire _212_;
	wire _213_;
	wire _214_;
	wire _215_;
	wire _216_;
	wire _217_;
	wire _218_;
	wire _219_;
	wire _220_;
	wire _221_;
	wire _222_;
	wire _223_;
	wire _224_;
	wire _225_;
	wire _226_;
	wire _227_;
	wire _228_;
	wire _229_;
	wire _230_;
	wire _231_;
	wire _232_;
	wire _233_;
	wire _234_;
	wire _235_;
	wire _236_;
	wire _237_;
	wire _238_;
	wire _239_;
	wire _240_;
	wire _241_;
	wire _242_;
	wire _243_;
	wire _244_;
	wire _245_;
	wire _246_;
	wire _247_;
	wire _248_;
	wire _249_;
	wire _250_;
	wire _251_;
	wire _252_;
	wire _253_;
	wire _254_;
	wire _255_;
	wire _256_;
	wire _257_;
	wire _258_;
	wire _259_;
	wire _260_;
	wire _261_;
	wire _262_;
	wire _263_;
	wire _264_;
	wire _265_;
	wire _266_;
	wire _267_;
	wire _268_;
	wire _269_;
	wire _270_;
	wire _271_;
	wire _272_;
	wire _273_;
	wire _274_;
	wire _275_;
	wire _276_;
	wire _277_;
	wire _278_;
	wire _279_;
	wire _280_;
	wire _281_;
	wire _282_;
	wire _283_;
	wire _284_;
	wire _285_;
	wire _286_;
	wire _287_;
	wire _288_;
	wire _289_;
	wire _290_;
	wire _291_;
	wire _292_;
	wire _293_;
	wire _294_;
	wire _295_;
	wire _296_;
	wire _297_;
	wire _298_;
	wire _299_;
	wire _300_;
	wire _301_;
	wire _302_;
	wire _303_;
	wire _304_;
	wire _305_;
	wire _306_;
	wire _307_;
	wire _308_;
	wire _309_;
	wire _310_;
	wire _311_;
	wire _312_;
	wire _313_;
	wire _314_;
	wire _315_;
	wire _316_;
	wire _317_;
	wire _318_;
	wire _319_;
	wire _320_;
	wire _321_;
	wire _322_;
	wire _323_;
	wire _324_;
	wire _325_;
	wire _326_;
	wire _327_;
	wire _328_;
	wire _329_;
	wire _330_;
	wire _331_;
	wire _332_;
	wire _333_;
	wire _334_;
	wire _335_;
	wire _336_;
	wire _337_;
	wire _338_;
	wire _339_;
	wire _340_;
	wire _341_;
	wire _342_;
	wire _343_;
	wire _344_;
	wire _345_;
	wire _346_;
	wire _347_;
	wire _348_;
	wire _349_;
	wire _350_;
	wire _351_;
	wire _352_;
	input wire [13:0] io_in;
	output wire [13:0] io_out;
	wire [7:0] \mchip.TPU.KERNAL_MAT.D ;
	wire [7:0] \mchip.TPU.KERNAL_MAT.Q ;
	wire \mchip.TPU.KERNAL_MAT.clk ;
	reg [7:0] \mchip.TPU.KERNAL_MAT.data ;
	wire \mchip.TPU.KERNAL_MAT.rst ;
	wire \mchip.TPU.KERNAL_MAT.we ;
	wire [7:0] \mchip.TPU.MATRIX_MAT.D ;
	wire [7:0] \mchip.TPU.MATRIX_MAT.Q ;
	wire \mchip.TPU.MATRIX_MAT.clk ;
	reg [7:0] \mchip.TPU.MATRIX_MAT.data ;
	wire \mchip.TPU.MATRIX_MAT.rst ;
	wire \mchip.TPU.MATRIX_MAT.we ;
	wire [9:0] \mchip.TPU.base_addr ;
	reg [9:0] \mchip.TPU.base_addr_x_counter.Q ;
	wire [9:0] \mchip.TPU.base_addr_x_counter.Q_next ;
	wire \mchip.TPU.base_addr_x_counter.clk ;
	wire \mchip.TPU.base_addr_x_counter.rst ;
	reg [9:0] \mchip.TPU.base_addr_y_counter.Q ;
	wire [9:0] \mchip.TPU.base_addr_y_counter.Q_next ;
	wire \mchip.TPU.base_addr_y_counter.clk ;
	wire \mchip.TPU.base_addr_y_counter.rst ;
	wire \mchip.TPU.clk ;
	wire [7:0] \mchip.TPU.conv_mac.a ;
	wire [7:0] \mchip.TPU.conv_mac.b ;
	wire \mchip.TPU.conv_mac.clk ;
	wire \mchip.TPU.conv_mac.en ;
	wire [7:0] \mchip.TPU.conv_mac.new_sum ;
	wire [7:0] \mchip.TPU.conv_mac.prod ;
	wire \mchip.TPU.conv_mac.rst ;
	wire [7:0] \mchip.TPU.conv_mac.sum ;
	wire [7:0] \mchip.TPU.conv_mac.sum_reg.D ;
	reg [7:0] \mchip.TPU.conv_mac.sum_reg.Q ;
	wire \mchip.TPU.conv_mac.sum_reg.clk ;
	wire \mchip.TPU.conv_mac.sum_reg.rst ;
	wire \mchip.TPU.conv_mac.sum_reg.we ;
	wire [7:0] \mchip.TPU.data_in ;
	wire [7:0] \mchip.TPU.data_out ;
	wire \mchip.TPU.done ;
	wire \mchip.TPU.insert_kernal ;
	wire [3:0] \mchip.TPU.kernal_addr ;
	reg [3:0] \mchip.TPU.kernal_addr_x_counter.Q ;
	wire [3:0] \mchip.TPU.kernal_addr_x_counter.Q_next ;
	wire \mchip.TPU.kernal_addr_x_counter.clk ;
	wire \mchip.TPU.kernal_addr_x_counter.en ;
	wire \mchip.TPU.kernal_addr_x_counter.rst ;
	reg [3:0] \mchip.TPU.kernal_addr_y_counter.Q ;
	wire [3:0] \mchip.TPU.kernal_addr_y_counter.Q_next ;
	wire \mchip.TPU.kernal_addr_y_counter.clk ;
	wire \mchip.TPU.kernal_addr_y_counter.rst ;
	wire [7:0] \mchip.TPU.kernal_data ;
	wire \mchip.TPU.kernal_x_incr ;
	wire \mchip.TPU.mac_en ;
	wire \mchip.TPU.mac_rst ;
	wire [7:0] \mchip.TPU.matrix_data ;
	wire \mchip.TPU.ready ;
	wire \mchip.TPU.rst ;
	wire \mchip.TPU.write ;
	wire \mchip.TPU.write_mode ;
	wire \mchip.clock ;
	wire [11:0] \mchip.io_in ;
	wire [11:0] \mchip.io_out ;
	wire \mchip.reset ;
	assign _000_ = \mchip.TPU.kernal_addr_x_counter.Q [0] | ~\mchip.TPU.kernal_addr_x_counter.Q [1];
	assign _019_ = ~\mchip.TPU.base_addr_x_counter.Q [4];
	assign _020_ = \mchip.TPU.base_addr_x_counter.Q [0] & \mchip.TPU.base_addr_x_counter.Q [1];
	assign _021_ = \mchip.TPU.base_addr_x_counter.Q [2] & \mchip.TPU.base_addr_x_counter.Q [3];
	assign _022_ = _021_ & _020_;
	assign _017_ = _022_ & ~_019_;
	assign _023_ = \mchip.TPU.kernal_addr_x_counter.Q [2] | \mchip.TPU.kernal_addr_x_counter.Q [3];
	assign _024_ = ~(_023_ | _000_);
	assign \mchip.TPU.kernal_addr_x_counter.Q_next [0] = ~(_024_ | \mchip.TPU.kernal_addr_x_counter.Q [0]);
	assign _025_ = \mchip.TPU.kernal_addr_x_counter.Q [0] & ~\mchip.TPU.kernal_addr_x_counter.Q [1];
	assign \mchip.TPU.kernal_addr_x_counter.Q_next [1] = (_000_ ? _025_ : _023_);
	assign _026_ = \mchip.TPU.kernal_addr_x_counter.Q [1] & \mchip.TPU.kernal_addr_x_counter.Q [0];
	assign _027_ = _026_ ^ \mchip.TPU.kernal_addr_x_counter.Q [2];
	assign \mchip.TPU.kernal_addr_x_counter.Q_next [2] = _027_ & ~_024_;
	assign _028_ = ~(_026_ & \mchip.TPU.kernal_addr_x_counter.Q [2]);
	assign _029_ = ~(_028_ ^ \mchip.TPU.kernal_addr_x_counter.Q [3]);
	assign \mchip.TPU.kernal_addr_x_counter.Q_next [3] = _029_ & ~_024_;
	assign _030_ = ~\mchip.TPU.kernal_addr_y_counter.Q [0];
	assign _031_ = ~(\mchip.TPU.kernal_addr_y_counter.Q [2] | \mchip.TPU.kernal_addr_y_counter.Q [3]);
	assign _032_ = \mchip.TPU.kernal_addr_y_counter.Q [1] & ~\mchip.TPU.kernal_addr_y_counter.Q [0];
	assign _033_ = _032_ & _031_;
	assign \mchip.TPU.kernal_addr_y_counter.Q_next [0] = _030_ & ~_033_;
	assign _034_ = ~_031_;
	assign _035_ = \mchip.TPU.kernal_addr_y_counter.Q [0] & ~\mchip.TPU.kernal_addr_y_counter.Q [1];
	assign \mchip.TPU.kernal_addr_y_counter.Q_next [1] = (_032_ ? _034_ : _035_);
	assign _036_ = \mchip.TPU.kernal_addr_y_counter.Q [0] & \mchip.TPU.kernal_addr_y_counter.Q [1];
	assign _037_ = _036_ ^ \mchip.TPU.kernal_addr_y_counter.Q [2];
	assign \mchip.TPU.kernal_addr_y_counter.Q_next [2] = _037_ & ~_033_;
	assign _038_ = ~(_036_ & \mchip.TPU.kernal_addr_y_counter.Q [2]);
	assign _039_ = ~(_038_ ^ \mchip.TPU.kernal_addr_y_counter.Q [3]);
	assign \mchip.TPU.kernal_addr_y_counter.Q_next [3] = _039_ & ~_033_;
	assign _040_ = \mchip.TPU.base_addr_x_counter.Q [9] & \mchip.TPU.base_addr_x_counter.Q [8];
	assign _041_ = ~(\mchip.TPU.base_addr_x_counter.Q [6] & \mchip.TPU.base_addr_x_counter.Q [7]);
	assign _042_ = ~(\mchip.TPU.base_addr_x_counter.Q [5] & \mchip.TPU.base_addr_x_counter.Q [4]);
	assign _043_ = ~(_042_ | _041_);
	assign _044_ = ~(_043_ & _022_);
	assign _045_ = _044_ | ~_040_;
	assign \mchip.TPU.base_addr_x_counter.Q_next [0] = _045_ & ~\mchip.TPU.base_addr_x_counter.Q [0];
	assign \mchip.TPU.base_addr_x_counter.Q_next [1] = \mchip.TPU.base_addr_x_counter.Q [0] ^ \mchip.TPU.base_addr_x_counter.Q [1];
	assign _046_ = ~\mchip.TPU.base_addr_x_counter.Q [2];
	assign _047_ = _020_ ^ _046_;
	assign \mchip.TPU.base_addr_x_counter.Q_next [2] = _045_ & ~_047_;
	assign _048_ = ~(_020_ & \mchip.TPU.base_addr_x_counter.Q [2]);
	assign _049_ = _048_ ^ \mchip.TPU.base_addr_x_counter.Q [3];
	assign \mchip.TPU.base_addr_x_counter.Q_next [3] = _045_ & ~_049_;
	assign _050_ = _022_ ^ _019_;
	assign \mchip.TPU.base_addr_x_counter.Q_next [4] = _045_ & ~_050_;
	assign _051_ = ~(_017_ ^ \mchip.TPU.base_addr_x_counter.Q [5]);
	assign \mchip.TPU.base_addr_x_counter.Q_next [5] = _045_ & ~_051_;
	assign _052_ = _022_ & ~_042_;
	assign _053_ = ~(_052_ ^ \mchip.TPU.base_addr_x_counter.Q [6]);
	assign \mchip.TPU.base_addr_x_counter.Q_next [6] = _045_ & ~_053_;
	assign _054_ = ~(_052_ & \mchip.TPU.base_addr_x_counter.Q [6]);
	assign _055_ = _054_ ^ \mchip.TPU.base_addr_x_counter.Q [7];
	assign \mchip.TPU.base_addr_x_counter.Q_next [7] = _045_ & ~_055_;
	assign _056_ = _044_ ^ \mchip.TPU.base_addr_x_counter.Q [8];
	assign \mchip.TPU.base_addr_x_counter.Q_next [8] = _045_ & ~_056_;
	assign _057_ = _044_ | ~\mchip.TPU.base_addr_x_counter.Q [8];
	assign _058_ = _057_ ^ \mchip.TPU.base_addr_x_counter.Q [9];
	assign \mchip.TPU.base_addr_x_counter.Q_next [9] = _045_ & ~_058_;
	assign _059_ = \mchip.TPU.base_addr_y_counter.Q [9] & \mchip.TPU.base_addr_y_counter.Q [8];
	assign _060_ = \mchip.TPU.base_addr_y_counter.Q [0] & \mchip.TPU.base_addr_y_counter.Q [1];
	assign _061_ = \mchip.TPU.base_addr_y_counter.Q [2] & \mchip.TPU.base_addr_y_counter.Q [3];
	assign _062_ = _061_ & _060_;
	assign _063_ = ~(\mchip.TPU.base_addr_y_counter.Q [6] & \mchip.TPU.base_addr_y_counter.Q [7]);
	assign _064_ = ~(\mchip.TPU.base_addr_y_counter.Q [4] & \mchip.TPU.base_addr_y_counter.Q [5]);
	assign _065_ = ~(_064_ | _063_);
	assign _066_ = ~(_065_ & _062_);
	assign _067_ = _066_ | ~_059_;
	assign \mchip.TPU.base_addr_y_counter.Q_next [0] = _067_ & ~\mchip.TPU.base_addr_y_counter.Q [0];
	assign \mchip.TPU.base_addr_y_counter.Q_next [1] = \mchip.TPU.base_addr_y_counter.Q [0] ^ \mchip.TPU.base_addr_y_counter.Q [1];
	assign _068_ = ~\mchip.TPU.base_addr_y_counter.Q [2];
	assign _069_ = _060_ ^ _068_;
	assign \mchip.TPU.base_addr_y_counter.Q_next [2] = _067_ & ~_069_;
	assign _070_ = ~(_060_ & \mchip.TPU.base_addr_y_counter.Q [2]);
	assign _071_ = _070_ ^ \mchip.TPU.base_addr_y_counter.Q [3];
	assign \mchip.TPU.base_addr_y_counter.Q_next [3] = _067_ & ~_071_;
	assign _072_ = ~\mchip.TPU.base_addr_y_counter.Q [4];
	assign _073_ = _062_ ^ _072_;
	assign \mchip.TPU.base_addr_y_counter.Q_next [4] = _067_ & ~_073_;
	assign _074_ = ~(_062_ & \mchip.TPU.base_addr_y_counter.Q [4]);
	assign _075_ = _074_ ^ \mchip.TPU.base_addr_y_counter.Q [5];
	assign \mchip.TPU.base_addr_y_counter.Q_next [5] = _067_ & ~_075_;
	assign _076_ = _062_ & ~_064_;
	assign _077_ = ~(_076_ ^ \mchip.TPU.base_addr_y_counter.Q [6]);
	assign \mchip.TPU.base_addr_y_counter.Q_next [6] = _067_ & ~_077_;
	assign _078_ = ~(_076_ & \mchip.TPU.base_addr_y_counter.Q [6]);
	assign _079_ = _078_ ^ \mchip.TPU.base_addr_y_counter.Q [7];
	assign \mchip.TPU.base_addr_y_counter.Q_next [7] = _067_ & ~_079_;
	assign _080_ = _066_ ^ \mchip.TPU.base_addr_y_counter.Q [8];
	assign \mchip.TPU.base_addr_y_counter.Q_next [8] = _067_ & ~_080_;
	assign _081_ = _066_ | ~\mchip.TPU.base_addr_y_counter.Q [8];
	assign _082_ = _081_ ^ \mchip.TPU.base_addr_y_counter.Q [9];
	assign \mchip.TPU.base_addr_y_counter.Q_next [9] = _067_ & ~_082_;
	assign _083_ = ~\mchip.TPU.MATRIX_MAT.data [4];
	assign _084_ = ~\mchip.TPU.MATRIX_MAT.data [5];
	assign _085_ = ~\mchip.TPU.base_addr_x_counter.Q [0];
	assign _086_ = ~(\mchip.TPU.base_addr_x_counter.Q [0] ^ \mchip.TPU.kernal_addr_x_counter.Q [0]);
	assign _087_ = io_in[2] & ~io_in[0];
	assign _088_ = (_087_ ? _085_ : _086_);
	assign _089_ = (_088_ ? _083_ : _084_);
	assign _090_ = \mchip.TPU.base_addr_x_counter.Q [0] & \mchip.TPU.kernal_addr_x_counter.Q [0];
	assign _091_ = ~(\mchip.TPU.base_addr_x_counter.Q [1] ^ \mchip.TPU.kernal_addr_x_counter.Q [1]);
	assign _092_ = ~(_091_ ^ _090_);
	assign _093_ = (_087_ ? \mchip.TPU.base_addr_x_counter.Q [1] : _092_);
	assign _094_ = ~\mchip.TPU.MATRIX_MAT.data [6];
	assign _095_ = ~\mchip.TPU.MATRIX_MAT.data [7];
	assign _096_ = (_088_ ? _094_ : _095_);
	assign _097_ = (_093_ ? _096_ : _089_);
	assign _098_ = ~(\mchip.TPU.base_addr_x_counter.Q [1] & \mchip.TPU.kernal_addr_x_counter.Q [1]);
	assign _099_ = _090_ & ~_091_;
	assign _100_ = _098_ & ~_099_;
	assign _101_ = _100_ ^ _046_;
	assign _102_ = (_087_ ? \mchip.TPU.base_addr_x_counter.Q [2] : _101_);
	assign _103_ = ~\mchip.TPU.MATRIX_MAT.data [0];
	assign _104_ = ~\mchip.TPU.MATRIX_MAT.data [1];
	assign _105_ = (_088_ ? _103_ : _104_);
	assign _106_ = ~\mchip.TPU.MATRIX_MAT.data [2];
	assign _107_ = ~\mchip.TPU.MATRIX_MAT.data [3];
	assign _108_ = (_088_ ? _106_ : _107_);
	assign _109_ = (_093_ ? _108_ : _105_);
	assign _110_ = (_102_ ? _097_ : _109_);
	assign _111_ = ~\mchip.TPU.KERNAL_MAT.data [6];
	assign _112_ = ~\mchip.TPU.KERNAL_MAT.data [7];
	assign _113_ = \mchip.TPU.kernal_addr_y_counter.Q [0] ^ \mchip.TPU.kernal_addr_x_counter.Q [0];
	assign _114_ = (_113_ ? _112_ : _111_);
	assign _115_ = \mchip.TPU.kernal_addr_y_counter.Q [0] & \mchip.TPU.kernal_addr_x_counter.Q [0];
	assign _116_ = \mchip.TPU.kernal_addr_y_counter.Q [1] ^ \mchip.TPU.kernal_addr_x_counter.Q [1];
	assign _117_ = _116_ ^ \mchip.TPU.kernal_addr_y_counter.Q [0];
	assign _118_ = _117_ ^ _115_;
	assign _119_ = ~\mchip.TPU.KERNAL_MAT.data [4];
	assign _120_ = ~\mchip.TPU.KERNAL_MAT.data [5];
	assign _121_ = (_113_ ? _120_ : _119_);
	assign _122_ = (_118_ ? _114_ : _121_);
	assign _123_ = _117_ & _115_;
	assign _124_ = ~(\mchip.TPU.kernal_addr_y_counter.Q [1] & \mchip.TPU.kernal_addr_x_counter.Q [1]);
	assign _125_ = _116_ & ~_030_;
	assign _126_ = _124_ & ~_125_;
	assign _127_ = ~(_126_ ^ \mchip.TPU.kernal_addr_y_counter.Q [1]);
	assign _128_ = _127_ ^ _123_;
	assign _129_ = ~\mchip.TPU.KERNAL_MAT.data [2];
	assign _130_ = ~\mchip.TPU.KERNAL_MAT.data [3];
	assign _131_ = (_113_ ? _130_ : _129_);
	assign _132_ = ~\mchip.TPU.KERNAL_MAT.data [0];
	assign _133_ = ~\mchip.TPU.KERNAL_MAT.data [1];
	assign _134_ = (_113_ ? _133_ : _132_);
	assign _135_ = (_118_ ? _131_ : _134_);
	assign _136_ = (_128_ ? _122_ : _135_);
	assign _137_ = _136_ | _110_;
	assign _138_ = \mchip.TPU.conv_mac.sum_reg.Q [0] & ~_137_;
	assign \mchip.TPU.conv_mac.sum_reg.D [1] = _138_ ^ \mchip.TPU.conv_mac.sum_reg.Q [1];
	assign _139_ = _138_ & \mchip.TPU.conv_mac.sum_reg.Q [1];
	assign \mchip.TPU.conv_mac.sum_reg.D [2] = _139_ ^ \mchip.TPU.conv_mac.sum_reg.Q [2];
	assign _140_ = _139_ & \mchip.TPU.conv_mac.sum_reg.Q [2];
	assign \mchip.TPU.conv_mac.sum_reg.D [3] = _140_ ^ \mchip.TPU.conv_mac.sum_reg.Q [3];
	assign _141_ = ~(\mchip.TPU.conv_mac.sum_reg.Q [3] & \mchip.TPU.conv_mac.sum_reg.Q [2]);
	assign _142_ = _139_ & ~_141_;
	assign \mchip.TPU.conv_mac.sum_reg.D [4] = _142_ ^ \mchip.TPU.conv_mac.sum_reg.Q [4];
	assign _143_ = _142_ & \mchip.TPU.conv_mac.sum_reg.Q [4];
	assign \mchip.TPU.conv_mac.sum_reg.D [5] = _143_ ^ \mchip.TPU.conv_mac.sum_reg.Q [5];
	assign _144_ = ~(\mchip.TPU.conv_mac.sum_reg.Q [5] & \mchip.TPU.conv_mac.sum_reg.Q [4]);
	assign _145_ = _142_ & ~_144_;
	assign \mchip.TPU.conv_mac.sum_reg.D [6] = _145_ ^ \mchip.TPU.conv_mac.sum_reg.Q [6];
	assign _146_ = _145_ & \mchip.TPU.conv_mac.sum_reg.Q [6];
	assign \mchip.TPU.conv_mac.sum_reg.D [7] = _146_ ^ \mchip.TPU.conv_mac.sum_reg.Q [7];
	assign \mchip.TPU.conv_mac.sum_reg.D [0] = ~(_137_ ^ \mchip.TPU.conv_mac.sum_reg.Q [0]);
	assign \mchip.TPU.KERNAL_MAT.we  = io_in[1] & io_in[0];
	assign \mchip.TPU.MATRIX_MAT.we  = io_in[1] & ~io_in[0];
	assign _147_ = ~io_in[2];
	assign _148_ = ~(io_in[1] & io_in[2]);
	assign _149_ = _148_ | ~io_in[0];
	assign _150_ = io_in[3] & ~_149_;
	assign \mchip.TPU.kernal_addr_x_counter.en  = _150_ | _147_;
	assign _151_ = _148_ | io_in[0];
	assign _152_ = _147_ & ~_000_;
	assign _018_ = _151_ & ~_152_;
	assign _153_ = io_in[3] & ~_018_;
	assign \mchip.TPU.mac_rst  = _153_ | io_in[13];
	assign \mchip.TPU.done  = _153_ & ~io_in[13];
	assign _154_ = ~(\mchip.TPU.base_addr_y_counter.Q [1] & \mchip.TPU.kernal_addr_y_counter.Q [1]);
	assign _155_ = \mchip.TPU.base_addr_y_counter.Q [1] ^ \mchip.TPU.kernal_addr_y_counter.Q [1];
	assign _156_ = ~(\mchip.TPU.base_addr_y_counter.Q [0] & \mchip.TPU.kernal_addr_y_counter.Q [0]);
	assign _157_ = _155_ & ~_156_;
	assign _158_ = _154_ & ~_157_;
	assign _159_ = _061_ & ~_158_;
	assign _160_ = _159_ & ~_072_;
	assign _161_ = _021_ & ~_100_;
	assign _162_ = _161_ & ~_019_;
	assign _163_ = _162_ | _160_;
	assign \mchip.TPU.conv_mac.en  = _147_ & ~_163_;
	assign _164_ = ~_113_;
	assign _165_ = \mchip.TPU.kernal_addr_y_counter.Q [1] & ~_126_;
	assign _166_ = _127_ & _123_;
	assign _167_ = ~(_166_ | _165_);
	assign _168_ = _167_ & ~_128_;
	assign _169_ = _164_ & ~_118_;
	assign _170_ = ~_169_;
	assign _171_ = _168_ & ~_170_;
	assign _172_ = ~(_171_ & io_in[4]);
	assign _173_ = _164_ & ~_172_;
	assign _174_ = ~(_118_ & _113_);
	assign _175_ = _174_ & ~_169_;
	assign _176_ = _173_ & ~_175_;
	assign _177_ = _170_ ^ _128_;
	assign _178_ = _176_ & ~_177_;
	assign _179_ = _169_ & ~_128_;
	assign _180_ = ~(_179_ ^ _167_);
	assign _181_ = ~_180_;
	assign _182_ = _178_ & ~_181_;
	assign _183_ = ~(_171_ & _164_);
	assign _184_ = _183_ | _175_;
	assign _185_ = _184_ | _177_;
	assign _186_ = _180_ & ~_185_;
	assign _187_ = \mchip.TPU.KERNAL_MAT.data [0] & ~_186_;
	assign _001_ = _187_ | _182_;
	assign _188_ = ~(_113_ & io_in[4]);
	assign _189_ = _188_ | ~_175_;
	assign _190_ = _177_ & ~_189_;
	assign _191_ = _190_ & ~_180_;
	assign _192_ = _118_ | _164_;
	assign _193_ = _177_ & ~_192_;
	assign _194_ = _193_ & ~_180_;
	assign _195_ = \mchip.TPU.KERNAL_MAT.data [1] & ~_194_;
	assign _002_ = _195_ | _191_;
	assign _196_ = ~_177_;
	assign _197_ = ~io_in[4];
	assign _198_ = _171_ | _197_;
	assign _199_ = _198_ | _113_;
	assign _200_ = _199_ | ~_175_;
	assign _201_ = _200_ | _196_;
	assign _202_ = _181_ & ~_201_;
	assign _203_ = ~(_118_ & _164_);
	assign _204_ = _177_ & ~_203_;
	assign _205_ = _204_ & ~_180_;
	assign _206_ = \mchip.TPU.KERNAL_MAT.data [2] & ~_205_;
	assign _003_ = _206_ | _202_;
	assign _207_ = _188_ | _175_;
	assign _208_ = _177_ & ~_207_;
	assign _209_ = _208_ & ~_180_;
	assign _210_ = _177_ & ~_174_;
	assign _211_ = _210_ & ~_180_;
	assign _212_ = \mchip.TPU.KERNAL_MAT.data [3] & ~_211_;
	assign _004_ = _212_ | _209_;
	assign _213_ = _199_ | _175_;
	assign _214_ = _213_ | _196_;
	assign _215_ = _181_ & ~_214_;
	assign _216_ = _171_ | _113_;
	assign _217_ = _216_ | _175_;
	assign _218_ = _217_ | _196_;
	assign _219_ = _181_ & ~_218_;
	assign _220_ = \mchip.TPU.KERNAL_MAT.data [4] & ~_219_;
	assign _005_ = _220_ | _215_;
	assign _221_ = ~(_189_ | _177_);
	assign _222_ = _221_ & ~_180_;
	assign _223_ = ~(_192_ | _177_);
	assign _224_ = _223_ & ~_180_;
	assign _225_ = \mchip.TPU.KERNAL_MAT.data [5] & ~_224_;
	assign _006_ = _225_ | _222_;
	assign _226_ = _200_ | _177_;
	assign _227_ = _181_ & ~_226_;
	assign _228_ = ~(_203_ | _177_);
	assign _229_ = _228_ & ~_180_;
	assign _230_ = \mchip.TPU.KERNAL_MAT.data [6] & ~_229_;
	assign _007_ = _230_ | _227_;
	assign _231_ = ~(_207_ | _177_);
	assign _232_ = _231_ & ~_180_;
	assign _233_ = ~(_177_ | _174_);
	assign _234_ = _233_ & ~_180_;
	assign _235_ = \mchip.TPU.KERNAL_MAT.data [7] & ~_234_;
	assign _008_ = _235_ | _232_;
	assign _236_ = _088_ & ~_093_;
	assign _237_ = _236_ & ~_102_;
	assign _238_ = \mchip.TPU.base_addr_x_counter.Q [2] & ~_100_;
	assign _239_ = _238_ ^ \mchip.TPU.base_addr_x_counter.Q [3];
	assign _240_ = (_087_ ? \mchip.TPU.base_addr_x_counter.Q [3] : _239_);
	assign _241_ = ~(_240_ ^ _237_);
	assign _242_ = ~_241_;
	assign _243_ = ~_088_;
	assign _244_ = _240_ | _102_;
	assign _245_ = _236_ & ~_244_;
	assign _246_ = _161_ ^ \mchip.TPU.base_addr_x_counter.Q [4];
	assign _247_ = (_087_ ? \mchip.TPU.base_addr_x_counter.Q [4] : _246_);
	assign _248_ = ~(_247_ ^ _245_);
	assign _249_ = _158_ ^ _068_;
	assign _250_ = (_087_ ? \mchip.TPU.base_addr_y_counter.Q [2] : _249_);
	assign _251_ = ~(_156_ ^ _155_);
	assign _252_ = (_087_ ? \mchip.TPU.base_addr_y_counter.Q [1] : _251_);
	assign _253_ = _252_ | _250_;
	assign _254_ = ~\mchip.TPU.base_addr_y_counter.Q [0];
	assign _255_ = ~(\mchip.TPU.base_addr_y_counter.Q [0] ^ \mchip.TPU.kernal_addr_y_counter.Q [0]);
	assign _256_ = (_087_ ? _254_ : _255_);
	assign _257_ = _247_ | ~_256_;
	assign _258_ = _257_ | _253_;
	assign _259_ = _245_ & ~_258_;
	assign _260_ = \mchip.TPU.base_addr_y_counter.Q [2] & ~_158_;
	assign _261_ = _260_ ^ \mchip.TPU.base_addr_y_counter.Q [3];
	assign _262_ = (_087_ ? \mchip.TPU.base_addr_y_counter.Q [3] : _261_);
	assign _263_ = _259_ & ~_262_;
	assign _264_ = _159_ ^ _072_;
	assign _265_ = (_087_ ? _072_ : _264_);
	assign _266_ = _265_ ^ _263_;
	assign _267_ = _266_ ^ _248_;
	assign _268_ = ~(_262_ ^ _259_);
	assign _269_ = _268_ ^ _248_;
	assign _270_ = _245_ & ~_257_;
	assign _271_ = _270_ & ~_252_;
	assign _272_ = ~(_271_ ^ _250_);
	assign _273_ = _272_ ^ _248_;
	assign _274_ = ~(_270_ ^ _252_);
	assign _275_ = _274_ ^ _248_;
	assign _276_ = _245_ & ~_247_;
	assign _277_ = _256_ ^ _276_;
	assign _278_ = _277_ ^ _248_;
	assign _279_ = _278_ | _275_;
	assign _280_ = _279_ | _273_;
	assign _281_ = _280_ | _269_;
	assign _282_ = _281_ | _267_;
	assign _283_ = ~_248_;
	assign _284_ = _262_ | ~_265_;
	assign _285_ = _259_ & ~_284_;
	assign _286_ = _285_ ^ _283_;
	assign _287_ = _286_ | _282_;
	assign _288_ = _287_ | _197_;
	assign _289_ = _288_ | _248_;
	assign _290_ = _289_ | _243_;
	assign _291_ = _093_ ^ _243_;
	assign _292_ = _291_ | _290_;
	assign _293_ = ~(_236_ ^ _102_);
	assign _294_ = _293_ | _292_;
	assign _295_ = _242_ & ~_294_;
	assign _296_ = _287_ | _248_;
	assign _297_ = _296_ | _243_;
	assign _298_ = _297_ | _291_;
	assign _299_ = _298_ | _293_;
	assign _300_ = _242_ & ~_299_;
	assign _301_ = \mchip.TPU.MATRIX_MAT.data [0] & ~_300_;
	assign _009_ = _301_ | _295_;
	assign _302_ = ~_293_;
	assign _303_ = ~_291_;
	assign _304_ = _288_ | _283_;
	assign _305_ = _304_ | _088_;
	assign _306_ = _305_ | _303_;
	assign _307_ = _306_ | _302_;
	assign _308_ = _241_ & ~_307_;
	assign _309_ = _287_ | _283_;
	assign _310_ = _309_ | _088_;
	assign _311_ = _310_ | _303_;
	assign _312_ = _311_ | _302_;
	assign _313_ = _241_ & ~_312_;
	assign _314_ = \mchip.TPU.MATRIX_MAT.data [1] & ~_313_;
	assign _010_ = _314_ | _308_;
	assign _315_ = _304_ | _243_;
	assign _316_ = _315_ | _303_;
	assign _317_ = _316_ | _302_;
	assign _318_ = _241_ & ~_317_;
	assign _319_ = _309_ | _243_;
	assign _320_ = _319_ | _303_;
	assign _321_ = _320_ | _302_;
	assign _322_ = _241_ & ~_321_;
	assign _323_ = \mchip.TPU.MATRIX_MAT.data [2] & ~_322_;
	assign _011_ = _323_ | _318_;
	assign _324_ = _305_ | _291_;
	assign _325_ = _324_ | _302_;
	assign _326_ = _241_ & ~_325_;
	assign _327_ = _310_ | _291_;
	assign _328_ = _327_ | _302_;
	assign _329_ = _241_ & ~_328_;
	assign _330_ = \mchip.TPU.MATRIX_MAT.data [3] & ~_329_;
	assign _012_ = _330_ | _326_;
	assign _331_ = _315_ | _291_;
	assign _332_ = _331_ | _302_;
	assign _333_ = _241_ & ~_332_;
	assign _334_ = _319_ | _291_;
	assign _335_ = _334_ | _302_;
	assign _336_ = _241_ & ~_335_;
	assign _337_ = \mchip.TPU.MATRIX_MAT.data [4] & ~_336_;
	assign _013_ = _337_ | _333_;
	assign _338_ = _306_ | _293_;
	assign _339_ = _241_ & ~_338_;
	assign _340_ = _311_ | _293_;
	assign _341_ = _241_ & ~_340_;
	assign _342_ = \mchip.TPU.MATRIX_MAT.data [5] & ~_341_;
	assign _014_ = _342_ | _339_;
	assign _343_ = _316_ | _293_;
	assign _344_ = _241_ & ~_343_;
	assign _345_ = _320_ | _293_;
	assign _346_ = _241_ & ~_345_;
	assign _347_ = \mchip.TPU.MATRIX_MAT.data [6] & ~_346_;
	assign _015_ = _347_ | _344_;
	assign _348_ = _324_ | _293_;
	assign _349_ = _241_ & ~_348_;
	assign _350_ = _327_ | _293_;
	assign _351_ = _241_ & ~_350_;
	assign _352_ = \mchip.TPU.MATRIX_MAT.data [7] & ~_351_;
	assign _016_ = _352_ | _349_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.TPU.KERNAL_MAT.data [0] <= 1'h0;
		else if (\mchip.TPU.KERNAL_MAT.we )
			\mchip.TPU.KERNAL_MAT.data [0] <= _001_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.TPU.KERNAL_MAT.data [1] <= 1'h0;
		else if (\mchip.TPU.KERNAL_MAT.we )
			\mchip.TPU.KERNAL_MAT.data [1] <= _002_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.TPU.KERNAL_MAT.data [2] <= 1'h0;
		else if (\mchip.TPU.KERNAL_MAT.we )
			\mchip.TPU.KERNAL_MAT.data [2] <= _003_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.TPU.KERNAL_MAT.data [3] <= 1'h0;
		else if (\mchip.TPU.KERNAL_MAT.we )
			\mchip.TPU.KERNAL_MAT.data [3] <= _004_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.TPU.KERNAL_MAT.data [4] <= 1'h0;
		else if (\mchip.TPU.KERNAL_MAT.we )
			\mchip.TPU.KERNAL_MAT.data [4] <= _005_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.TPU.KERNAL_MAT.data [5] <= 1'h0;
		else if (\mchip.TPU.KERNAL_MAT.we )
			\mchip.TPU.KERNAL_MAT.data [5] <= _006_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.TPU.KERNAL_MAT.data [6] <= 1'h0;
		else if (\mchip.TPU.KERNAL_MAT.we )
			\mchip.TPU.KERNAL_MAT.data [6] <= _007_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.TPU.KERNAL_MAT.data [7] <= 1'h0;
		else if (\mchip.TPU.KERNAL_MAT.we )
			\mchip.TPU.KERNAL_MAT.data [7] <= _008_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.TPU.MATRIX_MAT.data [0] <= 1'h0;
		else if (\mchip.TPU.MATRIX_MAT.we )
			\mchip.TPU.MATRIX_MAT.data [0] <= _009_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.TPU.MATRIX_MAT.data [1] <= 1'h0;
		else if (\mchip.TPU.MATRIX_MAT.we )
			\mchip.TPU.MATRIX_MAT.data [1] <= _010_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.TPU.MATRIX_MAT.data [2] <= 1'h0;
		else if (\mchip.TPU.MATRIX_MAT.we )
			\mchip.TPU.MATRIX_MAT.data [2] <= _011_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.TPU.MATRIX_MAT.data [3] <= 1'h0;
		else if (\mchip.TPU.MATRIX_MAT.we )
			\mchip.TPU.MATRIX_MAT.data [3] <= _012_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.TPU.MATRIX_MAT.data [4] <= 1'h0;
		else if (\mchip.TPU.MATRIX_MAT.we )
			\mchip.TPU.MATRIX_MAT.data [4] <= _013_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.TPU.MATRIX_MAT.data [5] <= 1'h0;
		else if (\mchip.TPU.MATRIX_MAT.we )
			\mchip.TPU.MATRIX_MAT.data [5] <= _014_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.TPU.MATRIX_MAT.data [6] <= 1'h0;
		else if (\mchip.TPU.MATRIX_MAT.we )
			\mchip.TPU.MATRIX_MAT.data [6] <= _015_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.TPU.MATRIX_MAT.data [7] <= 1'h0;
		else if (\mchip.TPU.MATRIX_MAT.we )
			\mchip.TPU.MATRIX_MAT.data [7] <= _016_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.TPU.kernal_addr_x_counter.Q [0] <= 1'h0;
		else if (\mchip.TPU.kernal_addr_x_counter.en )
			\mchip.TPU.kernal_addr_x_counter.Q [0] <= \mchip.TPU.kernal_addr_x_counter.Q_next [0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.TPU.kernal_addr_x_counter.Q [1] <= 1'h0;
		else if (\mchip.TPU.kernal_addr_x_counter.en )
			\mchip.TPU.kernal_addr_x_counter.Q [1] <= \mchip.TPU.kernal_addr_x_counter.Q_next [1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.TPU.kernal_addr_x_counter.Q [2] <= 1'h0;
		else if (\mchip.TPU.kernal_addr_x_counter.en )
			\mchip.TPU.kernal_addr_x_counter.Q [2] <= \mchip.TPU.kernal_addr_x_counter.Q_next [2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.TPU.kernal_addr_x_counter.Q [3] <= 1'h0;
		else if (\mchip.TPU.kernal_addr_x_counter.en )
			\mchip.TPU.kernal_addr_x_counter.Q [3] <= \mchip.TPU.kernal_addr_x_counter.Q_next [3];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.TPU.kernal_addr_y_counter.Q [0] <= 1'h0;
		else if (!_000_)
			\mchip.TPU.kernal_addr_y_counter.Q [0] <= \mchip.TPU.kernal_addr_y_counter.Q_next [0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.TPU.kernal_addr_y_counter.Q [1] <= 1'h0;
		else if (!_000_)
			\mchip.TPU.kernal_addr_y_counter.Q [1] <= \mchip.TPU.kernal_addr_y_counter.Q_next [1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.TPU.kernal_addr_y_counter.Q [2] <= 1'h0;
		else if (!_000_)
			\mchip.TPU.kernal_addr_y_counter.Q [2] <= \mchip.TPU.kernal_addr_y_counter.Q_next [2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.TPU.kernal_addr_y_counter.Q [3] <= 1'h0;
		else if (!_000_)
			\mchip.TPU.kernal_addr_y_counter.Q [3] <= \mchip.TPU.kernal_addr_y_counter.Q_next [3];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.TPU.base_addr_x_counter.Q [0] <= 1'h0;
		else if (!_018_)
			\mchip.TPU.base_addr_x_counter.Q [0] <= \mchip.TPU.base_addr_x_counter.Q_next [0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.TPU.base_addr_x_counter.Q [1] <= 1'h0;
		else if (!_018_)
			\mchip.TPU.base_addr_x_counter.Q [1] <= \mchip.TPU.base_addr_x_counter.Q_next [1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.TPU.base_addr_x_counter.Q [2] <= 1'h0;
		else if (!_018_)
			\mchip.TPU.base_addr_x_counter.Q [2] <= \mchip.TPU.base_addr_x_counter.Q_next [2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.TPU.base_addr_x_counter.Q [3] <= 1'h0;
		else if (!_018_)
			\mchip.TPU.base_addr_x_counter.Q [3] <= \mchip.TPU.base_addr_x_counter.Q_next [3];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.TPU.base_addr_x_counter.Q [4] <= 1'h0;
		else if (!_018_)
			\mchip.TPU.base_addr_x_counter.Q [4] <= \mchip.TPU.base_addr_x_counter.Q_next [4];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.TPU.base_addr_x_counter.Q [5] <= 1'h0;
		else if (!_018_)
			\mchip.TPU.base_addr_x_counter.Q [5] <= \mchip.TPU.base_addr_x_counter.Q_next [5];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.TPU.base_addr_x_counter.Q [6] <= 1'h0;
		else if (!_018_)
			\mchip.TPU.base_addr_x_counter.Q [6] <= \mchip.TPU.base_addr_x_counter.Q_next [6];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.TPU.base_addr_x_counter.Q [7] <= 1'h0;
		else if (!_018_)
			\mchip.TPU.base_addr_x_counter.Q [7] <= \mchip.TPU.base_addr_x_counter.Q_next [7];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.TPU.base_addr_x_counter.Q [8] <= 1'h0;
		else if (!_018_)
			\mchip.TPU.base_addr_x_counter.Q [8] <= \mchip.TPU.base_addr_x_counter.Q_next [8];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.TPU.base_addr_x_counter.Q [9] <= 1'h0;
		else if (!_018_)
			\mchip.TPU.base_addr_x_counter.Q [9] <= \mchip.TPU.base_addr_x_counter.Q_next [9];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.TPU.base_addr_y_counter.Q [0] <= 1'h0;
		else if (_017_)
			\mchip.TPU.base_addr_y_counter.Q [0] <= \mchip.TPU.base_addr_y_counter.Q_next [0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.TPU.base_addr_y_counter.Q [1] <= 1'h0;
		else if (_017_)
			\mchip.TPU.base_addr_y_counter.Q [1] <= \mchip.TPU.base_addr_y_counter.Q_next [1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.TPU.base_addr_y_counter.Q [2] <= 1'h0;
		else if (_017_)
			\mchip.TPU.base_addr_y_counter.Q [2] <= \mchip.TPU.base_addr_y_counter.Q_next [2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.TPU.base_addr_y_counter.Q [3] <= 1'h0;
		else if (_017_)
			\mchip.TPU.base_addr_y_counter.Q [3] <= \mchip.TPU.base_addr_y_counter.Q_next [3];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.TPU.base_addr_y_counter.Q [4] <= 1'h0;
		else if (_017_)
			\mchip.TPU.base_addr_y_counter.Q [4] <= \mchip.TPU.base_addr_y_counter.Q_next [4];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.TPU.base_addr_y_counter.Q [5] <= 1'h0;
		else if (_017_)
			\mchip.TPU.base_addr_y_counter.Q [5] <= \mchip.TPU.base_addr_y_counter.Q_next [5];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.TPU.base_addr_y_counter.Q [6] <= 1'h0;
		else if (_017_)
			\mchip.TPU.base_addr_y_counter.Q [6] <= \mchip.TPU.base_addr_y_counter.Q_next [6];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.TPU.base_addr_y_counter.Q [7] <= 1'h0;
		else if (_017_)
			\mchip.TPU.base_addr_y_counter.Q [7] <= \mchip.TPU.base_addr_y_counter.Q_next [7];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.TPU.base_addr_y_counter.Q [8] <= 1'h0;
		else if (_017_)
			\mchip.TPU.base_addr_y_counter.Q [8] <= \mchip.TPU.base_addr_y_counter.Q_next [8];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.TPU.base_addr_y_counter.Q [9] <= 1'h0;
		else if (_017_)
			\mchip.TPU.base_addr_y_counter.Q [9] <= \mchip.TPU.base_addr_y_counter.Q_next [9];
	always @(posedge io_in[12])
		if (\mchip.TPU.mac_rst )
			\mchip.TPU.conv_mac.sum_reg.Q [0] <= 1'h0;
		else if (\mchip.TPU.conv_mac.en )
			\mchip.TPU.conv_mac.sum_reg.Q [0] <= \mchip.TPU.conv_mac.sum_reg.D [0];
	always @(posedge io_in[12])
		if (\mchip.TPU.mac_rst )
			\mchip.TPU.conv_mac.sum_reg.Q [1] <= 1'h0;
		else if (\mchip.TPU.conv_mac.en )
			\mchip.TPU.conv_mac.sum_reg.Q [1] <= \mchip.TPU.conv_mac.sum_reg.D [1];
	always @(posedge io_in[12])
		if (\mchip.TPU.mac_rst )
			\mchip.TPU.conv_mac.sum_reg.Q [2] <= 1'h0;
		else if (\mchip.TPU.conv_mac.en )
			\mchip.TPU.conv_mac.sum_reg.Q [2] <= \mchip.TPU.conv_mac.sum_reg.D [2];
	always @(posedge io_in[12])
		if (\mchip.TPU.mac_rst )
			\mchip.TPU.conv_mac.sum_reg.Q [3] <= 1'h0;
		else if (\mchip.TPU.conv_mac.en )
			\mchip.TPU.conv_mac.sum_reg.Q [3] <= \mchip.TPU.conv_mac.sum_reg.D [3];
	always @(posedge io_in[12])
		if (\mchip.TPU.mac_rst )
			\mchip.TPU.conv_mac.sum_reg.Q [4] <= 1'h0;
		else if (\mchip.TPU.conv_mac.en )
			\mchip.TPU.conv_mac.sum_reg.Q [4] <= \mchip.TPU.conv_mac.sum_reg.D [4];
	always @(posedge io_in[12])
		if (\mchip.TPU.mac_rst )
			\mchip.TPU.conv_mac.sum_reg.Q [5] <= 1'h0;
		else if (\mchip.TPU.conv_mac.en )
			\mchip.TPU.conv_mac.sum_reg.Q [5] <= \mchip.TPU.conv_mac.sum_reg.D [5];
	always @(posedge io_in[12])
		if (\mchip.TPU.mac_rst )
			\mchip.TPU.conv_mac.sum_reg.Q [6] <= 1'h0;
		else if (\mchip.TPU.conv_mac.en )
			\mchip.TPU.conv_mac.sum_reg.Q [6] <= \mchip.TPU.conv_mac.sum_reg.D [6];
	always @(posedge io_in[12])
		if (\mchip.TPU.mac_rst )
			\mchip.TPU.conv_mac.sum_reg.Q [7] <= 1'h0;
		else if (\mchip.TPU.conv_mac.en )
			\mchip.TPU.conv_mac.sum_reg.Q [7] <= \mchip.TPU.conv_mac.sum_reg.D [7];
	assign io_out = {2'h0, \mchip.TPU.conv_mac.sum_reg.Q , 3'h0, \mchip.TPU.done };
	assign \mchip.TPU.KERNAL_MAT.D  = io_in[11:4];
	assign \mchip.TPU.KERNAL_MAT.Q  = 8'h00;
	assign \mchip.TPU.KERNAL_MAT.clk  = io_in[12];
	assign \mchip.TPU.KERNAL_MAT.rst  = io_in[13];
	assign \mchip.TPU.MATRIX_MAT.D  = io_in[11:4];
	assign \mchip.TPU.MATRIX_MAT.Q  = 8'h00;
	assign \mchip.TPU.MATRIX_MAT.clk  = io_in[12];
	assign \mchip.TPU.MATRIX_MAT.rst  = io_in[13];
	assign \mchip.TPU.base_addr  = {\mchip.TPU.base_addr_x_counter.Q [4:0], \mchip.TPU.base_addr_y_counter.Q [4:0]};
	assign \mchip.TPU.base_addr_x_counter.clk  = io_in[12];
	assign \mchip.TPU.base_addr_x_counter.rst  = io_in[13];
	assign \mchip.TPU.base_addr_y_counter.clk  = io_in[12];
	assign \mchip.TPU.base_addr_y_counter.rst  = io_in[13];
	assign \mchip.TPU.clk  = io_in[12];
	assign \mchip.TPU.conv_mac.a  = 8'h00;
	assign \mchip.TPU.conv_mac.b  = 8'h00;
	assign \mchip.TPU.conv_mac.clk  = io_in[12];
	assign \mchip.TPU.conv_mac.new_sum  = \mchip.TPU.conv_mac.sum_reg.D ;
	assign \mchip.TPU.conv_mac.prod  = 8'h00;
	assign \mchip.TPU.conv_mac.rst  = \mchip.TPU.mac_rst ;
	assign \mchip.TPU.conv_mac.sum  = \mchip.TPU.conv_mac.sum_reg.Q ;
	assign \mchip.TPU.conv_mac.sum_reg.clk  = io_in[12];
	assign \mchip.TPU.conv_mac.sum_reg.rst  = \mchip.TPU.mac_rst ;
	assign \mchip.TPU.conv_mac.sum_reg.we  = \mchip.TPU.conv_mac.en ;
	assign \mchip.TPU.data_in  = io_in[11:4];
	assign \mchip.TPU.data_out  = \mchip.TPU.conv_mac.sum_reg.Q ;
	assign \mchip.TPU.insert_kernal  = io_in[0];
	assign \mchip.TPU.kernal_addr  = {\mchip.TPU.kernal_addr_x_counter.Q [1:0], \mchip.TPU.kernal_addr_y_counter.Q [1:0]};
	assign \mchip.TPU.kernal_addr_x_counter.clk  = io_in[12];
	assign \mchip.TPU.kernal_addr_x_counter.rst  = io_in[13];
	assign \mchip.TPU.kernal_addr_y_counter.clk  = io_in[12];
	assign \mchip.TPU.kernal_addr_y_counter.rst  = io_in[13];
	assign \mchip.TPU.kernal_data  = 8'h00;
	assign \mchip.TPU.kernal_x_incr  = \mchip.TPU.kernal_addr_x_counter.en ;
	assign \mchip.TPU.mac_en  = \mchip.TPU.conv_mac.en ;
	assign \mchip.TPU.matrix_data  = 8'h00;
	assign \mchip.TPU.ready  = io_in[3];
	assign \mchip.TPU.rst  = io_in[13];
	assign \mchip.TPU.write  = io_in[1];
	assign \mchip.TPU.write_mode  = io_in[2];
	assign \mchip.clock  = io_in[12];
	assign \mchip.io_in  = io_in[11:0];
	assign \mchip.io_out  = {\mchip.TPU.conv_mac.sum_reg.Q , 3'h0, \mchip.TPU.done };
	assign \mchip.reset  = io_in[13];
endmodule
module d25_araghave_huffman (
	io_in,
	io_out
);
	wire _0000_;
	wire _0001_;
	wire _0002_;
	wire _0003_;
	wire _0004_;
	wire _0005_;
	wire _0006_;
	wire _0007_;
	wire _0008_;
	wire _0009_;
	wire _0010_;
	wire _0011_;
	wire _0012_;
	wire _0013_;
	wire _0014_;
	wire _0015_;
	wire _0016_;
	wire _0017_;
	wire _0018_;
	wire _0019_;
	wire _0020_;
	wire _0021_;
	wire _0022_;
	wire _0023_;
	wire _0024_;
	wire _0025_;
	wire _0026_;
	wire _0027_;
	wire _0028_;
	wire _0029_;
	wire _0030_;
	wire _0031_;
	wire _0032_;
	wire _0033_;
	wire _0034_;
	wire _0035_;
	wire _0036_;
	wire _0037_;
	wire _0038_;
	wire _0039_;
	wire _0040_;
	wire _0041_;
	wire _0042_;
	wire _0043_;
	wire _0044_;
	wire _0045_;
	wire _0046_;
	wire _0047_;
	wire _0048_;
	wire _0049_;
	wire _0050_;
	wire _0051_;
	wire _0052_;
	wire _0053_;
	wire _0054_;
	wire _0055_;
	wire _0056_;
	wire _0057_;
	wire _0058_;
	wire _0059_;
	wire _0060_;
	wire _0061_;
	wire _0062_;
	wire _0063_;
	wire _0064_;
	wire _0065_;
	wire _0066_;
	wire _0067_;
	wire _0068_;
	wire _0069_;
	wire _0070_;
	wire _0071_;
	wire _0072_;
	wire _0073_;
	wire _0074_;
	wire _0075_;
	wire _0076_;
	wire _0077_;
	wire _0078_;
	wire _0079_;
	wire _0080_;
	wire _0081_;
	wire _0082_;
	wire _0083_;
	wire _0084_;
	wire _0085_;
	wire _0086_;
	wire _0087_;
	wire _0088_;
	wire _0089_;
	wire _0090_;
	wire _0091_;
	wire _0092_;
	wire _0093_;
	wire _0094_;
	wire _0095_;
	wire _0096_;
	wire _0097_;
	wire _0098_;
	wire _0099_;
	wire _0100_;
	wire _0101_;
	wire _0102_;
	wire _0103_;
	wire _0104_;
	wire _0105_;
	wire _0106_;
	wire _0107_;
	wire _0108_;
	wire _0109_;
	wire _0110_;
	wire _0111_;
	wire _0112_;
	wire _0113_;
	wire _0114_;
	wire _0115_;
	wire _0116_;
	wire _0117_;
	wire _0118_;
	wire _0119_;
	wire _0120_;
	wire _0121_;
	wire _0122_;
	wire _0123_;
	wire _0124_;
	wire _0125_;
	wire _0126_;
	wire _0127_;
	wire _0128_;
	wire _0129_;
	wire _0130_;
	wire _0131_;
	wire _0132_;
	wire _0133_;
	wire _0134_;
	wire _0135_;
	wire _0136_;
	wire _0137_;
	wire _0138_;
	wire _0139_;
	wire _0140_;
	wire _0141_;
	wire _0142_;
	wire _0143_;
	wire _0144_;
	wire _0145_;
	wire _0146_;
	wire _0147_;
	wire _0148_;
	wire _0149_;
	wire _0150_;
	wire _0151_;
	wire _0152_;
	wire _0153_;
	wire _0154_;
	wire _0155_;
	wire _0156_;
	wire _0157_;
	wire _0158_;
	wire _0159_;
	wire _0160_;
	wire _0161_;
	wire _0162_;
	wire _0163_;
	wire _0164_;
	wire _0165_;
	wire _0166_;
	wire _0167_;
	wire _0168_;
	wire _0169_;
	wire _0170_;
	wire _0171_;
	wire _0172_;
	wire _0173_;
	wire _0174_;
	wire _0175_;
	wire _0176_;
	wire _0177_;
	wire _0178_;
	wire _0179_;
	wire _0180_;
	wire _0181_;
	wire _0182_;
	wire _0183_;
	wire _0184_;
	wire _0185_;
	wire _0186_;
	wire _0187_;
	wire _0188_;
	wire _0189_;
	wire _0190_;
	wire _0191_;
	wire _0192_;
	wire _0193_;
	wire _0194_;
	wire _0195_;
	wire _0196_;
	wire _0197_;
	wire _0198_;
	wire _0199_;
	wire _0200_;
	wire _0201_;
	wire _0202_;
	wire _0203_;
	wire _0204_;
	wire _0205_;
	wire _0206_;
	wire _0207_;
	wire _0208_;
	wire _0209_;
	wire _0210_;
	wire _0211_;
	wire _0212_;
	wire _0213_;
	wire _0214_;
	wire _0215_;
	wire _0216_;
	wire _0217_;
	wire _0218_;
	wire _0219_;
	wire _0220_;
	wire _0221_;
	wire _0222_;
	wire _0223_;
	wire _0224_;
	wire _0225_;
	wire _0226_;
	wire _0227_;
	wire _0228_;
	wire _0229_;
	wire _0230_;
	wire _0231_;
	wire _0232_;
	wire _0233_;
	wire _0234_;
	wire _0235_;
	wire _0236_;
	wire _0237_;
	wire _0238_;
	wire _0239_;
	wire _0240_;
	wire _0241_;
	wire _0242_;
	wire _0243_;
	wire _0244_;
	wire _0245_;
	wire _0246_;
	wire _0247_;
	wire _0248_;
	wire _0249_;
	wire _0250_;
	wire _0251_;
	wire _0252_;
	wire _0253_;
	wire _0254_;
	wire _0255_;
	wire _0256_;
	wire _0257_;
	wire _0258_;
	wire _0259_;
	wire _0260_;
	wire _0261_;
	wire _0262_;
	wire _0263_;
	wire _0264_;
	wire _0265_;
	wire _0266_;
	wire _0267_;
	wire _0268_;
	wire _0269_;
	wire _0270_;
	wire _0271_;
	wire _0272_;
	wire _0273_;
	wire _0274_;
	wire _0275_;
	wire _0276_;
	wire _0277_;
	wire _0278_;
	wire _0279_;
	wire _0280_;
	wire _0281_;
	wire _0282_;
	wire _0283_;
	wire _0284_;
	wire _0285_;
	wire _0286_;
	wire _0287_;
	wire _0288_;
	wire _0289_;
	wire _0290_;
	wire _0291_;
	wire _0292_;
	wire _0293_;
	wire _0294_;
	wire _0295_;
	wire _0296_;
	wire _0297_;
	wire _0298_;
	wire _0299_;
	wire _0300_;
	wire _0301_;
	wire _0302_;
	wire _0303_;
	wire _0304_;
	wire _0305_;
	wire _0306_;
	wire _0307_;
	wire _0308_;
	wire _0309_;
	wire _0310_;
	wire _0311_;
	wire _0312_;
	wire _0313_;
	wire _0314_;
	wire _0315_;
	wire _0316_;
	wire _0317_;
	wire _0318_;
	wire _0319_;
	wire _0320_;
	wire _0321_;
	wire _0322_;
	wire _0323_;
	wire _0324_;
	wire _0325_;
	wire _0326_;
	wire _0327_;
	wire _0328_;
	wire _0329_;
	wire _0330_;
	wire _0331_;
	wire _0332_;
	wire _0333_;
	wire _0334_;
	wire _0335_;
	wire _0336_;
	wire _0337_;
	wire _0338_;
	wire _0339_;
	wire _0340_;
	wire _0341_;
	wire _0342_;
	wire _0343_;
	wire _0344_;
	wire _0345_;
	wire _0346_;
	wire _0347_;
	wire _0348_;
	wire _0349_;
	wire _0350_;
	wire _0351_;
	wire _0352_;
	wire _0353_;
	wire _0354_;
	wire _0355_;
	wire _0356_;
	wire _0357_;
	wire _0358_;
	wire _0359_;
	wire _0360_;
	wire _0361_;
	wire _0362_;
	wire _0363_;
	wire _0364_;
	wire _0365_;
	wire _0366_;
	wire _0367_;
	wire _0368_;
	wire _0369_;
	wire _0370_;
	wire _0371_;
	wire _0372_;
	wire _0373_;
	wire _0374_;
	wire _0375_;
	wire _0376_;
	wire _0377_;
	wire _0378_;
	wire _0379_;
	wire _0380_;
	wire _0381_;
	wire _0382_;
	wire _0383_;
	wire _0384_;
	wire _0385_;
	wire _0386_;
	wire _0387_;
	wire _0388_;
	wire _0389_;
	wire _0390_;
	wire _0391_;
	wire _0392_;
	wire _0393_;
	wire _0394_;
	wire _0395_;
	wire _0396_;
	wire _0397_;
	wire _0398_;
	wire _0399_;
	wire _0400_;
	wire _0401_;
	wire _0402_;
	wire _0403_;
	wire _0404_;
	wire _0405_;
	wire _0406_;
	wire _0407_;
	wire _0408_;
	wire _0409_;
	wire _0410_;
	wire _0411_;
	wire _0412_;
	wire _0413_;
	wire _0414_;
	wire _0415_;
	wire _0416_;
	wire _0417_;
	wire _0418_;
	wire _0419_;
	wire _0420_;
	wire _0421_;
	wire _0422_;
	wire _0423_;
	wire _0424_;
	wire _0425_;
	wire _0426_;
	wire _0427_;
	wire _0428_;
	wire _0429_;
	wire _0430_;
	wire _0431_;
	wire _0432_;
	wire _0433_;
	wire _0434_;
	wire _0435_;
	wire _0436_;
	wire _0437_;
	wire _0438_;
	wire _0439_;
	wire _0440_;
	wire _0441_;
	wire _0442_;
	wire _0443_;
	wire _0444_;
	wire _0445_;
	wire _0446_;
	wire _0447_;
	wire _0448_;
	wire _0449_;
	wire _0450_;
	wire _0451_;
	wire _0452_;
	wire _0453_;
	wire _0454_;
	wire _0455_;
	wire _0456_;
	wire _0457_;
	wire _0458_;
	wire _0459_;
	wire _0460_;
	wire _0461_;
	wire _0462_;
	wire _0463_;
	wire _0464_;
	wire _0465_;
	wire _0466_;
	wire _0467_;
	wire _0468_;
	wire _0469_;
	wire _0470_;
	wire _0471_;
	wire _0472_;
	wire _0473_;
	wire _0474_;
	wire _0475_;
	wire _0476_;
	wire _0477_;
	wire _0478_;
	wire _0479_;
	wire _0480_;
	wire _0481_;
	wire _0482_;
	wire _0483_;
	wire _0484_;
	wire _0485_;
	wire _0486_;
	wire _0487_;
	wire _0488_;
	wire _0489_;
	wire _0490_;
	wire _0491_;
	wire _0492_;
	wire _0493_;
	wire _0494_;
	wire _0495_;
	wire _0496_;
	wire _0497_;
	wire _0498_;
	wire _0499_;
	wire _0500_;
	wire _0501_;
	wire _0502_;
	wire _0503_;
	wire _0504_;
	wire _0505_;
	wire _0506_;
	wire _0507_;
	wire _0508_;
	wire _0509_;
	wire _0510_;
	wire _0511_;
	wire _0512_;
	wire _0513_;
	wire _0514_;
	wire _0515_;
	wire _0516_;
	wire _0517_;
	wire _0518_;
	wire _0519_;
	wire _0520_;
	wire _0521_;
	wire _0522_;
	wire _0523_;
	wire _0524_;
	wire _0525_;
	wire _0526_;
	wire _0527_;
	wire _0528_;
	wire _0529_;
	wire _0530_;
	wire _0531_;
	wire _0532_;
	wire _0533_;
	wire _0534_;
	wire _0535_;
	wire _0536_;
	wire _0537_;
	wire _0538_;
	wire _0539_;
	wire _0540_;
	wire _0541_;
	wire _0542_;
	wire _0543_;
	wire _0544_;
	wire _0545_;
	wire _0546_;
	wire _0547_;
	wire _0548_;
	wire _0549_;
	wire _0550_;
	wire _0551_;
	wire _0552_;
	wire _0553_;
	wire _0554_;
	wire _0555_;
	wire _0556_;
	wire _0557_;
	wire _0558_;
	wire _0559_;
	wire _0560_;
	wire _0561_;
	wire _0562_;
	wire _0563_;
	wire _0564_;
	wire _0565_;
	wire _0566_;
	wire _0567_;
	wire _0568_;
	wire _0569_;
	wire _0570_;
	wire _0571_;
	wire _0572_;
	wire _0573_;
	wire _0574_;
	wire _0575_;
	wire _0576_;
	wire _0577_;
	wire _0578_;
	wire _0579_;
	wire _0580_;
	wire _0581_;
	wire _0582_;
	wire _0583_;
	wire _0584_;
	wire _0585_;
	wire _0586_;
	wire _0587_;
	wire _0588_;
	wire _0589_;
	wire _0590_;
	wire _0591_;
	wire _0592_;
	wire _0593_;
	wire _0594_;
	wire _0595_;
	wire _0596_;
	wire _0597_;
	wire _0598_;
	wire _0599_;
	wire _0600_;
	wire _0601_;
	wire _0602_;
	wire _0603_;
	wire _0604_;
	wire _0605_;
	wire _0606_;
	wire _0607_;
	wire _0608_;
	wire _0609_;
	wire _0610_;
	wire _0611_;
	wire _0612_;
	wire _0613_;
	wire _0614_;
	wire _0615_;
	wire _0616_;
	wire _0617_;
	wire _0618_;
	wire _0619_;
	wire _0620_;
	wire _0621_;
	wire _0622_;
	wire _0623_;
	wire _0624_;
	wire _0625_;
	wire _0626_;
	wire _0627_;
	wire _0628_;
	wire _0629_;
	wire _0630_;
	wire _0631_;
	wire _0632_;
	wire _0633_;
	wire _0634_;
	wire _0635_;
	wire _0636_;
	wire _0637_;
	wire _0638_;
	wire _0639_;
	wire _0640_;
	wire _0641_;
	wire _0642_;
	wire _0643_;
	wire _0644_;
	wire _0645_;
	wire _0646_;
	wire _0647_;
	wire _0648_;
	wire _0649_;
	wire _0650_;
	wire _0651_;
	wire _0652_;
	wire _0653_;
	wire _0654_;
	wire _0655_;
	wire _0656_;
	wire _0657_;
	wire _0658_;
	wire _0659_;
	wire _0660_;
	wire _0661_;
	wire _0662_;
	wire _0663_;
	wire _0664_;
	wire _0665_;
	wire _0666_;
	wire _0667_;
	wire _0668_;
	wire _0669_;
	wire _0670_;
	wire _0671_;
	wire _0672_;
	wire _0673_;
	wire _0674_;
	wire _0675_;
	wire _0676_;
	wire _0677_;
	wire _0678_;
	wire _0679_;
	wire _0680_;
	wire _0681_;
	wire _0682_;
	wire _0683_;
	wire _0684_;
	wire _0685_;
	wire _0686_;
	wire _0687_;
	wire _0688_;
	wire _0689_;
	wire _0690_;
	wire _0691_;
	wire _0692_;
	wire _0693_;
	wire _0694_;
	wire _0695_;
	wire _0696_;
	wire _0697_;
	wire _0698_;
	wire _0699_;
	wire _0700_;
	wire _0701_;
	wire _0702_;
	wire _0703_;
	wire _0704_;
	wire _0705_;
	wire _0706_;
	wire _0707_;
	wire _0708_;
	wire _0709_;
	wire _0710_;
	wire _0711_;
	wire _0712_;
	wire _0713_;
	wire _0714_;
	wire _0715_;
	wire _0716_;
	wire _0717_;
	wire _0718_;
	wire _0719_;
	wire _0720_;
	wire _0721_;
	wire _0722_;
	wire _0723_;
	wire _0724_;
	wire _0725_;
	wire _0726_;
	wire _0727_;
	wire _0728_;
	wire _0729_;
	wire _0730_;
	wire _0731_;
	wire _0732_;
	wire _0733_;
	wire _0734_;
	wire _0735_;
	wire _0736_;
	wire _0737_;
	wire _0738_;
	wire _0739_;
	wire _0740_;
	wire _0741_;
	wire _0742_;
	wire _0743_;
	wire _0744_;
	wire _0745_;
	wire _0746_;
	wire _0747_;
	wire _0748_;
	wire _0749_;
	wire _0750_;
	wire _0751_;
	wire _0752_;
	wire _0753_;
	wire _0754_;
	wire _0755_;
	wire _0756_;
	wire _0757_;
	wire _0758_;
	wire _0759_;
	wire _0760_;
	wire _0761_;
	wire _0762_;
	wire _0763_;
	wire _0764_;
	wire _0765_;
	wire _0766_;
	wire _0767_;
	wire _0768_;
	wire _0769_;
	wire _0770_;
	wire _0771_;
	wire _0772_;
	wire _0773_;
	wire _0774_;
	wire _0775_;
	wire _0776_;
	wire _0777_;
	wire _0778_;
	wire _0779_;
	wire _0780_;
	wire _0781_;
	wire _0782_;
	wire _0783_;
	wire _0784_;
	wire _0785_;
	wire _0786_;
	wire _0787_;
	wire _0788_;
	wire _0789_;
	wire _0790_;
	wire _0791_;
	wire _0792_;
	wire _0793_;
	wire _0794_;
	wire _0795_;
	wire _0796_;
	wire _0797_;
	wire _0798_;
	wire _0799_;
	wire _0800_;
	wire _0801_;
	wire _0802_;
	wire _0803_;
	wire _0804_;
	wire _0805_;
	wire _0806_;
	wire _0807_;
	wire _0808_;
	wire _0809_;
	wire _0810_;
	wire _0811_;
	wire _0812_;
	wire _0813_;
	wire _0814_;
	wire _0815_;
	wire _0816_;
	wire _0817_;
	wire _0818_;
	wire _0819_;
	wire _0820_;
	wire _0821_;
	wire _0822_;
	wire _0823_;
	wire _0824_;
	wire _0825_;
	wire _0826_;
	wire _0827_;
	wire _0828_;
	wire _0829_;
	wire _0830_;
	wire _0831_;
	wire _0832_;
	wire _0833_;
	wire _0834_;
	wire _0835_;
	wire _0836_;
	wire _0837_;
	wire _0838_;
	wire _0839_;
	wire _0840_;
	wire _0841_;
	wire _0842_;
	wire _0843_;
	wire _0844_;
	wire _0845_;
	wire _0846_;
	wire _0847_;
	wire _0848_;
	wire _0849_;
	wire _0850_;
	wire _0851_;
	wire _0852_;
	wire _0853_;
	wire _0854_;
	wire _0855_;
	wire _0856_;
	wire _0857_;
	wire _0858_;
	wire _0859_;
	wire _0860_;
	wire _0861_;
	wire _0862_;
	wire _0863_;
	wire _0864_;
	wire _0865_;
	wire _0866_;
	wire _0867_;
	wire _0868_;
	wire _0869_;
	wire _0870_;
	wire _0871_;
	wire _0872_;
	wire _0873_;
	wire _0874_;
	wire _0875_;
	wire _0876_;
	wire _0877_;
	wire _0878_;
	wire _0879_;
	wire _0880_;
	wire _0881_;
	wire _0882_;
	wire _0883_;
	wire _0884_;
	wire _0885_;
	wire _0886_;
	wire _0887_;
	wire _0888_;
	wire _0889_;
	wire _0890_;
	wire _0891_;
	wire _0892_;
	wire _0893_;
	wire _0894_;
	wire _0895_;
	wire _0896_;
	wire _0897_;
	wire _0898_;
	wire _0899_;
	wire _0900_;
	wire _0901_;
	wire _0902_;
	wire _0903_;
	wire _0904_;
	wire _0905_;
	wire _0906_;
	wire _0907_;
	wire _0908_;
	wire _0909_;
	wire _0910_;
	wire _0911_;
	wire _0912_;
	wire _0913_;
	wire _0914_;
	wire _0915_;
	wire _0916_;
	wire _0917_;
	wire _0918_;
	wire _0919_;
	wire _0920_;
	wire _0921_;
	wire _0922_;
	wire _0923_;
	wire _0924_;
	wire _0925_;
	wire _0926_;
	wire _0927_;
	wire _0928_;
	wire _0929_;
	wire _0930_;
	wire _0931_;
	wire _0932_;
	wire _0933_;
	wire _0934_;
	wire _0935_;
	wire _0936_;
	wire _0937_;
	wire _0938_;
	wire _0939_;
	wire _0940_;
	wire _0941_;
	wire _0942_;
	wire _0943_;
	wire _0944_;
	wire _0945_;
	wire _0946_;
	wire _0947_;
	wire _0948_;
	wire _0949_;
	wire _0950_;
	wire _0951_;
	wire _0952_;
	wire _0953_;
	wire _0954_;
	wire _0955_;
	wire _0956_;
	wire _0957_;
	wire _0958_;
	wire _0959_;
	wire _0960_;
	wire _0961_;
	wire _0962_;
	wire _0963_;
	wire _0964_;
	wire _0965_;
	wire _0966_;
	wire _0967_;
	wire _0968_;
	wire _0969_;
	wire _0970_;
	wire _0971_;
	wire _0972_;
	wire _0973_;
	wire _0974_;
	wire _0975_;
	wire _0976_;
	wire _0977_;
	wire _0978_;
	wire _0979_;
	wire _0980_;
	wire _0981_;
	wire _0982_;
	wire _0983_;
	wire _0984_;
	wire _0985_;
	wire _0986_;
	wire _0987_;
	wire _0988_;
	wire _0989_;
	wire _0990_;
	wire _0991_;
	wire _0992_;
	wire _0993_;
	wire _0994_;
	wire _0995_;
	wire _0996_;
	wire _0997_;
	wire _0998_;
	wire _0999_;
	wire _1000_;
	wire _1001_;
	wire _1002_;
	wire _1003_;
	wire _1004_;
	wire _1005_;
	wire _1006_;
	wire _1007_;
	wire _1008_;
	wire _1009_;
	wire _1010_;
	wire _1011_;
	wire _1012_;
	wire _1013_;
	wire _1014_;
	wire _1015_;
	wire _1016_;
	wire _1017_;
	wire _1018_;
	wire _1019_;
	wire _1020_;
	wire _1021_;
	wire _1022_;
	wire _1023_;
	wire _1024_;
	wire _1025_;
	wire _1026_;
	wire _1027_;
	wire _1028_;
	wire _1029_;
	wire _1030_;
	wire _1031_;
	wire _1032_;
	wire _1033_;
	wire _1034_;
	wire _1035_;
	wire _1036_;
	wire _1037_;
	wire _1038_;
	wire _1039_;
	wire _1040_;
	wire _1041_;
	wire _1042_;
	wire _1043_;
	wire _1044_;
	wire _1045_;
	wire _1046_;
	wire _1047_;
	wire _1048_;
	wire _1049_;
	wire _1050_;
	wire _1051_;
	wire _1052_;
	wire _1053_;
	wire _1054_;
	wire _1055_;
	wire _1056_;
	wire _1057_;
	wire _1058_;
	wire _1059_;
	wire _1060_;
	wire _1061_;
	wire _1062_;
	wire _1063_;
	wire _1064_;
	wire _1065_;
	wire _1066_;
	wire _1067_;
	wire _1068_;
	wire _1069_;
	wire _1070_;
	wire _1071_;
	wire _1072_;
	wire _1073_;
	wire _1074_;
	wire _1075_;
	wire _1076_;
	wire _1077_;
	wire _1078_;
	wire _1079_;
	wire _1080_;
	wire _1081_;
	wire _1082_;
	wire _1083_;
	wire _1084_;
	wire _1085_;
	wire _1086_;
	wire _1087_;
	wire _1088_;
	wire _1089_;
	wire _1090_;
	wire _1091_;
	wire _1092_;
	wire _1093_;
	wire _1094_;
	wire _1095_;
	wire _1096_;
	wire _1097_;
	wire _1098_;
	wire _1099_;
	wire _1100_;
	wire _1101_;
	wire _1102_;
	wire _1103_;
	wire _1104_;
	wire _1105_;
	wire _1106_;
	wire _1107_;
	wire _1108_;
	wire _1109_;
	wire _1110_;
	wire _1111_;
	wire _1112_;
	wire _1113_;
	wire _1114_;
	wire _1115_;
	wire _1116_;
	wire _1117_;
	wire _1118_;
	wire _1119_;
	wire _1120_;
	wire _1121_;
	wire _1122_;
	wire _1123_;
	wire _1124_;
	wire _1125_;
	wire _1126_;
	wire _1127_;
	wire _1128_;
	wire _1129_;
	wire _1130_;
	wire _1131_;
	wire _1132_;
	wire _1133_;
	wire _1134_;
	wire _1135_;
	wire _1136_;
	wire _1137_;
	wire _1138_;
	wire _1139_;
	wire _1140_;
	wire _1141_;
	wire _1142_;
	wire _1143_;
	wire _1144_;
	wire _1145_;
	wire _1146_;
	wire _1147_;
	wire _1148_;
	wire _1149_;
	wire _1150_;
	wire _1151_;
	wire _1152_;
	wire _1153_;
	wire _1154_;
	wire _1155_;
	wire _1156_;
	wire _1157_;
	wire _1158_;
	wire _1159_;
	wire _1160_;
	wire _1161_;
	wire _1162_;
	wire _1163_;
	wire _1164_;
	wire _1165_;
	wire _1166_;
	wire _1167_;
	wire _1168_;
	wire _1169_;
	wire _1170_;
	wire _1171_;
	wire _1172_;
	wire _1173_;
	wire _1174_;
	wire _1175_;
	wire _1176_;
	wire _1177_;
	wire _1178_;
	wire _1179_;
	wire _1180_;
	wire _1181_;
	wire _1182_;
	wire _1183_;
	wire _1184_;
	wire _1185_;
	wire _1186_;
	wire _1187_;
	wire _1188_;
	wire _1189_;
	wire _1190_;
	wire _1191_;
	wire _1192_;
	wire _1193_;
	wire _1194_;
	wire _1195_;
	wire _1196_;
	wire _1197_;
	wire _1198_;
	wire _1199_;
	wire _1200_;
	wire _1201_;
	wire _1202_;
	wire _1203_;
	wire _1204_;
	wire _1205_;
	wire _1206_;
	wire _1207_;
	wire _1208_;
	wire _1209_;
	wire _1210_;
	wire _1211_;
	wire _1212_;
	wire _1213_;
	wire _1214_;
	wire _1215_;
	wire _1216_;
	wire _1217_;
	wire _1218_;
	wire _1219_;
	wire _1220_;
	wire _1221_;
	wire _1222_;
	wire _1223_;
	wire _1224_;
	wire _1225_;
	wire _1226_;
	wire _1227_;
	wire _1228_;
	wire _1229_;
	wire _1230_;
	wire _1231_;
	wire _1232_;
	wire _1233_;
	wire _1234_;
	wire _1235_;
	wire _1236_;
	wire _1237_;
	wire _1238_;
	wire _1239_;
	wire _1240_;
	wire _1241_;
	wire _1242_;
	wire _1243_;
	wire _1244_;
	wire _1245_;
	wire _1246_;
	wire _1247_;
	wire _1248_;
	wire _1249_;
	wire _1250_;
	wire _1251_;
	wire _1252_;
	wire _1253_;
	wire _1254_;
	wire _1255_;
	wire _1256_;
	wire _1257_;
	wire _1258_;
	wire _1259_;
	wire _1260_;
	wire _1261_;
	wire _1262_;
	wire _1263_;
	wire _1264_;
	wire _1265_;
	wire _1266_;
	wire _1267_;
	wire _1268_;
	wire _1269_;
	wire _1270_;
	wire _1271_;
	wire _1272_;
	wire _1273_;
	wire _1274_;
	wire _1275_;
	wire _1276_;
	wire _1277_;
	wire _1278_;
	wire _1279_;
	wire _1280_;
	wire _1281_;
	wire _1282_;
	wire _1283_;
	wire _1284_;
	wire _1285_;
	wire _1286_;
	wire _1287_;
	wire _1288_;
	wire _1289_;
	wire _1290_;
	wire _1291_;
	wire _1292_;
	wire _1293_;
	wire _1294_;
	wire _1295_;
	wire _1296_;
	wire _1297_;
	wire _1298_;
	wire _1299_;
	wire _1300_;
	wire _1301_;
	wire _1302_;
	wire _1303_;
	wire _1304_;
	wire _1305_;
	wire _1306_;
	wire _1307_;
	wire _1308_;
	wire _1309_;
	wire _1310_;
	wire _1311_;
	wire _1312_;
	wire _1313_;
	wire _1314_;
	wire _1315_;
	wire _1316_;
	wire _1317_;
	wire _1318_;
	wire _1319_;
	wire _1320_;
	wire _1321_;
	wire _1322_;
	wire _1323_;
	wire _1324_;
	wire _1325_;
	wire _1326_;
	wire _1327_;
	wire _1328_;
	wire _1329_;
	wire _1330_;
	wire _1331_;
	wire _1332_;
	wire _1333_;
	wire _1334_;
	wire _1335_;
	wire _1336_;
	wire _1337_;
	wire _1338_;
	wire _1339_;
	wire _1340_;
	wire _1341_;
	wire _1342_;
	wire _1343_;
	wire _1344_;
	wire _1345_;
	wire _1346_;
	wire _1347_;
	wire _1348_;
	wire _1349_;
	wire _1350_;
	wire _1351_;
	wire _1352_;
	wire _1353_;
	wire _1354_;
	wire _1355_;
	wire _1356_;
	wire _1357_;
	wire _1358_;
	wire _1359_;
	wire _1360_;
	wire _1361_;
	wire _1362_;
	wire _1363_;
	wire _1364_;
	wire _1365_;
	wire _1366_;
	wire _1367_;
	wire _1368_;
	wire _1369_;
	wire _1370_;
	wire _1371_;
	wire _1372_;
	wire _1373_;
	wire _1374_;
	wire _1375_;
	wire _1376_;
	wire _1377_;
	wire _1378_;
	wire _1379_;
	wire _1380_;
	wire _1381_;
	wire _1382_;
	wire _1383_;
	wire _1384_;
	wire _1385_;
	wire _1386_;
	wire _1387_;
	wire _1388_;
	wire _1389_;
	wire _1390_;
	wire _1391_;
	wire _1392_;
	wire _1393_;
	wire _1394_;
	wire _1395_;
	wire _1396_;
	wire _1397_;
	wire _1398_;
	wire _1399_;
	wire _1400_;
	wire _1401_;
	wire _1402_;
	wire _1403_;
	wire _1404_;
	wire _1405_;
	wire _1406_;
	wire _1407_;
	wire _1408_;
	wire _1409_;
	wire _1410_;
	wire _1411_;
	wire _1412_;
	wire _1413_;
	wire _1414_;
	wire _1415_;
	wire _1416_;
	wire _1417_;
	wire _1418_;
	wire _1419_;
	wire _1420_;
	wire _1421_;
	wire _1422_;
	wire _1423_;
	wire _1424_;
	wire _1425_;
	wire _1426_;
	wire _1427_;
	wire _1428_;
	wire _1429_;
	wire _1430_;
	wire _1431_;
	wire _1432_;
	wire _1433_;
	wire _1434_;
	wire _1435_;
	wire _1436_;
	wire _1437_;
	wire _1438_;
	wire _1439_;
	wire _1440_;
	wire _1441_;
	wire _1442_;
	wire _1443_;
	wire _1444_;
	wire _1445_;
	wire _1446_;
	wire _1447_;
	wire _1448_;
	wire _1449_;
	wire _1450_;
	wire _1451_;
	wire _1452_;
	wire _1453_;
	wire _1454_;
	wire _1455_;
	wire _1456_;
	wire _1457_;
	wire _1458_;
	wire _1459_;
	wire _1460_;
	wire _1461_;
	wire _1462_;
	wire _1463_;
	wire _1464_;
	wire _1465_;
	wire _1466_;
	wire _1467_;
	wire _1468_;
	wire _1469_;
	wire _1470_;
	wire _1471_;
	wire _1472_;
	wire _1473_;
	wire _1474_;
	wire _1475_;
	wire _1476_;
	wire _1477_;
	wire _1478_;
	wire _1479_;
	wire _1480_;
	wire _1481_;
	wire _1482_;
	wire _1483_;
	wire _1484_;
	wire _1485_;
	wire _1486_;
	wire _1487_;
	wire _1488_;
	wire _1489_;
	wire _1490_;
	wire _1491_;
	wire _1492_;
	wire _1493_;
	wire _1494_;
	wire _1495_;
	wire _1496_;
	wire _1497_;
	wire _1498_;
	wire _1499_;
	wire _1500_;
	wire _1501_;
	wire _1502_;
	wire _1503_;
	wire _1504_;
	wire _1505_;
	wire _1506_;
	wire _1507_;
	wire _1508_;
	wire _1509_;
	wire _1510_;
	wire _1511_;
	wire _1512_;
	wire _1513_;
	wire _1514_;
	wire _1515_;
	wire _1516_;
	wire _1517_;
	wire _1518_;
	wire _1519_;
	wire _1520_;
	wire _1521_;
	wire _1522_;
	wire _1523_;
	wire _1524_;
	wire _1525_;
	wire _1526_;
	wire _1527_;
	wire _1528_;
	wire _1529_;
	wire _1530_;
	wire _1531_;
	wire _1532_;
	wire _1533_;
	wire _1534_;
	wire _1535_;
	wire _1536_;
	wire _1537_;
	wire _1538_;
	wire _1539_;
	wire _1540_;
	wire _1541_;
	wire _1542_;
	wire _1543_;
	wire _1544_;
	wire _1545_;
	wire _1546_;
	wire _1547_;
	wire _1548_;
	wire _1549_;
	wire _1550_;
	wire _1551_;
	wire _1552_;
	wire _1553_;
	wire _1554_;
	wire _1555_;
	wire _1556_;
	wire _1557_;
	wire _1558_;
	wire _1559_;
	wire _1560_;
	wire _1561_;
	wire _1562_;
	wire _1563_;
	wire _1564_;
	wire _1565_;
	wire _1566_;
	wire _1567_;
	wire _1568_;
	wire _1569_;
	wire _1570_;
	wire _1571_;
	wire _1572_;
	wire _1573_;
	wire _1574_;
	wire _1575_;
	wire _1576_;
	wire _1577_;
	wire _1578_;
	wire _1579_;
	wire _1580_;
	wire _1581_;
	wire _1582_;
	wire _1583_;
	wire _1584_;
	wire _1585_;
	wire _1586_;
	wire _1587_;
	wire _1588_;
	wire _1589_;
	wire _1590_;
	wire _1591_;
	wire _1592_;
	wire _1593_;
	wire _1594_;
	wire _1595_;
	wire _1596_;
	wire _1597_;
	wire _1598_;
	wire _1599_;
	wire _1600_;
	wire _1601_;
	wire _1602_;
	wire _1603_;
	wire _1604_;
	wire _1605_;
	wire _1606_;
	wire _1607_;
	wire _1608_;
	wire _1609_;
	wire _1610_;
	wire _1611_;
	wire _1612_;
	wire _1613_;
	wire _1614_;
	wire _1615_;
	wire _1616_;
	wire _1617_;
	wire _1618_;
	wire _1619_;
	wire _1620_;
	wire _1621_;
	wire _1622_;
	wire _1623_;
	wire _1624_;
	wire _1625_;
	wire _1626_;
	wire _1627_;
	wire _1628_;
	wire _1629_;
	wire _1630_;
	wire _1631_;
	wire _1632_;
	wire _1633_;
	wire _1634_;
	wire _1635_;
	wire _1636_;
	wire _1637_;
	wire _1638_;
	wire _1639_;
	wire _1640_;
	wire _1641_;
	wire _1642_;
	wire _1643_;
	wire _1644_;
	wire _1645_;
	wire _1646_;
	wire _1647_;
	wire _1648_;
	wire _1649_;
	wire _1650_;
	wire _1651_;
	wire _1652_;
	wire _1653_;
	wire _1654_;
	wire _1655_;
	wire _1656_;
	wire _1657_;
	wire _1658_;
	wire _1659_;
	wire _1660_;
	wire _1661_;
	wire _1662_;
	wire _1663_;
	wire _1664_;
	wire _1665_;
	wire _1666_;
	wire _1667_;
	wire _1668_;
	wire _1669_;
	wire _1670_;
	wire _1671_;
	wire _1672_;
	wire _1673_;
	wire _1674_;
	wire _1675_;
	wire _1676_;
	wire _1677_;
	wire _1678_;
	wire _1679_;
	wire _1680_;
	wire _1681_;
	wire _1682_;
	wire _1683_;
	wire _1684_;
	wire _1685_;
	wire _1686_;
	wire _1687_;
	wire _1688_;
	wire _1689_;
	wire _1690_;
	wire _1691_;
	wire _1692_;
	wire _1693_;
	wire _1694_;
	wire _1695_;
	wire _1696_;
	wire _1697_;
	wire _1698_;
	wire _1699_;
	wire _1700_;
	wire _1701_;
	wire _1702_;
	wire _1703_;
	wire _1704_;
	wire _1705_;
	wire _1706_;
	wire _1707_;
	wire _1708_;
	wire _1709_;
	wire _1710_;
	wire _1711_;
	wire _1712_;
	wire _1713_;
	wire _1714_;
	wire _1715_;
	wire _1716_;
	wire _1717_;
	wire _1718_;
	wire _1719_;
	wire _1720_;
	wire _1721_;
	wire _1722_;
	wire _1723_;
	wire _1724_;
	wire _1725_;
	wire _1726_;
	wire _1727_;
	wire _1728_;
	wire _1729_;
	wire _1730_;
	wire _1731_;
	wire _1732_;
	wire _1733_;
	wire _1734_;
	wire _1735_;
	wire _1736_;
	wire _1737_;
	wire _1738_;
	wire _1739_;
	wire _1740_;
	wire _1741_;
	wire _1742_;
	wire _1743_;
	wire _1744_;
	wire _1745_;
	wire _1746_;
	wire _1747_;
	wire _1748_;
	wire _1749_;
	wire _1750_;
	wire _1751_;
	wire _1752_;
	wire _1753_;
	wire _1754_;
	wire _1755_;
	wire _1756_;
	wire _1757_;
	wire _1758_;
	wire _1759_;
	wire _1760_;
	wire _1761_;
	wire _1762_;
	wire _1763_;
	wire _1764_;
	wire _1765_;
	wire [1:0] _1766_;
	wire [1:0] _1767_;
	wire [1:0] _1768_;
	wire [1:0] _1769_;
	wire [1:0] _1770_;
	wire [1:0] _1771_;
	wire [1:0] _1772_;
	wire [1:0] _1773_;
	wire [2:0] _1774_;
	wire [1:0] _1775_;
	wire [3:0] _1776_;
	input wire [13:0] io_in;
	output wire [13:0] io_out;
	reg [2:0] \mchip.DUT.a ;
	wire [2:0] \mchip.DUT.b ;
	reg [2:0] \mchip.DUT.c ;
	reg [14:0] \mchip.DUT.character ;
	wire \mchip.DUT.clk ;
	reg [1:0] \mchip.DUT.count ;
	wire [23:0] \mchip.DUT.data_in ;
	reg [8:0] \mchip.DUT.encoded_mask ;
	reg [8:0] \mchip.DUT.encoded_value ;
	wire [2:0] \mchip.DUT.encoded_value_h[0] ;
	wire [2:0] \mchip.DUT.encoded_value_h[1] ;
	reg [2:0] \mchip.DUT.encoded_value_h[2] ;
	reg [2:0] \mchip.DUT.encoded_value_h[3] ;
	reg [2:0] \mchip.DUT.encoded_value_h[4] ;
	reg [2:0] \mchip.DUT.encoded_value_h[5] ;
	wire [23:0] \mchip.DUT.freq_calc_ins.data_in ;
	wire [8:0] \mchip.DUT.freq_calc_ins.freq_in ;
	wire [56:0] \mchip.DUT.freq_calc_ins.node ;
	wire [31:0] \mchip.DUT.freq_calc_ins.sv2v_autoblock_1.i ;
	reg [8:0] \mchip.DUT.freq_in ;
	wire [19:0] \mchip.DUT.huff_tree[0] ;
	wire [19:0] \mchip.DUT.huff_tree[1] ;
	reg [19:0] \mchip.DUT.huff_tree[2] ;
	reg [19:0] \mchip.DUT.huff_tree[3] ;
	reg [19:0] \mchip.DUT.huff_tree[4] ;
	reg [19:0] \mchip.DUT.huff_tree[5] ;
	wire [56:0] \mchip.DUT.in_huff_tree ;
	wire [56:0] \mchip.DUT.initial_node ;
	wire [11:0] \mchip.DUT.io_in ;
	wire [11:0] \mchip.DUT.io_out ;
	wire [18:0] \mchip.DUT.merge_nodes_ins.merged_node ;
	wire [18:0] \mchip.DUT.merge_nodes_ins.min_node ;
	wire [18:0] \mchip.DUT.merge_nodes_ins.second_min_node ;
	wire [18:0] \mchip.DUT.merged_node ;
	wire \mchip.DUT.node_sorter_ins.clk ;
	wire [56:0] \mchip.DUT.node_sorter_ins.input_node ;
	reg [56:0] \mchip.DUT.node_sorter_ins.output_node ;
	wire [75:0] \mchip.DUT.out_huff_tree ;
	wire \mchip.DUT.reset ;
	reg [6:0] \mchip.DUT.state ;
	wire \mchip.clock ;
	wire [11:0] \mchip.io_in ;
	wire [11:0] \mchip.io_out ;
	wire \mchip.reset ;
	assign _1278_ = ~\mchip.DUT.huff_tree[1] [14];
	assign _1279_ = \mchip.DUT.huff_tree[1] [13] ^ \mchip.DUT.huff_tree[4] [19];
	assign _1280_ = \mchip.DUT.huff_tree[1] [12] ^ \mchip.DUT.huff_tree[4] [18];
	assign _1281_ = \mchip.DUT.huff_tree[1] [11] ^ \mchip.DUT.huff_tree[4] [17];
	assign _1282_ = _1281_ | _1280_;
	assign _1283_ = \mchip.DUT.huff_tree[1] [10] ^ \mchip.DUT.huff_tree[4] [16];
	assign _1284_ = \mchip.DUT.huff_tree[1] [9] ^ \mchip.DUT.huff_tree[4] [15];
	assign _1285_ = _1284_ | _1283_;
	assign _1286_ = _1285_ | _1282_;
	assign _1287_ = _1286_ | _1279_;
	assign _1288_ = ~(\mchip.DUT.huff_tree[1] [4] ^ \mchip.DUT.huff_tree[4] [15]);
	assign _1289_ = \mchip.DUT.huff_tree[1] [5] ^ \mchip.DUT.huff_tree[4] [16];
	assign _1290_ = _1288_ & ~_1289_;
	assign _1291_ = \mchip.DUT.huff_tree[1] [7] ^ \mchip.DUT.huff_tree[4] [18];
	assign _1292_ = \mchip.DUT.huff_tree[1] [6] ^ \mchip.DUT.huff_tree[4] [17];
	assign _1293_ = _1292_ | _1291_;
	assign _1294_ = _1290_ & ~_1293_;
	assign _1295_ = \mchip.DUT.huff_tree[1] [8] ^ \mchip.DUT.huff_tree[4] [19];
	assign _1296_ = _1294_ & ~_1295_;
	assign _1297_ = _1287_ & ~_1296_;
	assign _1298_ = _1278_ & ~_1297_;
	assign _1299_ = _1298_ | \mchip.DUT.huff_tree[4] [2];
	assign _1300_ = ~\mchip.DUT.huff_tree[2] [14];
	assign _1301_ = \mchip.DUT.huff_tree[2] [13] ^ \mchip.DUT.huff_tree[4] [19];
	assign _1302_ = \mchip.DUT.huff_tree[2] [12] ^ \mchip.DUT.huff_tree[4] [18];
	assign _1303_ = \mchip.DUT.huff_tree[2] [11] ^ \mchip.DUT.huff_tree[4] [17];
	assign _1304_ = _1303_ | _1302_;
	assign _1305_ = \mchip.DUT.huff_tree[2] [10] ^ \mchip.DUT.huff_tree[4] [16];
	assign _1306_ = \mchip.DUT.huff_tree[2] [9] ^ \mchip.DUT.huff_tree[4] [15];
	assign _1307_ = _1306_ | _1305_;
	assign _1308_ = _1307_ | _1304_;
	assign _1309_ = _1308_ | _1301_;
	assign _1310_ = ~(\mchip.DUT.huff_tree[2] [4] ^ \mchip.DUT.huff_tree[4] [15]);
	assign _1311_ = \mchip.DUT.huff_tree[2] [5] ^ \mchip.DUT.huff_tree[4] [16];
	assign _1312_ = _1310_ & ~_1311_;
	assign _1313_ = \mchip.DUT.huff_tree[2] [7] ^ \mchip.DUT.huff_tree[4] [18];
	assign _1314_ = \mchip.DUT.huff_tree[2] [6] ^ \mchip.DUT.huff_tree[4] [17];
	assign _1315_ = _1314_ | _1313_;
	assign _1316_ = _1312_ & ~_1315_;
	assign _1317_ = \mchip.DUT.huff_tree[2] [8] ^ \mchip.DUT.huff_tree[4] [19];
	assign _1318_ = _1316_ & ~_1317_;
	assign _1319_ = _1309_ & ~_1318_;
	assign _1320_ = _1300_ & ~_1319_;
	assign _1321_ = _1299_ & ~_1320_;
	assign _1322_ = ~\mchip.DUT.huff_tree[3] [14];
	assign _1323_ = \mchip.DUT.huff_tree[3] [13] ^ \mchip.DUT.huff_tree[4] [19];
	assign _1324_ = \mchip.DUT.huff_tree[3] [12] ^ \mchip.DUT.huff_tree[4] [18];
	assign _1325_ = \mchip.DUT.huff_tree[3] [11] ^ \mchip.DUT.huff_tree[4] [17];
	assign _1326_ = _1325_ | _1324_;
	assign _1327_ = \mchip.DUT.huff_tree[3] [10] ^ \mchip.DUT.huff_tree[4] [16];
	assign _1328_ = \mchip.DUT.huff_tree[3] [9] ^ \mchip.DUT.huff_tree[4] [15];
	assign _1329_ = _1328_ | _1327_;
	assign _1330_ = _1329_ | _1326_;
	assign _1331_ = _1330_ | _1323_;
	assign _1332_ = ~(\mchip.DUT.huff_tree[3] [4] ^ \mchip.DUT.huff_tree[4] [15]);
	assign _1333_ = \mchip.DUT.huff_tree[3] [5] ^ \mchip.DUT.huff_tree[4] [16];
	assign _1334_ = _1332_ & ~_1333_;
	assign _1335_ = \mchip.DUT.huff_tree[3] [7] ^ \mchip.DUT.huff_tree[4] [18];
	assign _1336_ = \mchip.DUT.huff_tree[3] [6] ^ \mchip.DUT.huff_tree[4] [17];
	assign _1337_ = _1336_ | _1335_;
	assign _1338_ = _1334_ & ~_1337_;
	assign _1339_ = \mchip.DUT.huff_tree[3] [8] ^ \mchip.DUT.huff_tree[4] [19];
	assign _1340_ = _1338_ & ~_1339_;
	assign _1341_ = _1331_ & ~_1340_;
	assign _1342_ = _1322_ & ~_1341_;
	assign _1343_ = _1342_ | _1321_;
	assign _1344_ = ~\mchip.DUT.huff_tree[4] [14];
	assign _1345_ = \mchip.DUT.huff_tree[4] [13] ^ \mchip.DUT.huff_tree[4] [19];
	assign _1346_ = \mchip.DUT.huff_tree[4] [12] ^ \mchip.DUT.huff_tree[4] [18];
	assign _1347_ = \mchip.DUT.huff_tree[4] [11] ^ \mchip.DUT.huff_tree[4] [17];
	assign _1348_ = _1347_ | _1346_;
	assign _1349_ = \mchip.DUT.huff_tree[4] [10] ^ \mchip.DUT.huff_tree[4] [16];
	assign _1350_ = \mchip.DUT.huff_tree[4] [9] ^ \mchip.DUT.huff_tree[4] [15];
	assign _1351_ = _1350_ | _1349_;
	assign _1352_ = _1351_ | _1348_;
	assign _1353_ = _1352_ | _1345_;
	assign _1354_ = ~(\mchip.DUT.huff_tree[4] [4] ^ \mchip.DUT.huff_tree[4] [15]);
	assign _1355_ = \mchip.DUT.huff_tree[4] [5] ^ \mchip.DUT.huff_tree[4] [16];
	assign _1356_ = _1354_ & ~_1355_;
	assign _1357_ = \mchip.DUT.huff_tree[4] [7] ^ \mchip.DUT.huff_tree[4] [18];
	assign _1358_ = \mchip.DUT.huff_tree[4] [6] ^ \mchip.DUT.huff_tree[4] [17];
	assign _1359_ = _1358_ | _1357_;
	assign _1360_ = _1356_ & ~_1359_;
	assign _1361_ = \mchip.DUT.huff_tree[4] [8] ^ \mchip.DUT.huff_tree[4] [19];
	assign _1362_ = _1360_ & ~_1361_;
	assign _1363_ = _1353_ & ~_1362_;
	assign _1364_ = _1344_ & ~_1363_;
	assign _1365_ = _1343_ & ~_1364_;
	assign _1366_ = ~\mchip.DUT.huff_tree[5] [14];
	assign _1367_ = \mchip.DUT.huff_tree[4] [19] ^ \mchip.DUT.huff_tree[5] [13];
	assign _1368_ = \mchip.DUT.huff_tree[4] [18] ^ \mchip.DUT.huff_tree[5] [12];
	assign _1369_ = \mchip.DUT.huff_tree[4] [17] ^ \mchip.DUT.huff_tree[5] [11];
	assign _1370_ = _1369_ | _1368_;
	assign _1371_ = \mchip.DUT.huff_tree[4] [16] ^ \mchip.DUT.huff_tree[5] [10];
	assign _1372_ = \mchip.DUT.huff_tree[4] [15] ^ \mchip.DUT.huff_tree[5] [9];
	assign _1373_ = _1372_ | _1371_;
	assign _1374_ = _1373_ | _1370_;
	assign _1375_ = _1374_ | _1367_;
	assign _1376_ = ~(\mchip.DUT.huff_tree[5] [4] ^ \mchip.DUT.huff_tree[4] [15]);
	assign _1377_ = \mchip.DUT.huff_tree[5] [5] ^ \mchip.DUT.huff_tree[4] [16];
	assign _1378_ = _1376_ & ~_1377_;
	assign _1379_ = \mchip.DUT.huff_tree[5] [7] ^ \mchip.DUT.huff_tree[4] [18];
	assign _1380_ = \mchip.DUT.huff_tree[5] [6] ^ \mchip.DUT.huff_tree[4] [17];
	assign _1381_ = _1380_ | _1379_;
	assign _1382_ = _1378_ & ~_1381_;
	assign _1383_ = \mchip.DUT.huff_tree[5] [8] ^ \mchip.DUT.huff_tree[4] [19];
	assign _1384_ = _1382_ & ~_1383_;
	assign _1385_ = _1375_ & ~_1384_;
	assign _1386_ = _1366_ & ~_1385_;
	assign _0017_ = _1386_ | _1365_;
	assign _1387_ = \mchip.DUT.huff_tree[4] [3] & ~_1298_;
	assign _1388_ = _1387_ | _1320_;
	assign _1389_ = ~(_1388_ | _1342_);
	assign _1390_ = _1389_ | _1364_;
	assign _0040_ = ~(_1390_ | _1386_);
	assign _1391_ = \mchip.DUT.huff_tree[3] [19] ^ \mchip.DUT.huff_tree[1] [13];
	assign _1392_ = \mchip.DUT.huff_tree[3] [18] ^ \mchip.DUT.huff_tree[1] [12];
	assign _1393_ = \mchip.DUT.huff_tree[3] [17] ^ \mchip.DUT.huff_tree[1] [11];
	assign _1394_ = _1393_ | _1392_;
	assign _1395_ = \mchip.DUT.huff_tree[3] [16] ^ \mchip.DUT.huff_tree[1] [10];
	assign _1396_ = \mchip.DUT.huff_tree[3] [15] ^ \mchip.DUT.huff_tree[1] [9];
	assign _1397_ = _1396_ | _1395_;
	assign _1398_ = _1397_ | _1394_;
	assign _1399_ = _1398_ | _1391_;
	assign _1400_ = ~(\mchip.DUT.huff_tree[3] [15] ^ \mchip.DUT.huff_tree[1] [4]);
	assign _1401_ = \mchip.DUT.huff_tree[3] [16] ^ \mchip.DUT.huff_tree[1] [5];
	assign _1402_ = _1400_ & ~_1401_;
	assign _1403_ = \mchip.DUT.huff_tree[3] [18] ^ \mchip.DUT.huff_tree[1] [7];
	assign _1404_ = \mchip.DUT.huff_tree[3] [17] ^ \mchip.DUT.huff_tree[1] [6];
	assign _1405_ = _1404_ | _1403_;
	assign _1406_ = _1402_ & ~_1405_;
	assign _1407_ = \mchip.DUT.huff_tree[3] [19] ^ \mchip.DUT.huff_tree[1] [8];
	assign _1408_ = _1406_ & ~_1407_;
	assign _1409_ = _1399_ & ~_1408_;
	assign _1410_ = _1278_ & ~_1409_;
	assign _1411_ = _1410_ | \mchip.DUT.huff_tree[3] [2];
	assign _1412_ = \mchip.DUT.huff_tree[3] [19] ^ \mchip.DUT.huff_tree[2] [13];
	assign _1413_ = \mchip.DUT.huff_tree[3] [18] ^ \mchip.DUT.huff_tree[2] [12];
	assign _1414_ = \mchip.DUT.huff_tree[3] [17] ^ \mchip.DUT.huff_tree[2] [11];
	assign _1415_ = _1414_ | _1413_;
	assign _1416_ = \mchip.DUT.huff_tree[3] [16] ^ \mchip.DUT.huff_tree[2] [10];
	assign _1417_ = \mchip.DUT.huff_tree[3] [15] ^ \mchip.DUT.huff_tree[2] [9];
	assign _1418_ = _1417_ | _1416_;
	assign _1419_ = _1418_ | _1415_;
	assign _1420_ = _1419_ | _1412_;
	assign _1421_ = ~(\mchip.DUT.huff_tree[3] [15] ^ \mchip.DUT.huff_tree[2] [4]);
	assign _1422_ = \mchip.DUT.huff_tree[3] [16] ^ \mchip.DUT.huff_tree[2] [5];
	assign _1423_ = _1421_ & ~_1422_;
	assign _1424_ = \mchip.DUT.huff_tree[3] [18] ^ \mchip.DUT.huff_tree[2] [7];
	assign _1425_ = \mchip.DUT.huff_tree[3] [17] ^ \mchip.DUT.huff_tree[2] [6];
	assign _1426_ = _1425_ | _1424_;
	assign _1427_ = _1423_ & ~_1426_;
	assign _1428_ = \mchip.DUT.huff_tree[3] [19] ^ \mchip.DUT.huff_tree[2] [8];
	assign _1429_ = _1427_ & ~_1428_;
	assign _1430_ = _1420_ & ~_1429_;
	assign _1431_ = _1300_ & ~_1430_;
	assign _1432_ = _1411_ & ~_1431_;
	assign _1433_ = \mchip.DUT.huff_tree[3] [19] ^ \mchip.DUT.huff_tree[3] [13];
	assign _1434_ = \mchip.DUT.huff_tree[3] [18] ^ \mchip.DUT.huff_tree[3] [12];
	assign _1435_ = \mchip.DUT.huff_tree[3] [17] ^ \mchip.DUT.huff_tree[3] [11];
	assign _1436_ = _1435_ | _1434_;
	assign _1437_ = \mchip.DUT.huff_tree[3] [16] ^ \mchip.DUT.huff_tree[3] [10];
	assign _1438_ = \mchip.DUT.huff_tree[3] [15] ^ \mchip.DUT.huff_tree[3] [9];
	assign _1439_ = _1438_ | _1437_;
	assign _1440_ = _1439_ | _1436_;
	assign _1441_ = _1440_ | _1433_;
	assign _1442_ = ~(\mchip.DUT.huff_tree[3] [15] ^ \mchip.DUT.huff_tree[3] [4]);
	assign _1443_ = \mchip.DUT.huff_tree[3] [16] ^ \mchip.DUT.huff_tree[3] [5];
	assign _1444_ = _1442_ & ~_1443_;
	assign _1445_ = \mchip.DUT.huff_tree[3] [18] ^ \mchip.DUT.huff_tree[3] [7];
	assign _1446_ = \mchip.DUT.huff_tree[3] [17] ^ \mchip.DUT.huff_tree[3] [6];
	assign _1447_ = _1446_ | _1445_;
	assign _1448_ = _1444_ & ~_1447_;
	assign _1449_ = \mchip.DUT.huff_tree[3] [19] ^ \mchip.DUT.huff_tree[3] [8];
	assign _1450_ = _1448_ & ~_1449_;
	assign _1451_ = _1441_ & ~_1450_;
	assign _1452_ = _1322_ & ~_1451_;
	assign _1453_ = _1452_ | _1432_;
	assign _1454_ = \mchip.DUT.huff_tree[3] [19] ^ \mchip.DUT.huff_tree[4] [13];
	assign _1455_ = \mchip.DUT.huff_tree[3] [18] ^ \mchip.DUT.huff_tree[4] [12];
	assign _1456_ = \mchip.DUT.huff_tree[3] [17] ^ \mchip.DUT.huff_tree[4] [11];
	assign _1457_ = _1456_ | _1455_;
	assign _1458_ = \mchip.DUT.huff_tree[3] [16] ^ \mchip.DUT.huff_tree[4] [10];
	assign _1459_ = \mchip.DUT.huff_tree[3] [15] ^ \mchip.DUT.huff_tree[4] [9];
	assign _1460_ = _1459_ | _1458_;
	assign _1461_ = _1460_ | _1457_;
	assign _1462_ = _1461_ | _1454_;
	assign _1463_ = ~(\mchip.DUT.huff_tree[3] [15] ^ \mchip.DUT.huff_tree[4] [4]);
	assign _1464_ = \mchip.DUT.huff_tree[3] [16] ^ \mchip.DUT.huff_tree[4] [5];
	assign _1465_ = _1463_ & ~_1464_;
	assign _1466_ = \mchip.DUT.huff_tree[3] [18] ^ \mchip.DUT.huff_tree[4] [7];
	assign _1467_ = \mchip.DUT.huff_tree[3] [17] ^ \mchip.DUT.huff_tree[4] [6];
	assign _1468_ = _1467_ | _1466_;
	assign _1469_ = _1465_ & ~_1468_;
	assign _1470_ = \mchip.DUT.huff_tree[3] [19] ^ \mchip.DUT.huff_tree[4] [8];
	assign _1471_ = _1469_ & ~_1470_;
	assign _1472_ = _1462_ & ~_1471_;
	assign _1473_ = _1344_ & ~_1472_;
	assign _1474_ = _1453_ & ~_1473_;
	assign _1475_ = \mchip.DUT.huff_tree[3] [19] ^ \mchip.DUT.huff_tree[5] [13];
	assign _1476_ = \mchip.DUT.huff_tree[3] [18] ^ \mchip.DUT.huff_tree[5] [12];
	assign _1477_ = \mchip.DUT.huff_tree[3] [17] ^ \mchip.DUT.huff_tree[5] [11];
	assign _1478_ = _1477_ | _1476_;
	assign _1479_ = \mchip.DUT.huff_tree[3] [16] ^ \mchip.DUT.huff_tree[5] [10];
	assign _1480_ = \mchip.DUT.huff_tree[3] [15] ^ \mchip.DUT.huff_tree[5] [9];
	assign _1481_ = _1480_ | _1479_;
	assign _1482_ = _1481_ | _1478_;
	assign _1483_ = _1482_ | _1475_;
	assign _1484_ = ~(\mchip.DUT.huff_tree[3] [15] ^ \mchip.DUT.huff_tree[5] [4]);
	assign _1485_ = \mchip.DUT.huff_tree[3] [16] ^ \mchip.DUT.huff_tree[5] [5];
	assign _1486_ = _1484_ & ~_1485_;
	assign _1487_ = \mchip.DUT.huff_tree[3] [18] ^ \mchip.DUT.huff_tree[5] [7];
	assign _1488_ = \mchip.DUT.huff_tree[3] [17] ^ \mchip.DUT.huff_tree[5] [6];
	assign _1489_ = _1488_ | _1487_;
	assign _1490_ = _1486_ & ~_1489_;
	assign _1491_ = \mchip.DUT.huff_tree[3] [19] ^ \mchip.DUT.huff_tree[5] [8];
	assign _1492_ = _1490_ & ~_1491_;
	assign _1493_ = _1483_ & ~_1492_;
	assign _1494_ = _1366_ & ~_1493_;
	assign _0018_ = _1494_ | _1474_;
	assign _1495_ = \mchip.DUT.huff_tree[3] [3] & ~_1410_;
	assign _1496_ = _1495_ | _1431_;
	assign _1497_ = ~(_1496_ | _1452_);
	assign _1498_ = _1497_ | _1473_;
	assign _0039_ = ~(_1498_ | _1494_);
	assign _1499_ = \mchip.DUT.huff_tree[2] [19] ^ \mchip.DUT.huff_tree[1] [13];
	assign _1500_ = \mchip.DUT.huff_tree[2] [18] ^ \mchip.DUT.huff_tree[1] [12];
	assign _1501_ = \mchip.DUT.huff_tree[2] [17] ^ \mchip.DUT.huff_tree[1] [11];
	assign _1502_ = _1501_ | _1500_;
	assign _1503_ = \mchip.DUT.huff_tree[2] [16] ^ \mchip.DUT.huff_tree[1] [10];
	assign _1504_ = \mchip.DUT.huff_tree[2] [15] ^ \mchip.DUT.huff_tree[1] [9];
	assign _1505_ = _1504_ | _1503_;
	assign _1506_ = _1505_ | _1502_;
	assign _1507_ = _1506_ | _1499_;
	assign _1508_ = ~(\mchip.DUT.huff_tree[2] [15] ^ \mchip.DUT.huff_tree[1] [4]);
	assign _1509_ = \mchip.DUT.huff_tree[2] [16] ^ \mchip.DUT.huff_tree[1] [5];
	assign _1510_ = _1508_ & ~_1509_;
	assign _1511_ = \mchip.DUT.huff_tree[2] [18] ^ \mchip.DUT.huff_tree[1] [7];
	assign _1512_ = \mchip.DUT.huff_tree[2] [17] ^ \mchip.DUT.huff_tree[1] [6];
	assign _1513_ = _1512_ | _1511_;
	assign _1514_ = _1510_ & ~_1513_;
	assign _1515_ = \mchip.DUT.huff_tree[2] [19] ^ \mchip.DUT.huff_tree[1] [8];
	assign _1516_ = _1514_ & ~_1515_;
	assign _1517_ = _1507_ & ~_1516_;
	assign _1518_ = _1278_ & ~_1517_;
	assign _1519_ = _1518_ | \mchip.DUT.huff_tree[2] [2];
	assign _1520_ = \mchip.DUT.huff_tree[2] [19] ^ \mchip.DUT.huff_tree[2] [13];
	assign _1521_ = \mchip.DUT.huff_tree[2] [18] ^ \mchip.DUT.huff_tree[2] [12];
	assign _1522_ = \mchip.DUT.huff_tree[2] [17] ^ \mchip.DUT.huff_tree[2] [11];
	assign _1523_ = _1522_ | _1521_;
	assign _1524_ = \mchip.DUT.huff_tree[2] [16] ^ \mchip.DUT.huff_tree[2] [10];
	assign _1525_ = \mchip.DUT.huff_tree[2] [15] ^ \mchip.DUT.huff_tree[2] [9];
	assign _1526_ = _1525_ | _1524_;
	assign _1527_ = _1526_ | _1523_;
	assign _1528_ = _1527_ | _1520_;
	assign _1529_ = ~(\mchip.DUT.huff_tree[2] [15] ^ \mchip.DUT.huff_tree[2] [4]);
	assign _1530_ = \mchip.DUT.huff_tree[2] [16] ^ \mchip.DUT.huff_tree[2] [5];
	assign _1531_ = _1529_ & ~_1530_;
	assign _1532_ = \mchip.DUT.huff_tree[2] [18] ^ \mchip.DUT.huff_tree[2] [7];
	assign _1533_ = \mchip.DUT.huff_tree[2] [17] ^ \mchip.DUT.huff_tree[2] [6];
	assign _1534_ = _1533_ | _1532_;
	assign _1535_ = _1531_ & ~_1534_;
	assign _1536_ = \mchip.DUT.huff_tree[2] [19] ^ \mchip.DUT.huff_tree[2] [8];
	assign _1537_ = _1535_ & ~_1536_;
	assign _1538_ = _1528_ & ~_1537_;
	assign _1539_ = _1300_ & ~_1538_;
	assign _1540_ = _1519_ & ~_1539_;
	assign _1541_ = \mchip.DUT.huff_tree[2] [19] ^ \mchip.DUT.huff_tree[3] [13];
	assign _1542_ = \mchip.DUT.huff_tree[2] [18] ^ \mchip.DUT.huff_tree[3] [12];
	assign _1543_ = \mchip.DUT.huff_tree[2] [17] ^ \mchip.DUT.huff_tree[3] [11];
	assign _1544_ = _1543_ | _1542_;
	assign _1545_ = \mchip.DUT.huff_tree[2] [16] ^ \mchip.DUT.huff_tree[3] [10];
	assign _1546_ = \mchip.DUT.huff_tree[2] [15] ^ \mchip.DUT.huff_tree[3] [9];
	assign _1547_ = _1546_ | _1545_;
	assign _1548_ = _1547_ | _1544_;
	assign _1549_ = _1548_ | _1541_;
	assign _1550_ = ~(\mchip.DUT.huff_tree[2] [15] ^ \mchip.DUT.huff_tree[3] [4]);
	assign _1551_ = \mchip.DUT.huff_tree[2] [16] ^ \mchip.DUT.huff_tree[3] [5];
	assign _1552_ = _1550_ & ~_1551_;
	assign _1553_ = \mchip.DUT.huff_tree[2] [18] ^ \mchip.DUT.huff_tree[3] [7];
	assign _1554_ = \mchip.DUT.huff_tree[2] [17] ^ \mchip.DUT.huff_tree[3] [6];
	assign _1555_ = _1554_ | _1553_;
	assign _1556_ = _1552_ & ~_1555_;
	assign _1557_ = \mchip.DUT.huff_tree[2] [19] ^ \mchip.DUT.huff_tree[3] [8];
	assign _1558_ = _1556_ & ~_1557_;
	assign _1559_ = _1549_ & ~_1558_;
	assign _1560_ = _1322_ & ~_1559_;
	assign _1561_ = _1560_ | _1540_;
	assign _1562_ = \mchip.DUT.huff_tree[2] [19] ^ \mchip.DUT.huff_tree[4] [13];
	assign _1563_ = \mchip.DUT.huff_tree[2] [18] ^ \mchip.DUT.huff_tree[4] [12];
	assign _1564_ = \mchip.DUT.huff_tree[2] [17] ^ \mchip.DUT.huff_tree[4] [11];
	assign _1565_ = _1564_ | _1563_;
	assign _1566_ = \mchip.DUT.huff_tree[2] [16] ^ \mchip.DUT.huff_tree[4] [10];
	assign _1567_ = \mchip.DUT.huff_tree[2] [15] ^ \mchip.DUT.huff_tree[4] [9];
	assign _1568_ = _1567_ | _1566_;
	assign _1569_ = _1568_ | _1565_;
	assign _1570_ = _1569_ | _1562_;
	assign _1571_ = ~(\mchip.DUT.huff_tree[2] [15] ^ \mchip.DUT.huff_tree[4] [4]);
	assign _1572_ = \mchip.DUT.huff_tree[2] [16] ^ \mchip.DUT.huff_tree[4] [5];
	assign _1573_ = _1571_ & ~_1572_;
	assign _1574_ = \mchip.DUT.huff_tree[2] [18] ^ \mchip.DUT.huff_tree[4] [7];
	assign _1575_ = \mchip.DUT.huff_tree[2] [17] ^ \mchip.DUT.huff_tree[4] [6];
	assign _1576_ = _1575_ | _1574_;
	assign _1577_ = _1573_ & ~_1576_;
	assign _1578_ = \mchip.DUT.huff_tree[2] [19] ^ \mchip.DUT.huff_tree[4] [8];
	assign _1579_ = _1577_ & ~_1578_;
	assign _1580_ = _1570_ & ~_1579_;
	assign _1581_ = _1344_ & ~_1580_;
	assign _1582_ = _1561_ & ~_1581_;
	assign _1583_ = \mchip.DUT.huff_tree[2] [19] ^ \mchip.DUT.huff_tree[5] [13];
	assign _1584_ = \mchip.DUT.huff_tree[2] [18] ^ \mchip.DUT.huff_tree[5] [12];
	assign _1585_ = \mchip.DUT.huff_tree[2] [17] ^ \mchip.DUT.huff_tree[5] [11];
	assign _1586_ = _1585_ | _1584_;
	assign _1587_ = \mchip.DUT.huff_tree[2] [16] ^ \mchip.DUT.huff_tree[5] [10];
	assign _1588_ = \mchip.DUT.huff_tree[2] [15] ^ \mchip.DUT.huff_tree[5] [9];
	assign _1589_ = _1588_ | _1587_;
	assign _1590_ = _1589_ | _1586_;
	assign _1591_ = _1590_ | _1583_;
	assign _1592_ = ~(\mchip.DUT.huff_tree[2] [15] ^ \mchip.DUT.huff_tree[5] [4]);
	assign _1593_ = \mchip.DUT.huff_tree[2] [16] ^ \mchip.DUT.huff_tree[5] [5];
	assign _1594_ = _1592_ & ~_1593_;
	assign _1595_ = \mchip.DUT.huff_tree[2] [18] ^ \mchip.DUT.huff_tree[5] [7];
	assign _1596_ = \mchip.DUT.huff_tree[2] [17] ^ \mchip.DUT.huff_tree[5] [6];
	assign _1597_ = _1596_ | _1595_;
	assign _1598_ = _1594_ & ~_1597_;
	assign _1599_ = \mchip.DUT.huff_tree[2] [19] ^ \mchip.DUT.huff_tree[5] [8];
	assign _1600_ = _1598_ & ~_1599_;
	assign _1601_ = _1591_ & ~_1600_;
	assign _1602_ = _1366_ & ~_1601_;
	assign _0019_ = _1602_ | _1582_;
	assign _1603_ = \mchip.DUT.huff_tree[2] [3] & ~_1518_;
	assign _1604_ = _1603_ | _1539_;
	assign _1605_ = ~(_1604_ | _1560_);
	assign _1606_ = _1605_ | _1581_;
	assign _0038_ = ~(_1606_ | _1602_);
	assign _1775_[0] = ~\mchip.DUT.count [0];
	assign _1775_[1] = ~(\mchip.DUT.count [1] ^ \mchip.DUT.count [0]);
	assign _1607_ = \mchip.DUT.huff_tree[5] [19] ^ \mchip.DUT.huff_tree[1] [13];
	assign _1608_ = \mchip.DUT.huff_tree[5] [18] ^ \mchip.DUT.huff_tree[1] [12];
	assign _1609_ = \mchip.DUT.huff_tree[5] [17] ^ \mchip.DUT.huff_tree[1] [11];
	assign _1610_ = _1609_ | _1608_;
	assign _1611_ = \mchip.DUT.huff_tree[5] [16] ^ \mchip.DUT.huff_tree[1] [10];
	assign _1612_ = \mchip.DUT.huff_tree[5] [15] ^ \mchip.DUT.huff_tree[1] [9];
	assign _1613_ = _1612_ | _1611_;
	assign _1614_ = _1613_ | _1610_;
	assign _1615_ = _1614_ | _1607_;
	assign _1616_ = ~(\mchip.DUT.huff_tree[5] [15] ^ \mchip.DUT.huff_tree[1] [4]);
	assign _1617_ = \mchip.DUT.huff_tree[5] [16] ^ \mchip.DUT.huff_tree[1] [5];
	assign _1618_ = _1616_ & ~_1617_;
	assign _1619_ = \mchip.DUT.huff_tree[5] [18] ^ \mchip.DUT.huff_tree[1] [7];
	assign _1620_ = \mchip.DUT.huff_tree[5] [17] ^ \mchip.DUT.huff_tree[1] [6];
	assign _1621_ = _1620_ | _1619_;
	assign _1622_ = _1618_ & ~_1621_;
	assign _1623_ = \mchip.DUT.huff_tree[5] [19] ^ \mchip.DUT.huff_tree[1] [8];
	assign _1624_ = _1622_ & ~_1623_;
	assign _1625_ = _1615_ & ~_1624_;
	assign _1626_ = _1278_ & ~_1625_;
	assign _1627_ = _1626_ | \mchip.DUT.huff_tree[5] [2];
	assign _1628_ = \mchip.DUT.huff_tree[5] [19] ^ \mchip.DUT.huff_tree[2] [13];
	assign _1629_ = \mchip.DUT.huff_tree[5] [18] ^ \mchip.DUT.huff_tree[2] [12];
	assign _1630_ = \mchip.DUT.huff_tree[5] [17] ^ \mchip.DUT.huff_tree[2] [11];
	assign _1631_ = _1630_ | _1629_;
	assign _1632_ = \mchip.DUT.huff_tree[5] [16] ^ \mchip.DUT.huff_tree[2] [10];
	assign _1633_ = \mchip.DUT.huff_tree[5] [15] ^ \mchip.DUT.huff_tree[2] [9];
	assign _1634_ = _1633_ | _1632_;
	assign _1635_ = _1634_ | _1631_;
	assign _1636_ = _1635_ | _1628_;
	assign _1637_ = ~(\mchip.DUT.huff_tree[5] [15] ^ \mchip.DUT.huff_tree[2] [4]);
	assign _1638_ = \mchip.DUT.huff_tree[5] [16] ^ \mchip.DUT.huff_tree[2] [5];
	assign _1639_ = _1637_ & ~_1638_;
	assign _1640_ = \mchip.DUT.huff_tree[5] [18] ^ \mchip.DUT.huff_tree[2] [7];
	assign _1641_ = \mchip.DUT.huff_tree[5] [17] ^ \mchip.DUT.huff_tree[2] [6];
	assign _1642_ = _1641_ | _1640_;
	assign _1643_ = _1639_ & ~_1642_;
	assign _1644_ = \mchip.DUT.huff_tree[5] [19] ^ \mchip.DUT.huff_tree[2] [8];
	assign _1645_ = _1643_ & ~_1644_;
	assign _1646_ = _1636_ & ~_1645_;
	assign _1647_ = _1300_ & ~_1646_;
	assign _1648_ = _1627_ & ~_1647_;
	assign _1649_ = \mchip.DUT.huff_tree[5] [19] ^ \mchip.DUT.huff_tree[3] [13];
	assign _1650_ = \mchip.DUT.huff_tree[5] [18] ^ \mchip.DUT.huff_tree[3] [12];
	assign _1651_ = \mchip.DUT.huff_tree[5] [17] ^ \mchip.DUT.huff_tree[3] [11];
	assign _1652_ = _1651_ | _1650_;
	assign _1653_ = \mchip.DUT.huff_tree[5] [16] ^ \mchip.DUT.huff_tree[3] [10];
	assign _1654_ = \mchip.DUT.huff_tree[5] [15] ^ \mchip.DUT.huff_tree[3] [9];
	assign _1655_ = _1654_ | _1653_;
	assign _1656_ = _1655_ | _1652_;
	assign _1657_ = _1656_ | _1649_;
	assign _1658_ = ~(\mchip.DUT.huff_tree[5] [15] ^ \mchip.DUT.huff_tree[3] [4]);
	assign _1659_ = \mchip.DUT.huff_tree[5] [16] ^ \mchip.DUT.huff_tree[3] [5];
	assign _1660_ = _1658_ & ~_1659_;
	assign _1661_ = \mchip.DUT.huff_tree[5] [18] ^ \mchip.DUT.huff_tree[3] [7];
	assign _1662_ = \mchip.DUT.huff_tree[5] [17] ^ \mchip.DUT.huff_tree[3] [6];
	assign _1663_ = _1662_ | _1661_;
	assign _1664_ = _1660_ & ~_1663_;
	assign _1665_ = \mchip.DUT.huff_tree[5] [19] ^ \mchip.DUT.huff_tree[3] [8];
	assign _1666_ = _1664_ & ~_1665_;
	assign _1667_ = _1657_ & ~_1666_;
	assign _1668_ = _1322_ & ~_1667_;
	assign _1669_ = _1668_ | _1648_;
	assign _1670_ = \mchip.DUT.huff_tree[5] [19] ^ \mchip.DUT.huff_tree[4] [13];
	assign _1671_ = \mchip.DUT.huff_tree[5] [18] ^ \mchip.DUT.huff_tree[4] [12];
	assign _1672_ = \mchip.DUT.huff_tree[5] [17] ^ \mchip.DUT.huff_tree[4] [11];
	assign _1673_ = _1672_ | _1671_;
	assign _1674_ = \mchip.DUT.huff_tree[5] [16] ^ \mchip.DUT.huff_tree[4] [10];
	assign _1675_ = \mchip.DUT.huff_tree[5] [15] ^ \mchip.DUT.huff_tree[4] [9];
	assign _1676_ = _1675_ | _1674_;
	assign _1677_ = _1676_ | _1673_;
	assign _1678_ = _1677_ | _1670_;
	assign _1679_ = ~(\mchip.DUT.huff_tree[5] [15] ^ \mchip.DUT.huff_tree[4] [4]);
	assign _1680_ = \mchip.DUT.huff_tree[5] [16] ^ \mchip.DUT.huff_tree[4] [5];
	assign _1681_ = _1679_ & ~_1680_;
	assign _1682_ = \mchip.DUT.huff_tree[5] [18] ^ \mchip.DUT.huff_tree[4] [7];
	assign _1683_ = \mchip.DUT.huff_tree[5] [17] ^ \mchip.DUT.huff_tree[4] [6];
	assign _1684_ = _1683_ | _1682_;
	assign _1685_ = _1681_ & ~_1684_;
	assign _1686_ = \mchip.DUT.huff_tree[5] [19] ^ \mchip.DUT.huff_tree[4] [8];
	assign _1687_ = _1685_ & ~_1686_;
	assign _1688_ = _1678_ & ~_1687_;
	assign _1689_ = _1344_ & ~_1688_;
	assign _1690_ = _1669_ & ~_1689_;
	assign _1691_ = \mchip.DUT.huff_tree[5] [19] ^ \mchip.DUT.huff_tree[5] [13];
	assign _1692_ = \mchip.DUT.huff_tree[5] [18] ^ \mchip.DUT.huff_tree[5] [12];
	assign _1693_ = \mchip.DUT.huff_tree[5] [17] ^ \mchip.DUT.huff_tree[5] [11];
	assign _1694_ = _1693_ | _1692_;
	assign _1695_ = \mchip.DUT.huff_tree[5] [16] ^ \mchip.DUT.huff_tree[5] [10];
	assign _1696_ = \mchip.DUT.huff_tree[5] [15] ^ \mchip.DUT.huff_tree[5] [9];
	assign _1697_ = _1696_ | _1695_;
	assign _1698_ = _1697_ | _1694_;
	assign _1699_ = _1698_ | _1691_;
	assign _1700_ = ~(\mchip.DUT.huff_tree[5] [15] ^ \mchip.DUT.huff_tree[5] [4]);
	assign _1701_ = \mchip.DUT.huff_tree[5] [16] ^ \mchip.DUT.huff_tree[5] [5];
	assign _1702_ = _1700_ & ~_1701_;
	assign _1703_ = \mchip.DUT.huff_tree[5] [18] ^ \mchip.DUT.huff_tree[5] [7];
	assign _1704_ = \mchip.DUT.huff_tree[5] [17] ^ \mchip.DUT.huff_tree[5] [6];
	assign _1705_ = _1704_ | _1703_;
	assign _1706_ = _1702_ & ~_1705_;
	assign _1707_ = \mchip.DUT.huff_tree[5] [19] ^ \mchip.DUT.huff_tree[5] [8];
	assign _1708_ = _1706_ & ~_1707_;
	assign _1709_ = _1699_ & ~_1708_;
	assign _1710_ = _1366_ & ~_1709_;
	assign _0020_ = _1710_ | _1690_;
	assign _1711_ = \mchip.DUT.huff_tree[5] [3] & ~_1626_;
	assign _1712_ = _1711_ | _1647_;
	assign _1713_ = ~(_1712_ | _1668_);
	assign _1714_ = _1713_ | _1689_;
	assign _0041_ = ~(_1714_ | _1710_);
	assign _1774_[0] = ~\mchip.DUT.b [0];
	assign _1715_ = ~(_0038_ & _0019_);
	assign _1716_ = _0019_ | ~_0038_;
	assign _1717_ = ~(_1716_ & _1715_);
	assign _1718_ = ~\mchip.DUT.huff_tree[3] [0];
	assign _1719_ = _1715_ | _1718_;
	assign _1720_ = \mchip.DUT.huff_tree[2] [0] & ~_1716_;
	assign _1721_ = _1719_ & ~_1720_;
	assign _1722_ = _1717_ & ~_1721_;
	assign _1766_[0] = ~_1722_;
	assign _1723_ = ~(_0039_ & _0018_);
	assign _1724_ = _0039_ & ~_0018_;
	assign _1725_ = _1724_ | ~_1723_;
	assign _1726_ = _1723_ | _1718_;
	assign _1727_ = _1724_ & ~_1722_;
	assign _1728_ = _1726_ & ~_1727_;
	assign _1768_[0] = _1728_ | ~_1725_;
	assign _1729_ = ~(_0041_ & _0020_);
	assign _1730_ = _0041_ & ~_0020_;
	assign _1731_ = _1730_ | ~_1729_;
	assign _1732_ = _1722_ | ~_1730_;
	assign _1733_ = _1768_[0] & ~_1729_;
	assign _1734_ = _1732_ & ~_1733_;
	assign _1735_ = _1731_ & ~_1734_;
	assign _1772_[0] = ~_1735_;
	assign _1736_ = ~(_0040_ & _0017_);
	assign _1737_ = _0040_ & ~_0017_;
	assign _1738_ = _1737_ | ~_1736_;
	assign _1739_ = _1722_ | ~_1737_;
	assign _1740_ = _1768_[0] & ~_1736_;
	assign _1741_ = _1739_ & ~_1740_;
	assign _1742_ = _1738_ & ~_1741_;
	assign _1770_[0] = ~_1742_;
	assign _1743_ = \mchip.DUT.c [0] & \mchip.DUT.c [1];
	assign _1744_ = _1743_ & ~\mchip.DUT.c [2];
	assign _1745_ = _1744_ | io_in[13];
	assign _1746_ = \mchip.DUT.state [0] & ~_1745_;
	assign _1747_ = ~\mchip.DUT.a [2];
	assign _1748_ = \mchip.DUT.a [0] & \mchip.DUT.a [1];
	assign _1749_ = _1747_ & ~_1748_;
	assign _1750_ = _1749_ | io_in[13];
	assign _1751_ = \mchip.DUT.state [6] & ~_1750_;
	assign _1752_ = _1751_ | io_in[13];
	assign _0004_ = _1752_ | _1746_;
	assign _1753_ = ~(\mchip.DUT.count [1] & \mchip.DUT.count [0]);
	assign _0007_ = \mchip.DUT.state [1] & ~_1753_;
	assign _1754_ = \mchip.DUT.state [2] & ~io_in[13];
	assign _1755_ = \mchip.DUT.count [0] & ~\mchip.DUT.count [1];
	assign _1756_ = _1755_ | io_in[13];
	assign _1757_ = \mchip.DUT.state [1] & ~_1756_;
	assign _0005_ = _1757_ | _1754_;
	assign _1758_ = \mchip.DUT.state [3] & ~io_in[13];
	assign _1759_ = ~io_in[13];
	assign _1760_ = ~(_1749_ & _1759_);
	assign _1761_ = \mchip.DUT.state [6] & ~_1760_;
	assign _0006_ = _1761_ | _1758_;
	assign _1762_ = \mchip.DUT.count [0] | ~\mchip.DUT.count [1];
	assign _0008_ = \mchip.DUT.state [1] & ~_1762_;
	assign _0199_ = ~(\mchip.DUT.state [0] | \mchip.DUT.state [6]);
	assign _0009_ = (\mchip.DUT.state [0] ? io_in[11] : \mchip.DUT.state [6]);
	assign _0010_ = (\mchip.DUT.state [6] ? \mchip.DUT.b [0] : \mchip.DUT.state [0]);
	assign _1763_ = \mchip.DUT.huff_tree[1] [18] ^ \mchip.DUT.data_in [19];
	assign _1764_ = \mchip.DUT.huff_tree[1] [17] ^ \mchip.DUT.data_in [18];
	assign _1765_ = _1764_ | _1763_;
	assign _0200_ = \mchip.DUT.huff_tree[1] [16] ^ \mchip.DUT.data_in [17];
	assign _0201_ = \mchip.DUT.huff_tree[1] [15] ^ \mchip.DUT.data_in [16];
	assign _0202_ = _0201_ | _0200_;
	assign _0203_ = _0202_ | _1765_;
	assign _0204_ = _0203_ | \mchip.DUT.huff_tree[1] [19];
	assign _0205_ = _0204_ | _1278_;
	assign _0206_ = \mchip.DUT.data_in [19] ^ \mchip.DUT.huff_tree[2] [18];
	assign _0207_ = \mchip.DUT.data_in [18] ^ \mchip.DUT.huff_tree[2] [17];
	assign _0208_ = _0207_ | _0206_;
	assign _0209_ = \mchip.DUT.data_in [17] ^ \mchip.DUT.huff_tree[2] [16];
	assign _0210_ = \mchip.DUT.data_in [16] ^ \mchip.DUT.huff_tree[2] [15];
	assign _0211_ = _0210_ | _0209_;
	assign _0212_ = _0211_ | _0208_;
	assign _0213_ = _0212_ | \mchip.DUT.huff_tree[2] [19];
	assign _0214_ = \mchip.DUT.huff_tree[2] [14] & ~_0213_;
	assign _0215_ = _0205_ & ~_0214_;
	assign _0216_ = \mchip.DUT.data_in [19] ^ \mchip.DUT.huff_tree[4] [18];
	assign _0217_ = \mchip.DUT.data_in [18] ^ \mchip.DUT.huff_tree[4] [17];
	assign _0218_ = _0217_ | _0216_;
	assign _0219_ = \mchip.DUT.data_in [17] ^ \mchip.DUT.huff_tree[4] [16];
	assign _0220_ = \mchip.DUT.data_in [16] ^ \mchip.DUT.huff_tree[4] [15];
	assign _0221_ = _0220_ | _0219_;
	assign _0222_ = _0221_ | _0218_;
	assign _0223_ = _0222_ | \mchip.DUT.huff_tree[4] [19];
	assign _0224_ = \mchip.DUT.huff_tree[4] [14] & ~_0223_;
	assign _0225_ = \mchip.DUT.data_in [19] ^ \mchip.DUT.huff_tree[3] [18];
	assign _0226_ = \mchip.DUT.data_in [18] ^ \mchip.DUT.huff_tree[3] [17];
	assign _0227_ = _0226_ | _0225_;
	assign _0228_ = \mchip.DUT.data_in [17] ^ \mchip.DUT.huff_tree[3] [16];
	assign _0229_ = \mchip.DUT.data_in [16] ^ \mchip.DUT.huff_tree[3] [15];
	assign _0230_ = _0229_ | _0228_;
	assign _0231_ = _0230_ | _0227_;
	assign _0232_ = _0231_ | \mchip.DUT.huff_tree[3] [19];
	assign _0233_ = \mchip.DUT.huff_tree[3] [14] & ~_0232_;
	assign _0234_ = _0233_ | _0224_;
	assign _0235_ = _0215_ & ~_0234_;
	assign _0236_ = \mchip.DUT.data_in [19] ^ \mchip.DUT.huff_tree[5] [18];
	assign _0237_ = \mchip.DUT.data_in [18] ^ \mchip.DUT.huff_tree[5] [17];
	assign _0238_ = _0237_ | _0236_;
	assign _0239_ = \mchip.DUT.data_in [17] ^ \mchip.DUT.huff_tree[5] [16];
	assign _0240_ = \mchip.DUT.data_in [16] ^ \mchip.DUT.huff_tree[5] [15];
	assign _0241_ = _0240_ | _0239_;
	assign _0242_ = _0241_ | _0238_;
	assign _0243_ = _0242_ | \mchip.DUT.huff_tree[5] [19];
	assign _0244_ = \mchip.DUT.huff_tree[5] [14] & ~_0243_;
	assign _0245_ = _0235_ & ~_0244_;
	assign _0011_ = \mchip.DUT.state [3] & ~_0245_;
	assign _0246_ = \mchip.DUT.data_in [11] ^ \mchip.DUT.huff_tree[1] [18];
	assign _0247_ = \mchip.DUT.data_in [10] ^ \mchip.DUT.huff_tree[1] [17];
	assign _0248_ = _0247_ | _0246_;
	assign _0249_ = \mchip.DUT.data_in [9] ^ \mchip.DUT.huff_tree[1] [16];
	assign _0250_ = \mchip.DUT.data_in [8] ^ \mchip.DUT.huff_tree[1] [15];
	assign _0251_ = _0250_ | _0249_;
	assign _0252_ = _0251_ | _0248_;
	assign _0253_ = _0252_ | \mchip.DUT.huff_tree[1] [19];
	assign _0254_ = _0253_ | _1278_;
	assign _0255_ = \mchip.DUT.data_in [11] ^ \mchip.DUT.huff_tree[2] [18];
	assign _0256_ = \mchip.DUT.data_in [10] ^ \mchip.DUT.huff_tree[2] [17];
	assign _0257_ = _0256_ | _0255_;
	assign _0258_ = \mchip.DUT.data_in [9] ^ \mchip.DUT.huff_tree[2] [16];
	assign _0259_ = \mchip.DUT.data_in [8] ^ \mchip.DUT.huff_tree[2] [15];
	assign _0260_ = _0259_ | _0258_;
	assign _0261_ = _0260_ | _0257_;
	assign _0262_ = _0261_ | \mchip.DUT.huff_tree[2] [19];
	assign _0263_ = \mchip.DUT.huff_tree[2] [14] & ~_0262_;
	assign _0264_ = _0254_ & ~_0263_;
	assign _0265_ = \mchip.DUT.data_in [11] ^ \mchip.DUT.huff_tree[4] [18];
	assign _0266_ = \mchip.DUT.data_in [10] ^ \mchip.DUT.huff_tree[4] [17];
	assign _0267_ = _0266_ | _0265_;
	assign _0268_ = \mchip.DUT.data_in [9] ^ \mchip.DUT.huff_tree[4] [16];
	assign _0269_ = \mchip.DUT.data_in [8] ^ \mchip.DUT.huff_tree[4] [15];
	assign _0270_ = _0269_ | _0268_;
	assign _0271_ = _0270_ | _0267_;
	assign _0272_ = _0271_ | \mchip.DUT.huff_tree[4] [19];
	assign _0273_ = \mchip.DUT.huff_tree[4] [14] & ~_0272_;
	assign _0274_ = \mchip.DUT.data_in [11] ^ \mchip.DUT.huff_tree[3] [18];
	assign _0275_ = \mchip.DUT.data_in [10] ^ \mchip.DUT.huff_tree[3] [17];
	assign _0276_ = _0275_ | _0274_;
	assign _0277_ = \mchip.DUT.data_in [9] ^ \mchip.DUT.huff_tree[3] [16];
	assign _0278_ = \mchip.DUT.data_in [8] ^ \mchip.DUT.huff_tree[3] [15];
	assign _0279_ = _0278_ | _0277_;
	assign _0280_ = _0279_ | _0276_;
	assign _0281_ = _0280_ | \mchip.DUT.huff_tree[3] [19];
	assign _0282_ = \mchip.DUT.huff_tree[3] [14] & ~_0281_;
	assign _0283_ = _0282_ | _0273_;
	assign _0284_ = _0264_ & ~_0283_;
	assign _0285_ = \mchip.DUT.data_in [11] ^ \mchip.DUT.huff_tree[5] [18];
	assign _0286_ = \mchip.DUT.data_in [10] ^ \mchip.DUT.huff_tree[5] [17];
	assign _0287_ = _0286_ | _0285_;
	assign _0288_ = \mchip.DUT.data_in [9] ^ \mchip.DUT.huff_tree[5] [16];
	assign _0289_ = \mchip.DUT.data_in [8] ^ \mchip.DUT.huff_tree[5] [15];
	assign _0290_ = _0289_ | _0288_;
	assign _0291_ = _0290_ | _0287_;
	assign _0292_ = _0291_ | \mchip.DUT.huff_tree[5] [19];
	assign _0293_ = \mchip.DUT.huff_tree[5] [14] & ~_0292_;
	assign _0294_ = _0284_ & ~_0293_;
	assign _0012_ = \mchip.DUT.state [3] & ~_0294_;
	assign _0295_ = \mchip.DUT.data_in [3] ^ \mchip.DUT.huff_tree[1] [18];
	assign _0296_ = \mchip.DUT.data_in [2] ^ \mchip.DUT.huff_tree[1] [17];
	assign _0297_ = _0296_ | _0295_;
	assign _0298_ = \mchip.DUT.data_in [1] ^ \mchip.DUT.huff_tree[1] [16];
	assign _0299_ = \mchip.DUT.data_in [0] ^ \mchip.DUT.huff_tree[1] [15];
	assign _0300_ = _0299_ | _0298_;
	assign _0301_ = _0300_ | _0297_;
	assign _0302_ = _0301_ | \mchip.DUT.huff_tree[1] [19];
	assign _0303_ = _0302_ | _1278_;
	assign _0304_ = \mchip.DUT.data_in [3] ^ \mchip.DUT.huff_tree[2] [18];
	assign _0305_ = \mchip.DUT.data_in [2] ^ \mchip.DUT.huff_tree[2] [17];
	assign _0306_ = _0305_ | _0304_;
	assign _0307_ = \mchip.DUT.data_in [1] ^ \mchip.DUT.huff_tree[2] [16];
	assign _0308_ = \mchip.DUT.data_in [0] ^ \mchip.DUT.huff_tree[2] [15];
	assign _0309_ = _0308_ | _0307_;
	assign _0310_ = _0309_ | _0306_;
	assign _0311_ = _0310_ | \mchip.DUT.huff_tree[2] [19];
	assign _0312_ = \mchip.DUT.huff_tree[2] [14] & ~_0311_;
	assign _0313_ = _0303_ & ~_0312_;
	assign _0314_ = \mchip.DUT.data_in [3] ^ \mchip.DUT.huff_tree[4] [18];
	assign _0315_ = \mchip.DUT.data_in [2] ^ \mchip.DUT.huff_tree[4] [17];
	assign _0316_ = _0315_ | _0314_;
	assign _0317_ = \mchip.DUT.data_in [1] ^ \mchip.DUT.huff_tree[4] [16];
	assign _0318_ = \mchip.DUT.data_in [0] ^ \mchip.DUT.huff_tree[4] [15];
	assign _0319_ = _0318_ | _0317_;
	assign _0320_ = _0319_ | _0316_;
	assign _0321_ = _0320_ | \mchip.DUT.huff_tree[4] [19];
	assign _0322_ = \mchip.DUT.huff_tree[4] [14] & ~_0321_;
	assign _0323_ = \mchip.DUT.data_in [3] ^ \mchip.DUT.huff_tree[3] [18];
	assign _0324_ = \mchip.DUT.data_in [2] ^ \mchip.DUT.huff_tree[3] [17];
	assign _0325_ = _0324_ | _0323_;
	assign _0326_ = \mchip.DUT.data_in [1] ^ \mchip.DUT.huff_tree[3] [16];
	assign _0327_ = \mchip.DUT.data_in [0] ^ \mchip.DUT.huff_tree[3] [15];
	assign _0328_ = _0327_ | _0326_;
	assign _0329_ = _0328_ | _0325_;
	assign _0330_ = _0329_ | \mchip.DUT.huff_tree[3] [19];
	assign _0331_ = \mchip.DUT.huff_tree[3] [14] & ~_0330_;
	assign _0332_ = _0331_ | _0322_;
	assign _0333_ = _0313_ & ~_0332_;
	assign _0334_ = \mchip.DUT.data_in [3] ^ \mchip.DUT.huff_tree[5] [18];
	assign _0335_ = \mchip.DUT.data_in [2] ^ \mchip.DUT.huff_tree[5] [17];
	assign _0336_ = _0335_ | _0334_;
	assign _0337_ = \mchip.DUT.data_in [1] ^ \mchip.DUT.huff_tree[5] [16];
	assign _0338_ = \mchip.DUT.data_in [0] ^ \mchip.DUT.huff_tree[5] [15];
	assign _0339_ = _0338_ | _0337_;
	assign _0340_ = _0339_ | _0336_;
	assign _0341_ = _0340_ | \mchip.DUT.huff_tree[5] [19];
	assign _0342_ = \mchip.DUT.huff_tree[5] [14] & ~_0341_;
	assign _0343_ = _0333_ & ~_0342_;
	assign _0013_ = \mchip.DUT.state [3] & ~_0343_;
	assign _0198_ = ~(\mchip.DUT.state [2] | \mchip.DUT.state [1]);
	assign _0014_ = _1759_ & ~_0198_;
	assign _0344_ = io_in[13] | ~io_in[11];
	assign _0015_ = \mchip.DUT.state [0] & ~_0344_;
	assign _0016_ = _1759_ & ~_0199_;
	assign _0345_ = _1748_ & ~_1747_;
	assign _0346_ = _0345_ | _1749_;
	assign _0347_ = \mchip.DUT.a [0] & ~_0346_;
	assign _0348_ = ~(\mchip.DUT.a [0] ^ \mchip.DUT.a [1]);
	assign _0349_ = ~_0348_;
	assign _0350_ = _0349_ ^ _1749_;
	assign _0351_ = _0350_ & _0347_;
	assign _0352_ = _0348_ & ~_1749_;
	assign _0353_ = _0352_ ^ _0345_;
	assign _0354_ = _0353_ ^ _0351_;
	assign _0355_ = ~\mchip.DUT.a [0];
	assign _0356_ = ~_0345_;
	assign _0357_ = _0352_ & ~_0356_;
	assign _0358_ = _0353_ & _0351_;
	assign _0359_ = _0358_ | _0357_;
	assign _0360_ = ~(_0345_ | _1749_);
	assign _0361_ = _0360_ ^ _0359_;
	assign _0362_ = _0361_ | ~\mchip.DUT.character [14];
	assign _0363_ = _0355_ & ~_0362_;
	assign _0364_ = \mchip.DUT.character [12] & ~_0361_;
	assign _0365_ = \mchip.DUT.character [13] & ~_0361_;
	assign _0366_ = (\mchip.DUT.a [0] ? _0365_ : _0364_);
	assign _0367_ = (_0348_ ? _0363_ : _0366_);
	assign _0368_ = ~_0367_;
	assign _0369_ = _0346_ ^ _0355_;
	assign _0370_ = \mchip.DUT.character [10] & ~_0361_;
	assign _0371_ = \mchip.DUT.character [11] & ~_0361_;
	assign _0372_ = (\mchip.DUT.a [0] ? _0371_ : _0370_);
	assign _0373_ = \mchip.DUT.character [8] & ~_0361_;
	assign _0374_ = \mchip.DUT.character [9] & ~_0361_;
	assign _0375_ = (\mchip.DUT.a [0] ? _0374_ : _0373_);
	assign _0376_ = (_0348_ ? _0372_ : _0375_);
	assign _0377_ = ~_0376_;
	assign _0378_ = (_0369_ ? _0368_ : _0377_);
	assign _0379_ = _0350_ ^ _0347_;
	assign _0380_ = \mchip.DUT.character [6] & ~_0361_;
	assign _0381_ = \mchip.DUT.character [7] & ~_0361_;
	assign _0382_ = (\mchip.DUT.a [0] ? _0381_ : _0380_);
	assign _0383_ = \mchip.DUT.character [4] & ~_0361_;
	assign _0384_ = \mchip.DUT.character [5] & ~_0361_;
	assign _0385_ = (\mchip.DUT.a [0] ? _0384_ : _0383_);
	assign _0386_ = (_0348_ ? _0382_ : _0385_);
	assign _0387_ = ~_0386_;
	assign _0388_ = \mchip.DUT.character [2] & ~_0361_;
	assign _0389_ = \mchip.DUT.character [3] & ~_0361_;
	assign _0390_ = (\mchip.DUT.a [0] ? _0389_ : _0388_);
	assign _0391_ = ~_0390_;
	assign _0392_ = _0361_ | ~\mchip.DUT.character [0];
	assign _0393_ = \mchip.DUT.character [1] & ~_0361_;
	assign _0394_ = ~_0393_;
	assign _0395_ = (\mchip.DUT.a [0] ? _0394_ : _0392_);
	assign _0396_ = (_0348_ ? _0391_ : _0395_);
	assign _0397_ = (_0369_ ? _0387_ : _0396_);
	assign _0398_ = (_0379_ ? _0378_ : _0397_);
	assign _0399_ = ~(_0398_ | _0354_);
	assign _0400_ = ~(_0348_ ^ _0346_);
	assign _0401_ = ~(_0400_ & _0345_);
	assign _0402_ = _1748_ & ~_0401_;
	assign _0403_ = _0346_ & ~_0402_;
	assign _0404_ = _0400_ ^ _1748_;
	assign _0405_ = ~(_1749_ & \mchip.DUT.encoded_value [8]);
	assign _0406_ = _0405_ | \mchip.DUT.a [0];
	assign _0407_ = _0348_ ^ \mchip.DUT.a [0];
	assign _0408_ = _0407_ | _0406_;
	assign _0409_ = _0408_ | _0404_;
	assign _0410_ = ~_1748_;
	assign _0411_ = (\mchip.DUT.a [2] ? _0349_ : _0410_);
	assign _0412_ = _0411_ ^ _0356_;
	assign _0413_ = ~(_1749_ & \mchip.DUT.encoded_value [6]);
	assign _0414_ = ~(_1749_ & \mchip.DUT.encoded_value [7]);
	assign _0415_ = (\mchip.DUT.a [0] ? _0414_ : _0413_);
	assign _0416_ = ~(_1749_ & \mchip.DUT.encoded_value [4]);
	assign _0417_ = ~(_1749_ & \mchip.DUT.encoded_value [5]);
	assign _0418_ = (\mchip.DUT.a [0] ? _0417_ : _0416_);
	assign _0419_ = (_0407_ ? _0415_ : _0418_);
	assign _0420_ = ~(_1749_ & \mchip.DUT.encoded_value [2]);
	assign _0421_ = ~(_1749_ & \mchip.DUT.encoded_value [3]);
	assign _0422_ = (\mchip.DUT.a [0] ? _0421_ : _0420_);
	assign _0423_ = ~(_1749_ & \mchip.DUT.encoded_value [0]);
	assign _0424_ = ~(_1749_ & \mchip.DUT.encoded_value [1]);
	assign _0425_ = (\mchip.DUT.a [0] ? _0424_ : _0423_);
	assign _0426_ = (_0407_ ? _0422_ : _0425_);
	assign _0427_ = (_0404_ ? _0419_ : _0426_);
	assign _0428_ = (_0412_ ? _0409_ : _0427_);
	assign _0429_ = _0403_ & ~_0428_;
	assign _0021_ = (\mchip.DUT.b [0] ? _0429_ : _0399_);
	assign _0430_ = ~_0369_;
	assign _0431_ = ~(_0361_ & \mchip.DUT.character [0]);
	assign _0432_ = _0431_ | _0355_;
	assign _0433_ = _0432_ | ~_0348_;
	assign _0434_ = _0433_ | _0430_;
	assign _0435_ = _0379_ & ~_0434_;
	assign _0436_ = ~_0365_;
	assign _0437_ = (\mchip.DUT.a [0] ? _0362_ : _0436_);
	assign _0438_ = ~(_0437_ | _0348_);
	assign _0439_ = (\mchip.DUT.a [0] ? _0364_ : _0371_);
	assign _0440_ = (\mchip.DUT.a [0] ? _0370_ : _0374_);
	assign _0441_ = (_0348_ ? _0439_ : _0440_);
	assign _0442_ = (_0369_ ? _0438_ : _0441_);
	assign _0443_ = (\mchip.DUT.a [0] ? _0373_ : _0381_);
	assign _0444_ = (\mchip.DUT.a [0] ? _0380_ : _0384_);
	assign _0445_ = (_0348_ ? _0443_ : _0444_);
	assign _0446_ = (\mchip.DUT.a [0] ? _0383_ : _0389_);
	assign _0447_ = (\mchip.DUT.a [0] ? _0388_ : _0393_);
	assign _0448_ = (_0348_ ? _0446_ : _0447_);
	assign _0449_ = (_0369_ ? _0445_ : _0448_);
	assign _0450_ = (_0379_ ? _0442_ : _0449_);
	assign _0451_ = (_0354_ ? _0435_ : _0450_);
	assign _0452_ = ~_0412_;
	assign _0453_ = ~_0407_;
	assign _0454_ = _1749_ | ~\mchip.DUT.encoded_value [0];
	assign _0455_ = _0454_ | _0355_;
	assign _0456_ = _0455_ | _0453_;
	assign _0457_ = _0404_ & ~_0456_;
	assign _0458_ = (\mchip.DUT.a [0] ? _0405_ : _0414_);
	assign _0459_ = (\mchip.DUT.a [0] ? _0413_ : _0417_);
	assign _0460_ = (_0407_ ? _0458_ : _0459_);
	assign _0461_ = (\mchip.DUT.a [0] ? _0416_ : _0421_);
	assign _0462_ = (\mchip.DUT.a [0] ? _0420_ : _0424_);
	assign _0463_ = (_0407_ ? _0461_ : _0462_);
	assign _0464_ = (_0404_ ? _0460_ : _0463_);
	assign _0465_ = (_0403_ ? _0464_ : _0457_);
	assign _0466_ = _0452_ & ~_0465_;
	assign _0022_ = (\mchip.DUT.b [0] ? _0466_ : _0451_);
	assign _0467_ = ~(_0361_ & \mchip.DUT.character [1]);
	assign _0468_ = (\mchip.DUT.a [0] ? _0467_ : _0431_);
	assign _0469_ = _0468_ | ~_0348_;
	assign _0470_ = _0469_ | _0430_;
	assign _0471_ = _0379_ & ~_0470_;
	assign _0472_ = _0363_ & ~_0348_;
	assign _0473_ = (_0348_ ? _0366_ : _0372_);
	assign _0474_ = (_0369_ ? _0472_ : _0473_);
	assign _0475_ = (_0348_ ? _0375_ : _0382_);
	assign _0476_ = (_0348_ ? _0385_ : _0390_);
	assign _0477_ = (_0369_ ? _0475_ : _0476_);
	assign _0478_ = (_0379_ ? _0474_ : _0477_);
	assign _0479_ = (_0354_ ? _0471_ : _0478_);
	assign _0480_ = _1749_ | ~\mchip.DUT.encoded_value [1];
	assign _0481_ = (\mchip.DUT.a [0] ? _0480_ : _0454_);
	assign _0482_ = _0481_ | _0453_;
	assign _0483_ = _0404_ & ~_0482_;
	assign _0484_ = (_0407_ ? _0406_ : _0415_);
	assign _0485_ = (_0407_ ? _0418_ : _0422_);
	assign _0486_ = (_0404_ ? _0484_ : _0485_);
	assign _0487_ = (_0403_ ? _0486_ : _0483_);
	assign _0488_ = _0452_ & ~_0487_;
	assign _0023_ = (\mchip.DUT.b [0] ? _0488_ : _0479_);
	assign _0489_ = ~(_0361_ & \mchip.DUT.character [2]);
	assign _0490_ = (\mchip.DUT.a [0] ? _0489_ : _0467_);
	assign _0491_ = (_0348_ ? _0490_ : _0432_);
	assign _0492_ = _0491_ | ~_0369_;
	assign _0493_ = _0379_ & ~_0492_;
	assign _0494_ = ~_0439_;
	assign _0495_ = (_0348_ ? _0437_ : _0494_);
	assign _0496_ = _0430_ & ~_0495_;
	assign _0497_ = (_0348_ ? _0440_ : _0443_);
	assign _0498_ = (_0348_ ? _0444_ : _0446_);
	assign _0499_ = (_0369_ ? _0497_ : _0498_);
	assign _0500_ = (_0379_ ? _0496_ : _0499_);
	assign _0501_ = (_0354_ ? _0493_ : _0500_);
	assign _0502_ = ~(_1749_ & \mchip.DUT.encoded_mask [8]);
	assign _0503_ = _0502_ | \mchip.DUT.a [0];
	assign _0504_ = _0503_ | _0407_;
	assign _0505_ = _0504_ | _0404_;
	assign _0506_ = ~(_1749_ & \mchip.DUT.encoded_mask [6]);
	assign _0507_ = ~(_1749_ & \mchip.DUT.encoded_mask [7]);
	assign _0508_ = (\mchip.DUT.a [0] ? _0507_ : _0506_);
	assign _0509_ = ~(_1749_ & \mchip.DUT.encoded_mask [4]);
	assign _0510_ = ~(_1749_ & \mchip.DUT.encoded_mask [5]);
	assign _0511_ = (\mchip.DUT.a [0] ? _0510_ : _0509_);
	assign _0512_ = (_0407_ ? _0508_ : _0511_);
	assign _0513_ = ~(_1749_ & \mchip.DUT.encoded_mask [2]);
	assign _0514_ = ~(_1749_ & \mchip.DUT.encoded_mask [3]);
	assign _0515_ = (\mchip.DUT.a [0] ? _0514_ : _0513_);
	assign _0516_ = ~(_1749_ & \mchip.DUT.encoded_mask [0]);
	assign _0517_ = ~(_1749_ & \mchip.DUT.encoded_mask [1]);
	assign _0518_ = (\mchip.DUT.a [0] ? _0517_ : _0516_);
	assign _0519_ = (_0407_ ? _0515_ : _0518_);
	assign _0520_ = (_0404_ ? _0512_ : _0519_);
	assign _0521_ = (_0412_ ? _0505_ : _0520_);
	assign _0522_ = _0403_ & ~_0521_;
	assign _0024_ = (\mchip.DUT.b [0] ? _0522_ : _0501_);
	assign _0523_ = ~(_0361_ & \mchip.DUT.character [3]);
	assign _0524_ = (\mchip.DUT.a [0] ? _0523_ : _0489_);
	assign _0525_ = (_0348_ ? _0524_ : _0468_);
	assign _0526_ = _0525_ | ~_0369_;
	assign _0527_ = _0379_ & ~_0526_;
	assign _0528_ = _0367_ & ~_0369_;
	assign _0529_ = (_0369_ ? _0376_ : _0386_);
	assign _0530_ = (_0379_ ? _0528_ : _0529_);
	assign _0531_ = (_0354_ ? _0527_ : _0530_);
	assign _0532_ = _1749_ | ~\mchip.DUT.encoded_mask [0];
	assign _0533_ = _0532_ | _0355_;
	assign _0534_ = _0533_ | _0453_;
	assign _0535_ = _0404_ & ~_0534_;
	assign _0536_ = (\mchip.DUT.a [0] ? _0502_ : _0507_);
	assign _0537_ = (\mchip.DUT.a [0] ? _0506_ : _0510_);
	assign _0538_ = (_0407_ ? _0536_ : _0537_);
	assign _0539_ = (\mchip.DUT.a [0] ? _0509_ : _0514_);
	assign _0540_ = (\mchip.DUT.a [0] ? _0513_ : _0517_);
	assign _0541_ = (_0407_ ? _0539_ : _0540_);
	assign _0542_ = (_0404_ ? _0538_ : _0541_);
	assign _0543_ = (_0403_ ? _0542_ : _0535_);
	assign _0544_ = _0452_ & ~_0543_;
	assign _0025_ = (\mchip.DUT.b [0] ? _0544_ : _0531_);
	assign _0545_ = _1749_ | ~\mchip.DUT.encoded_mask [1];
	assign _0546_ = (\mchip.DUT.a [0] ? _0545_ : _0532_);
	assign _0547_ = _0546_ | _0453_;
	assign _0548_ = _0404_ & ~_0547_;
	assign _0549_ = (_0407_ ? _0503_ : _0508_);
	assign _0550_ = (_0407_ ? _0511_ : _0515_);
	assign _0551_ = (_0404_ ? _0549_ : _0550_);
	assign _0552_ = (_0403_ ? _0551_ : _0548_);
	assign _0553_ = _0452_ & ~_0552_;
	assign _0026_ = _0553_ | _1774_[0];
	assign _0554_ = \mchip.DUT.huff_tree[5] [2] & ~\mchip.DUT.huff_tree[5] [3];
	assign _0555_ = ~(_0554_ | \mchip.DUT.encoded_value_h[5] [0]);
	assign _0096_ = ~(_0555_ & _0554_);
	assign _0556_ = \mchip.DUT.huff_tree[2] [2] & ~\mchip.DUT.huff_tree[2] [3];
	assign _0557_ = _0556_ | ~\mchip.DUT.encoded_value_h[2] [0];
	assign _1776_[2] = _0556_ & ~_0557_;
	assign _0558_ = \mchip.DUT.huff_tree[3] [2] & ~\mchip.DUT.huff_tree[3] [3];
	assign _0559_ = ~(_0558_ | \mchip.DUT.encoded_value_h[3] [0]);
	assign _1776_[0] = ~(_0559_ & _0558_);
	assign _0560_ = \mchip.DUT.huff_tree[4] [2] & ~\mchip.DUT.huff_tree[4] [3];
	assign _0561_ = _0560_ | ~\mchip.DUT.encoded_value_h[4] [0];
	assign _0093_ = _0560_ & ~_0561_;
	assign _0562_ = ~_1776_[2];
	assign _0563_ = _0312_ & ~_0562_;
	assign _0564_ = (_0331_ ? _1776_[0] : _0563_);
	assign _0565_ = (_0322_ ? _0093_ : _0564_);
	assign _0050_ = (_0342_ ? _0096_ : _0565_);
	assign _0566_ = \mchip.DUT.huff_tree[5] [3] & \mchip.DUT.huff_tree[5] [2];
	assign _0097_ = (_0554_ ? \mchip.DUT.encoded_value_h[5] [1] : _0566_);
	assign _0567_ = \mchip.DUT.huff_tree[2] [3] & \mchip.DUT.huff_tree[2] [2];
	assign _0568_ = \mchip.DUT.huff_tree[2] [3] & ~\mchip.DUT.huff_tree[2] [2];
	assign _0569_ = ~(_0568_ | _0567_);
	assign _0570_ = ~_0569_;
	assign _0571_ = ~(_0568_ & \mchip.DUT.encoded_value_h[2] [0]);
	assign _0572_ = _0567_ & \mchip.DUT.encoded_value_h[3] [0];
	assign _0573_ = _0571_ & ~_0572_;
	assign _0574_ = _0570_ & ~_0573_;
	assign _1776_[3] = (_0556_ ? \mchip.DUT.encoded_value_h[2] [1] : _0574_);
	assign _0575_ = \mchip.DUT.huff_tree[3] [3] & \mchip.DUT.huff_tree[3] [2];
	assign _0576_ = \mchip.DUT.huff_tree[3] [3] & ~\mchip.DUT.huff_tree[3] [2];
	assign _0577_ = _0576_ | _0575_;
	assign _0578_ = ~(_0576_ & _1776_[2]);
	assign _0579_ = _0575_ & \mchip.DUT.encoded_value_h[3] [0];
	assign _0580_ = _0578_ & ~_0579_;
	assign _0581_ = _0577_ & ~_0580_;
	assign _1776_[1] = (_0558_ ? \mchip.DUT.encoded_value_h[3] [1] : _0581_);
	assign _0582_ = \mchip.DUT.huff_tree[4] [3] & \mchip.DUT.huff_tree[4] [2];
	assign _0094_ = (_0560_ ? \mchip.DUT.encoded_value_h[4] [1] : _0582_);
	assign _0583_ = _1776_[3] & _0312_;
	assign _0584_ = (_0331_ ? _1776_[1] : _0583_);
	assign _0585_ = (_0322_ ? _0094_ : _0584_);
	assign _0051_ = (_0342_ ? _0097_ : _0585_);
	assign _0586_ = \mchip.DUT.huff_tree[5] [3] & ~\mchip.DUT.huff_tree[5] [2];
	assign _0587_ = _0566_ | _0586_;
	assign _0588_ = ~(_1776_[3] & _0586_);
	assign _0589_ = _1776_[1] & _0566_;
	assign _0590_ = _0588_ & ~_0589_;
	assign _0591_ = _0587_ & ~_0590_;
	assign _0098_ = (_0554_ ? \mchip.DUT.encoded_value_h[5] [2] : _0591_);
	assign _0592_ = ~(_0567_ & \mchip.DUT.encoded_value_h[3] [1]);
	assign _0593_ = _0568_ & \mchip.DUT.encoded_value_h[2] [1];
	assign _0594_ = _0592_ & ~_0593_;
	assign _0595_ = _0570_ & ~_0594_;
	assign _0091_ = (_0556_ ? \mchip.DUT.encoded_value_h[2] [2] : _0595_);
	assign _0596_ = ~(_0575_ & \mchip.DUT.encoded_value_h[3] [1]);
	assign _0597_ = _0576_ & _1776_[3];
	assign _0598_ = _0596_ & ~_0597_;
	assign _0599_ = _0577_ & ~_0598_;
	assign _0092_ = (_0558_ ? \mchip.DUT.encoded_value_h[3] [2] : _0599_);
	assign _0600_ = \mchip.DUT.huff_tree[4] [3] & ~\mchip.DUT.huff_tree[4] [2];
	assign _0601_ = _0582_ | _0600_;
	assign _0602_ = ~(_0600_ & _1776_[3]);
	assign _0603_ = _0582_ & _1776_[1];
	assign _0604_ = _0602_ & ~_0603_;
	assign _0605_ = _0601_ & ~_0604_;
	assign _0095_ = (_0560_ ? \mchip.DUT.encoded_value_h[4] [2] : _0605_);
	assign _0606_ = _0091_ & _0312_;
	assign _0607_ = (_0331_ ? _0092_ : _0606_);
	assign _0608_ = (_0322_ ? _0095_ : _0607_);
	assign _0052_ = (_0342_ ? _0098_ : _0608_);
	assign _0609_ = ~(\mchip.DUT.huff_tree[2] [1] | \mchip.DUT.huff_tree[2] [0]);
	assign _0610_ = _0312_ & ~_0609_;
	assign _0611_ = \mchip.DUT.huff_tree[3] [1] | \mchip.DUT.huff_tree[3] [0];
	assign _0612_ = (_0331_ ? _0611_ : _0610_);
	assign _0613_ = \mchip.DUT.huff_tree[4] [0] | \mchip.DUT.huff_tree[4] [1];
	assign _0614_ = (_0322_ ? _0613_ : _0612_);
	assign _0615_ = \mchip.DUT.huff_tree[5] [0] | \mchip.DUT.huff_tree[5] [1];
	assign _0047_ = (_0342_ ? _0615_ : _0614_);
	assign _0616_ = \mchip.DUT.huff_tree[2] [0] & ~\mchip.DUT.huff_tree[2] [1];
	assign _0617_ = _0616_ ^ _0609_;
	assign _0618_ = _0312_ & ~_0617_;
	assign _0619_ = \mchip.DUT.huff_tree[3] [0] & ~\mchip.DUT.huff_tree[3] [1];
	assign _0620_ = _0619_ ^ _0611_;
	assign _0621_ = (_0331_ ? _0620_ : _0618_);
	assign _0622_ = \mchip.DUT.huff_tree[4] [0] & ~\mchip.DUT.huff_tree[4] [1];
	assign _0623_ = _0622_ ^ _0613_;
	assign _0624_ = (_0322_ ? _0623_ : _0621_);
	assign _0625_ = \mchip.DUT.huff_tree[5] [0] & ~\mchip.DUT.huff_tree[5] [1];
	assign _0626_ = _0625_ ^ _0615_;
	assign _0048_ = (_0342_ ? _0626_ : _0624_);
	assign _0627_ = ~(\mchip.DUT.huff_tree[2] [1] & \mchip.DUT.huff_tree[2] [0]);
	assign _0628_ = _0312_ & ~_0627_;
	assign _0629_ = \mchip.DUT.huff_tree[3] [1] & \mchip.DUT.huff_tree[3] [0];
	assign _0630_ = (_0331_ ? _0629_ : _0628_);
	assign _0631_ = \mchip.DUT.huff_tree[4] [0] & \mchip.DUT.huff_tree[4] [1];
	assign _0632_ = (_0322_ ? _0631_ : _0630_);
	assign _0633_ = \mchip.DUT.huff_tree[5] [0] & \mchip.DUT.huff_tree[5] [1];
	assign _0049_ = (_0342_ ? _0633_ : _0632_);
	assign _0634_ = (_0263_ ? \mchip.DUT.huff_tree[2] [15] : \mchip.DUT.huff_tree[1] [15]);
	assign _0635_ = (_0282_ ? \mchip.DUT.huff_tree[3] [15] : _0634_);
	assign _0636_ = (_0273_ ? \mchip.DUT.huff_tree[4] [15] : _0635_);
	assign _0027_ = (_0293_ ? \mchip.DUT.huff_tree[5] [15] : _0636_);
	assign _0637_ = (_0263_ ? \mchip.DUT.huff_tree[2] [16] : \mchip.DUT.huff_tree[1] [16]);
	assign _0638_ = (_0282_ ? \mchip.DUT.huff_tree[3] [16] : _0637_);
	assign _0639_ = (_0273_ ? \mchip.DUT.huff_tree[4] [16] : _0638_);
	assign _0028_ = (_0293_ ? \mchip.DUT.huff_tree[5] [16] : _0639_);
	assign _0640_ = (_0263_ ? \mchip.DUT.huff_tree[2] [17] : \mchip.DUT.huff_tree[1] [17]);
	assign _0641_ = (_0282_ ? \mchip.DUT.huff_tree[3] [17] : _0640_);
	assign _0642_ = (_0273_ ? \mchip.DUT.huff_tree[4] [17] : _0641_);
	assign _0029_ = (_0293_ ? \mchip.DUT.huff_tree[5] [17] : _0642_);
	assign _0643_ = (_0263_ ? \mchip.DUT.huff_tree[2] [18] : \mchip.DUT.huff_tree[1] [18]);
	assign _0644_ = (_0282_ ? \mchip.DUT.huff_tree[3] [18] : _0643_);
	assign _0645_ = (_0273_ ? \mchip.DUT.huff_tree[4] [18] : _0644_);
	assign _0030_ = (_0293_ ? \mchip.DUT.huff_tree[5] [18] : _0645_);
	assign _0646_ = (_0263_ ? \mchip.DUT.huff_tree[2] [19] : \mchip.DUT.huff_tree[1] [19]);
	assign _0647_ = (_0282_ ? \mchip.DUT.huff_tree[3] [19] : _0646_);
	assign _0648_ = (_0273_ ? \mchip.DUT.huff_tree[4] [19] : _0647_);
	assign _0031_ = (_0293_ ? \mchip.DUT.huff_tree[5] [19] : _0648_);
	assign _0649_ = _0263_ & ~_0562_;
	assign _0650_ = (_0282_ ? _1776_[0] : _0649_);
	assign _0651_ = (_0273_ ? _0093_ : _0650_);
	assign _0035_ = (_0293_ ? _0096_ : _0651_);
	assign _0652_ = _1776_[3] & _0263_;
	assign _0653_ = (_0282_ ? _1776_[1] : _0652_);
	assign _0654_ = (_0273_ ? _0094_ : _0653_);
	assign _0036_ = (_0293_ ? _0097_ : _0654_);
	assign _0655_ = _0091_ & _0263_;
	assign _0656_ = (_0282_ ? _0092_ : _0655_);
	assign _0657_ = (_0273_ ? _0095_ : _0656_);
	assign _0037_ = (_0293_ ? _0098_ : _0657_);
	assign _0658_ = _0263_ & ~_0609_;
	assign _0659_ = (_0282_ ? _0611_ : _0658_);
	assign _0660_ = (_0273_ ? _0613_ : _0659_);
	assign _0032_ = (_0293_ ? _0615_ : _0660_);
	assign _0661_ = _0263_ & ~_0617_;
	assign _0662_ = (_0282_ ? _0620_ : _0661_);
	assign _0663_ = (_0273_ ? _0623_ : _0662_);
	assign _0033_ = (_0293_ ? _0626_ : _0663_);
	assign _0664_ = _0263_ & ~_0627_;
	assign _0665_ = (_0282_ ? _0629_ : _0664_);
	assign _0666_ = (_0273_ ? _0631_ : _0665_);
	assign _0034_ = (_0293_ ? _0633_ : _0666_);
	assign _0667_ = (_0214_ ? \mchip.DUT.huff_tree[2] [15] : \mchip.DUT.huff_tree[1] [15]);
	assign _0668_ = (_0233_ ? \mchip.DUT.huff_tree[3] [15] : _0667_);
	assign _0669_ = (_0224_ ? \mchip.DUT.huff_tree[4] [15] : _0668_);
	assign _0099_ = (_0244_ ? \mchip.DUT.huff_tree[5] [15] : _0669_);
	assign _0670_ = (_0214_ ? \mchip.DUT.huff_tree[2] [16] : \mchip.DUT.huff_tree[1] [16]);
	assign _0671_ = (_0233_ ? \mchip.DUT.huff_tree[3] [16] : _0670_);
	assign _0672_ = (_0224_ ? \mchip.DUT.huff_tree[4] [16] : _0671_);
	assign _0100_ = (_0244_ ? \mchip.DUT.huff_tree[5] [16] : _0672_);
	assign _0673_ = (_0214_ ? \mchip.DUT.huff_tree[2] [17] : \mchip.DUT.huff_tree[1] [17]);
	assign _0674_ = (_0233_ ? \mchip.DUT.huff_tree[3] [17] : _0673_);
	assign _0675_ = (_0224_ ? \mchip.DUT.huff_tree[4] [17] : _0674_);
	assign _0101_ = (_0244_ ? \mchip.DUT.huff_tree[5] [17] : _0675_);
	assign _0676_ = (_0214_ ? \mchip.DUT.huff_tree[2] [18] : \mchip.DUT.huff_tree[1] [18]);
	assign _0677_ = (_0233_ ? \mchip.DUT.huff_tree[3] [18] : _0676_);
	assign _0678_ = (_0224_ ? \mchip.DUT.huff_tree[4] [18] : _0677_);
	assign _0102_ = (_0244_ ? \mchip.DUT.huff_tree[5] [18] : _0678_);
	assign _0679_ = (_0214_ ? \mchip.DUT.huff_tree[2] [19] : \mchip.DUT.huff_tree[1] [19]);
	assign _0680_ = (_0233_ ? \mchip.DUT.huff_tree[3] [19] : _0679_);
	assign _0681_ = (_0224_ ? \mchip.DUT.huff_tree[4] [19] : _0680_);
	assign _0103_ = (_0244_ ? \mchip.DUT.huff_tree[5] [19] : _0681_);
	assign _0682_ = _0214_ & ~_0562_;
	assign _0683_ = (_0233_ ? _1776_[0] : _0682_);
	assign _0684_ = (_0224_ ? _0093_ : _0683_);
	assign _0107_ = (_0244_ ? _0096_ : _0684_);
	assign _0685_ = _1776_[3] & _0214_;
	assign _0686_ = (_0233_ ? _1776_[1] : _0685_);
	assign _0687_ = (_0224_ ? _0094_ : _0686_);
	assign _0108_ = (_0244_ ? _0097_ : _0687_);
	assign _0688_ = _0091_ & _0214_;
	assign _0689_ = (_0233_ ? _0092_ : _0688_);
	assign _0690_ = (_0224_ ? _0095_ : _0689_);
	assign _0109_ = (_0244_ ? _0098_ : _0690_);
	assign _0691_ = _0214_ & ~_0609_;
	assign _0692_ = (_0233_ ? _0611_ : _0691_);
	assign _0693_ = (_0224_ ? _0613_ : _0692_);
	assign _0104_ = (_0244_ ? _0615_ : _0693_);
	assign _0694_ = _0214_ & ~_0617_;
	assign _0695_ = (_0233_ ? _0620_ : _0694_);
	assign _0696_ = (_0224_ ? _0623_ : _0695_);
	assign _0105_ = (_0244_ ? _0626_ : _0696_);
	assign _0697_ = _0214_ & ~_0627_;
	assign _0698_ = (_0233_ ? _0629_ : _0697_);
	assign _0699_ = (_0224_ ? _0631_ : _0698_);
	assign _0106_ = (_0244_ ? _0633_ : _0699_);
	assign _0053_ = \mchip.DUT.node_sorter_ins.output_node [0] & \mchip.DUT.state [1];
	assign _0054_ = \mchip.DUT.node_sorter_ins.output_node [1] & \mchip.DUT.state [1];
	assign _0055_ = \mchip.DUT.node_sorter_ins.output_node [2] & \mchip.DUT.state [1];
	assign _0056_ = \mchip.DUT.node_sorter_ins.output_node [3] & \mchip.DUT.state [1];
	assign _0057_ = \mchip.DUT.node_sorter_ins.output_node [4] & \mchip.DUT.state [1];
	assign _0058_ = \mchip.DUT.node_sorter_ins.output_node [5] & \mchip.DUT.state [1];
	assign _0059_ = \mchip.DUT.node_sorter_ins.output_node [6] & \mchip.DUT.state [1];
	assign _0060_ = \mchip.DUT.node_sorter_ins.output_node [7] & \mchip.DUT.state [1];
	assign _0061_ = \mchip.DUT.node_sorter_ins.output_node [8] & \mchip.DUT.state [1];
	assign _0062_ = \mchip.DUT.node_sorter_ins.output_node [9] & \mchip.DUT.state [1];
	assign _0063_ = \mchip.DUT.node_sorter_ins.output_node [10] | ~\mchip.DUT.state [1];
	assign _0064_ = (\mchip.DUT.state [1] ? \mchip.DUT.node_sorter_ins.output_node [11] : \mchip.DUT.freq_in [3]);
	assign _0065_ = (\mchip.DUT.state [1] ? \mchip.DUT.node_sorter_ins.output_node [12] : \mchip.DUT.freq_in [4]);
	assign _0066_ = (\mchip.DUT.state [1] ? \mchip.DUT.node_sorter_ins.output_node [13] : \mchip.DUT.freq_in [5]);
	assign _0067_ = (\mchip.DUT.state [1] ? \mchip.DUT.node_sorter_ins.output_node [14] : \mchip.DUT.data_in [8]);
	assign _0068_ = (\mchip.DUT.state [1] ? \mchip.DUT.node_sorter_ins.output_node [15] : \mchip.DUT.data_in [9]);
	assign _0069_ = (\mchip.DUT.state [1] ? \mchip.DUT.node_sorter_ins.output_node [16] : \mchip.DUT.data_in [10]);
	assign _0070_ = (\mchip.DUT.state [1] ? \mchip.DUT.node_sorter_ins.output_node [17] : \mchip.DUT.data_in [11]);
	assign _0071_ = (\mchip.DUT.state [1] ? \mchip.DUT.node_sorter_ins.output_node [18] : \mchip.DUT.data_in [12]);
	assign _0072_ = \mchip.DUT.node_sorter_ins.output_node [33] & \mchip.DUT.state [1];
	assign _0073_ = \mchip.DUT.node_sorter_ins.output_node [34] & \mchip.DUT.state [1];
	assign _0074_ = \mchip.DUT.node_sorter_ins.output_node [35] & \mchip.DUT.state [1];
	assign _0075_ = \mchip.DUT.node_sorter_ins.output_node [36] & \mchip.DUT.state [1];
	assign _0076_ = \mchip.DUT.node_sorter_ins.output_node [37] & \mchip.DUT.state [1];
	assign _0077_ = \mchip.DUT.node_sorter_ins.output_node [52] & \mchip.DUT.state [1];
	assign _0078_ = \mchip.DUT.node_sorter_ins.output_node [53] & \mchip.DUT.state [1];
	assign _0079_ = \mchip.DUT.node_sorter_ins.output_node [54] & \mchip.DUT.state [1];
	assign _0080_ = \mchip.DUT.node_sorter_ins.output_node [55] & \mchip.DUT.state [1];
	assign _0081_ = \mchip.DUT.node_sorter_ins.output_node [56] & \mchip.DUT.state [1];
	assign _0082_ = ~\mchip.DUT.state [1];
	assign _0700_ = \mchip.DUT.node_sorter_ins.output_node [49] ^ \mchip.DUT.node_sorter_ins.output_node [30];
	assign _0083_ = (\mchip.DUT.state [1] ? _0700_ : \mchip.DUT.freq_in [6]);
	assign _0701_ = \mchip.DUT.node_sorter_ins.output_node [49] & \mchip.DUT.node_sorter_ins.output_node [30];
	assign _0702_ = ~(\mchip.DUT.node_sorter_ins.output_node [50] ^ \mchip.DUT.node_sorter_ins.output_node [31]);
	assign _0703_ = ~(_0702_ ^ _0701_);
	assign _0084_ = (\mchip.DUT.state [1] ? _0703_ : \mchip.DUT.freq_in [7]);
	assign _0704_ = \mchip.DUT.node_sorter_ins.output_node [50] & \mchip.DUT.node_sorter_ins.output_node [31];
	assign _0705_ = _0701_ & ~_0702_;
	assign _0706_ = _0705_ | _0704_;
	assign _0707_ = \mchip.DUT.node_sorter_ins.output_node [51] ^ \mchip.DUT.node_sorter_ins.output_node [32];
	assign _0708_ = _0707_ ^ _0706_;
	assign _0085_ = (\mchip.DUT.state [1] ? _0708_ : \mchip.DUT.freq_in [8]);
	assign _0709_ = \mchip.DUT.node_sorter_ins.output_node [52] ^ \mchip.DUT.node_sorter_ins.output_node [33];
	assign _0086_ = (\mchip.DUT.state [1] ? _0709_ : \mchip.DUT.data_in [16]);
	assign _0710_ = \mchip.DUT.node_sorter_ins.output_node [52] & \mchip.DUT.node_sorter_ins.output_node [33];
	assign _0711_ = ~(\mchip.DUT.node_sorter_ins.output_node [53] ^ \mchip.DUT.node_sorter_ins.output_node [34]);
	assign _0712_ = ~(_0711_ ^ _0710_);
	assign _0087_ = (\mchip.DUT.state [1] ? _0712_ : \mchip.DUT.data_in [17]);
	assign _0713_ = _0710_ & ~_0711_;
	assign _0714_ = \mchip.DUT.node_sorter_ins.output_node [53] & \mchip.DUT.node_sorter_ins.output_node [34];
	assign _0715_ = _0714_ | _0713_;
	assign _0716_ = \mchip.DUT.node_sorter_ins.output_node [54] ^ \mchip.DUT.node_sorter_ins.output_node [35];
	assign _0717_ = _0716_ ^ _0715_;
	assign _0088_ = (\mchip.DUT.state [1] ? _0717_ : \mchip.DUT.data_in [18]);
	assign _0718_ = \mchip.DUT.node_sorter_ins.output_node [54] & \mchip.DUT.node_sorter_ins.output_node [35];
	assign _0719_ = _0716_ & _0715_;
	assign _0720_ = _0719_ | _0718_;
	assign _0721_ = \mchip.DUT.node_sorter_ins.output_node [55] ^ \mchip.DUT.node_sorter_ins.output_node [36];
	assign _0722_ = _0721_ ^ _0720_;
	assign _0089_ = (\mchip.DUT.state [1] ? _0722_ : \mchip.DUT.data_in [19]);
	assign _0723_ = \mchip.DUT.node_sorter_ins.output_node [55] & \mchip.DUT.node_sorter_ins.output_node [36];
	assign _0724_ = _0721_ & _0718_;
	assign _0725_ = _0724_ | _0723_;
	assign _0726_ = ~(_0721_ & _0716_);
	assign _0727_ = _0715_ & ~_0726_;
	assign _0728_ = _0727_ | _0725_;
	assign _0729_ = \mchip.DUT.node_sorter_ins.output_node [56] ^ \mchip.DUT.node_sorter_ins.output_node [37];
	assign _0730_ = _0729_ ^ _0728_;
	assign _0090_ = (\mchip.DUT.state [1] ? _0730_ : \mchip.DUT.data_in [20]);
	assign _0731_ = (_0312_ ? \mchip.DUT.huff_tree[2] [15] : \mchip.DUT.huff_tree[1] [15]);
	assign _0732_ = (_0331_ ? \mchip.DUT.huff_tree[3] [15] : _0731_);
	assign _0733_ = (_0322_ ? \mchip.DUT.huff_tree[4] [15] : _0732_);
	assign _0042_ = (_0342_ ? \mchip.DUT.huff_tree[5] [15] : _0733_);
	assign _0734_ = (_0312_ ? \mchip.DUT.huff_tree[2] [16] : \mchip.DUT.huff_tree[1] [16]);
	assign _0735_ = (_0331_ ? \mchip.DUT.huff_tree[3] [16] : _0734_);
	assign _0736_ = (_0322_ ? \mchip.DUT.huff_tree[4] [16] : _0735_);
	assign _0043_ = (_0342_ ? \mchip.DUT.huff_tree[5] [16] : _0736_);
	assign _0737_ = (_0312_ ? \mchip.DUT.huff_tree[2] [17] : \mchip.DUT.huff_tree[1] [17]);
	assign _0738_ = (_0331_ ? \mchip.DUT.huff_tree[3] [17] : _0737_);
	assign _0739_ = (_0322_ ? \mchip.DUT.huff_tree[4] [17] : _0738_);
	assign _0044_ = (_0342_ ? \mchip.DUT.huff_tree[5] [17] : _0739_);
	assign _0740_ = (_0312_ ? \mchip.DUT.huff_tree[2] [18] : \mchip.DUT.huff_tree[1] [18]);
	assign _0741_ = (_0331_ ? \mchip.DUT.huff_tree[3] [18] : _0740_);
	assign _0742_ = (_0322_ ? \mchip.DUT.huff_tree[4] [18] : _0741_);
	assign _0045_ = (_0342_ ? \mchip.DUT.huff_tree[5] [18] : _0742_);
	assign _0743_ = (_0312_ ? \mchip.DUT.huff_tree[2] [19] : \mchip.DUT.huff_tree[1] [19]);
	assign _0744_ = (_0331_ ? \mchip.DUT.huff_tree[3] [19] : _0743_);
	assign _0745_ = (_0322_ ? \mchip.DUT.huff_tree[4] [19] : _0744_);
	assign _0046_ = (_0342_ ? \mchip.DUT.huff_tree[5] [19] : _0745_);
	assign _0134_ = ~(\mchip.DUT.c [0] | \mchip.DUT.state [6]);
	assign _0746_ = \mchip.DUT.c [0] ^ \mchip.DUT.c [1];
	assign _0135_ = _0746_ & ~\mchip.DUT.state [6];
	assign _0747_ = ~\mchip.DUT.c [2];
	assign _0748_ = _0747_ & ~_1743_;
	assign _0749_ = _1743_ & ~_0747_;
	assign _0750_ = ~(_0749_ | _0748_);
	assign _0136_ = _0750_ & ~\mchip.DUT.state [6];
	assign _0137_ = \mchip.DUT.state [6] & ~\mchip.DUT.b [0];
	assign _0138_ = \mchip.DUT.state [6] & ~\mchip.DUT.a [0];
	assign _0139_ = \mchip.DUT.state [6] & ~_0348_;
	assign _0140_ = \mchip.DUT.state [6] & ~_0346_;
	assign _0751_ = \mchip.DUT.in_huff_tree [56] | ~\mchip.DUT.in_huff_tree [37];
	assign _0752_ = ~(\mchip.DUT.in_huff_tree [37] ^ \mchip.DUT.in_huff_tree [56]);
	assign _0753_ = \mchip.DUT.in_huff_tree [55] | ~\mchip.DUT.in_huff_tree [36];
	assign _0754_ = ~(\mchip.DUT.in_huff_tree [36] ^ \mchip.DUT.in_huff_tree [55]);
	assign _0755_ = \mchip.DUT.in_huff_tree [54] | ~\mchip.DUT.in_huff_tree [35];
	assign _0756_ = _0754_ & ~_0755_;
	assign _0757_ = _0753_ & ~_0756_;
	assign _0758_ = \mchip.DUT.in_huff_tree [35] ^ \mchip.DUT.in_huff_tree [54];
	assign _0759_ = _0754_ & ~_0758_;
	assign _0760_ = \mchip.DUT.in_huff_tree [53] | ~\mchip.DUT.in_huff_tree [34];
	assign _0761_ = ~(\mchip.DUT.in_huff_tree [34] ^ \mchip.DUT.in_huff_tree [53]);
	assign _0762_ = \mchip.DUT.in_huff_tree [52] & ~\mchip.DUT.in_huff_tree [33];
	assign _0763_ = _0761_ & ~_0762_;
	assign _0764_ = _0760_ & ~_0763_;
	assign _0765_ = _0759_ & ~_0764_;
	assign _0766_ = _0757_ & ~_0765_;
	assign _0767_ = _0752_ & ~_0766_;
	assign _0768_ = _0751_ & ~_0767_;
	assign _0769_ = ~(\mchip.DUT.in_huff_tree [31] ^ \mchip.DUT.in_huff_tree [50]);
	assign _0770_ = ~(\mchip.DUT.in_huff_tree [30] ^ \mchip.DUT.in_huff_tree [49]);
	assign _0771_ = _0770_ & _0769_;
	assign _0772_ = ~(\mchip.DUT.in_huff_tree [32] ^ \mchip.DUT.in_huff_tree [51]);
	assign _0773_ = ~(_0772_ & _0771_);
	assign _0774_ = _0768_ & ~_0773_;
	assign _0775_ = \mchip.DUT.in_huff_tree [51] | ~\mchip.DUT.in_huff_tree [32];
	assign _0776_ = \mchip.DUT.in_huff_tree [50] | ~\mchip.DUT.in_huff_tree [31];
	assign _0777_ = \mchip.DUT.in_huff_tree [49] & ~\mchip.DUT.in_huff_tree [30];
	assign _0778_ = _0769_ & ~_0777_;
	assign _0779_ = _0776_ & ~_0778_;
	assign _0780_ = _0772_ & ~_0779_;
	assign _0781_ = _0775_ & ~_0780_;
	assign _0782_ = _0781_ | _0774_;
	assign _0783_ = (_0782_ ? \mchip.DUT.in_huff_tree [38] : \mchip.DUT.in_huff_tree [19]);
	assign _0784_ = ~(\mchip.DUT.in_huff_tree [32] | \mchip.DUT.in_huff_tree [51]);
	assign _0785_ = ~(_0784_ & \mchip.DUT.in_huff_tree [13]);
	assign _0786_ = (_0782_ ? \mchip.DUT.in_huff_tree [50] : \mchip.DUT.in_huff_tree [31]);
	assign _0787_ = _0786_ | ~\mchip.DUT.in_huff_tree [12];
	assign _0788_ = (_0782_ ? \mchip.DUT.in_huff_tree [49] : \mchip.DUT.in_huff_tree [30]);
	assign _0789_ = \mchip.DUT.in_huff_tree [11] | ~_0788_;
	assign _0790_ = _0786_ ^ \mchip.DUT.in_huff_tree [12];
	assign _0791_ = _0789_ & ~_0790_;
	assign _0792_ = _0787_ & ~_0791_;
	assign _0793_ = _0784_ ^ \mchip.DUT.in_huff_tree [13];
	assign _0794_ = _0793_ & ~_0792_;
	assign _0795_ = _0785_ & ~_0794_;
	assign _0796_ = _0788_ ^ \mchip.DUT.in_huff_tree [11];
	assign _0797_ = _0796_ | _0790_;
	assign _0798_ = _0793_ & ~_0797_;
	assign _0799_ = (_0782_ ? \mchip.DUT.in_huff_tree [56] : \mchip.DUT.in_huff_tree [37]);
	assign _0800_ = _0799_ ^ \mchip.DUT.in_huff_tree [18];
	assign _0801_ = ~\mchip.DUT.in_huff_tree [17];
	assign _0802_ = (_0782_ ? \mchip.DUT.in_huff_tree [55] : \mchip.DUT.in_huff_tree [36]);
	assign _0803_ = _0802_ | _0801_;
	assign _0804_ = _0802_ ^ _0801_;
	assign _0805_ = (_0782_ ? \mchip.DUT.in_huff_tree [54] : \mchip.DUT.in_huff_tree [35]);
	assign _0806_ = _0805_ | ~\mchip.DUT.in_huff_tree [16];
	assign _0807_ = _0804_ & ~_0806_;
	assign _0808_ = _0803_ & ~_0807_;
	assign _0809_ = _0805_ ^ \mchip.DUT.in_huff_tree [16];
	assign _0810_ = _0804_ & ~_0809_;
	assign _0811_ = ~\mchip.DUT.in_huff_tree [15];
	assign _0812_ = (_0782_ ? \mchip.DUT.in_huff_tree [53] : \mchip.DUT.in_huff_tree [34]);
	assign _0813_ = _0812_ | _0811_;
	assign _0814_ = _0812_ ^ _0811_;
	assign _0815_ = ~\mchip.DUT.in_huff_tree [14];
	assign _0816_ = ~\mchip.DUT.in_huff_tree [52];
	assign _0817_ = ~\mchip.DUT.in_huff_tree [33];
	assign _0818_ = (_0782_ ? _0816_ : _0817_);
	assign _0819_ = _0815_ & ~_0818_;
	assign _0820_ = _0814_ & ~_0819_;
	assign _0821_ = _0813_ & ~_0820_;
	assign _0822_ = _0810_ & ~_0821_;
	assign _0823_ = _0808_ & ~_0822_;
	assign _0824_ = _0823_ | _0800_;
	assign _0825_ = \mchip.DUT.in_huff_tree [18] & ~_0799_;
	assign _0826_ = _0824_ & ~_0825_;
	assign _0827_ = _0826_ & _0798_;
	assign _0828_ = _0827_ | _0795_;
	assign _0829_ = _0783_ & ~_0828_;
	assign _0830_ = (_0782_ ? \mchip.DUT.in_huff_tree [37] : \mchip.DUT.in_huff_tree [56]);
	assign _0831_ = ~_0830_;
	assign _0832_ = ~\mchip.DUT.in_huff_tree [18];
	assign _0833_ = ~_0799_;
	assign _0834_ = (_0828_ ? _0832_ : _0833_);
	assign _0835_ = _0834_ ^ _0831_;
	assign _0836_ = (_0782_ ? \mchip.DUT.in_huff_tree [36] : \mchip.DUT.in_huff_tree [55]);
	assign _0837_ = ~_0802_;
	assign _0838_ = (_0828_ ? _0801_ : _0837_);
	assign _0839_ = _0838_ | _0836_;
	assign _0840_ = _0838_ ^ _0836_;
	assign _0841_ = (_0782_ ? \mchip.DUT.in_huff_tree [35] : \mchip.DUT.in_huff_tree [54]);
	assign _0842_ = (_0828_ ? \mchip.DUT.in_huff_tree [16] : _0805_);
	assign _0843_ = _0841_ | ~_0842_;
	assign _0844_ = _0840_ & ~_0843_;
	assign _0845_ = _0839_ & ~_0844_;
	assign _0846_ = _0842_ ^ _0841_;
	assign _0847_ = _0840_ & ~_0846_;
	assign _0848_ = (_0782_ ? \mchip.DUT.in_huff_tree [34] : \mchip.DUT.in_huff_tree [53]);
	assign _0849_ = ~_0812_;
	assign _0850_ = (_0828_ ? _0811_ : _0849_);
	assign _0851_ = _0850_ | _0848_;
	assign _0852_ = _0850_ ^ _0848_;
	assign _0853_ = (_0828_ ? _0815_ : _0818_);
	assign _0854_ = (_0782_ ? \mchip.DUT.in_huff_tree [33] : \mchip.DUT.in_huff_tree [52]);
	assign _0855_ = _0854_ & _0853_;
	assign _0856_ = _0852_ & ~_0855_;
	assign _0857_ = _0851_ & ~_0856_;
	assign _0858_ = _0847_ & ~_0857_;
	assign _0859_ = _0845_ & ~_0858_;
	assign _0860_ = _0859_ | _0835_;
	assign _0861_ = _0831_ & ~_0834_;
	assign _0862_ = _0860_ & ~_0861_;
	assign _0863_ = \mchip.DUT.in_huff_tree [32] & \mchip.DUT.in_huff_tree [51];
	assign _0864_ = ~_0784_;
	assign _0865_ = (_0828_ ? \mchip.DUT.in_huff_tree [13] : _0864_);
	assign _0866_ = ~(_0865_ ^ _0863_);
	assign _0867_ = (_0782_ ? \mchip.DUT.in_huff_tree [31] : \mchip.DUT.in_huff_tree [50]);
	assign _0868_ = (_0828_ ? \mchip.DUT.in_huff_tree [12] : _0786_);
	assign _0869_ = ~(_0868_ ^ _0867_);
	assign _0870_ = (_0782_ ? \mchip.DUT.in_huff_tree [30] : \mchip.DUT.in_huff_tree [49]);
	assign _0871_ = (_0828_ ? \mchip.DUT.in_huff_tree [11] : _0788_);
	assign _0872_ = ~(_0871_ ^ _0870_);
	assign _0873_ = _0872_ & _0869_;
	assign _0874_ = ~(_0873_ & _0866_);
	assign _0875_ = _0862_ & ~_0874_;
	assign _0876_ = _0863_ | ~_0865_;
	assign _0877_ = _0867_ | ~_0868_;
	assign _0878_ = _0870_ & ~_0871_;
	assign _0879_ = _0869_ & ~_0878_;
	assign _0880_ = _0877_ & ~_0879_;
	assign _0881_ = _0866_ & ~_0880_;
	assign _0882_ = _0876_ & ~_0881_;
	assign _0883_ = _0882_ | _0875_;
	assign _0884_ = (_0782_ ? \mchip.DUT.in_huff_tree [19] : \mchip.DUT.in_huff_tree [38]);
	assign _0172_ = (_0883_ ? _0829_ : _0884_);
	assign _0885_ = ~\mchip.DUT.in_huff_tree [20];
	assign _0886_ = ~\mchip.DUT.in_huff_tree [39];
	assign _0887_ = (_0782_ ? _0886_ : _0885_);
	assign _0888_ = ~(_0887_ | _0828_);
	assign _0889_ = (_0782_ ? \mchip.DUT.in_huff_tree [20] : \mchip.DUT.in_huff_tree [39]);
	assign _0173_ = (_0883_ ? _0888_ : _0889_);
	assign _0890_ = ~\mchip.DUT.in_huff_tree [21];
	assign _0891_ = ~\mchip.DUT.in_huff_tree [40];
	assign _0892_ = (_0782_ ? _0891_ : _0890_);
	assign _0893_ = ~(_0892_ | _0828_);
	assign _0894_ = (_0782_ ? \mchip.DUT.in_huff_tree [21] : \mchip.DUT.in_huff_tree [40]);
	assign _0175_ = (_0883_ ? _0893_ : _0894_);
	assign _0895_ = ~\mchip.DUT.in_huff_tree [22];
	assign _0896_ = ~\mchip.DUT.in_huff_tree [41];
	assign _0897_ = (_0782_ ? _0896_ : _0895_);
	assign _0898_ = ~(_0897_ | _0828_);
	assign _0899_ = (_0782_ ? \mchip.DUT.in_huff_tree [22] : \mchip.DUT.in_huff_tree [41]);
	assign _0176_ = (_0883_ ? _0898_ : _0899_);
	assign _0900_ = ~\mchip.DUT.in_huff_tree [23];
	assign _0901_ = ~\mchip.DUT.in_huff_tree [42];
	assign _0902_ = (_0782_ ? _0901_ : _0900_);
	assign _0903_ = ~(_0902_ | _0828_);
	assign _0904_ = (_0782_ ? \mchip.DUT.in_huff_tree [23] : \mchip.DUT.in_huff_tree [42]);
	assign _0177_ = (_0883_ ? _0903_ : _0904_);
	assign _0905_ = ~\mchip.DUT.in_huff_tree [24];
	assign _0906_ = ~\mchip.DUT.in_huff_tree [43];
	assign _0907_ = (_0782_ ? _0906_ : _0905_);
	assign _0908_ = ~(_0907_ | _0828_);
	assign _0909_ = (_0782_ ? \mchip.DUT.in_huff_tree [24] : \mchip.DUT.in_huff_tree [43]);
	assign _0178_ = (_0883_ ? _0908_ : _0909_);
	assign _0910_ = ~\mchip.DUT.in_huff_tree [25];
	assign _0911_ = ~\mchip.DUT.in_huff_tree [44];
	assign _0912_ = (_0782_ ? _0911_ : _0910_);
	assign _0913_ = ~(_0912_ | _0828_);
	assign _0914_ = (_0782_ ? \mchip.DUT.in_huff_tree [25] : \mchip.DUT.in_huff_tree [44]);
	assign _0179_ = (_0883_ ? _0913_ : _0914_);
	assign _0915_ = ~\mchip.DUT.in_huff_tree [26];
	assign _0916_ = ~\mchip.DUT.in_huff_tree [45];
	assign _0917_ = (_0782_ ? _0916_ : _0915_);
	assign _0918_ = ~(_0917_ | _0828_);
	assign _0919_ = (_0782_ ? \mchip.DUT.in_huff_tree [26] : \mchip.DUT.in_huff_tree [45]);
	assign _0180_ = (_0883_ ? _0918_ : _0919_);
	assign _0920_ = ~\mchip.DUT.in_huff_tree [27];
	assign _0921_ = ~\mchip.DUT.in_huff_tree [46];
	assign _0922_ = (_0782_ ? _0921_ : _0920_);
	assign _0923_ = ~(_0922_ | _0828_);
	assign _0924_ = (_0782_ ? \mchip.DUT.in_huff_tree [27] : \mchip.DUT.in_huff_tree [46]);
	assign _0181_ = (_0883_ ? _0923_ : _0924_);
	assign _0925_ = ~\mchip.DUT.in_huff_tree [28];
	assign _0926_ = ~\mchip.DUT.in_huff_tree [47];
	assign _0927_ = (_0782_ ? _0926_ : _0925_);
	assign _0928_ = ~(_0927_ | _0828_);
	assign _0929_ = (_0782_ ? \mchip.DUT.in_huff_tree [28] : \mchip.DUT.in_huff_tree [47]);
	assign _0182_ = (_0883_ ? _0928_ : _0929_);
	assign _0930_ = (_0782_ ? \mchip.DUT.in_huff_tree [48] : \mchip.DUT.in_huff_tree [29]);
	assign _0931_ = (_0828_ ? \mchip.DUT.in_huff_tree [10] : _0930_);
	assign _0932_ = (_0782_ ? \mchip.DUT.in_huff_tree [29] : \mchip.DUT.in_huff_tree [48]);
	assign _0183_ = (_0883_ ? _0931_ : _0932_);
	assign _0184_ = (_0883_ ? _0871_ : _0870_);
	assign _0186_ = (_0883_ ? _0868_ : _0867_);
	assign _0187_ = (_0883_ ? _0865_ : _0863_);
	assign _0933_ = ~_0853_;
	assign _0188_ = (_0883_ ? _0933_ : _0854_);
	assign _0934_ = ~_0850_;
	assign _0189_ = (_0883_ ? _0934_ : _0848_);
	assign _0190_ = (_0883_ ? _0842_ : _0841_);
	assign _0935_ = ~_0838_;
	assign _0191_ = (_0883_ ? _0935_ : _0836_);
	assign _0936_ = ~_0834_;
	assign _0192_ = (_0883_ ? _0936_ : _0830_);
	assign _0937_ = (_0883_ ? _0884_ : _0829_);
	assign _0938_ = (_0828_ ? _0864_ : \mchip.DUT.in_huff_tree [13]);
	assign _0939_ = (_0883_ ? _0863_ : _0865_);
	assign _0940_ = _0939_ & ~_0938_;
	assign _0941_ = (_0828_ ? _0786_ : \mchip.DUT.in_huff_tree [12]);
	assign _0942_ = ~_0941_;
	assign _0943_ = ~_0867_;
	assign _0944_ = ~_0868_;
	assign _0945_ = (_0883_ ? _0943_ : _0944_);
	assign _0946_ = _0945_ ^ _0942_;
	assign _0947_ = (_0883_ ? _0870_ : _0871_);
	assign _0948_ = (_0828_ ? _0788_ : \mchip.DUT.in_huff_tree [11]);
	assign _0949_ = _0948_ & ~_0947_;
	assign _0950_ = _0949_ | _0946_;
	assign _0951_ = _0942_ & ~_0945_;
	assign _0952_ = _0950_ & ~_0951_;
	assign _0953_ = _0939_ ^ _0938_;
	assign _0954_ = ~(_0953_ | _0952_);
	assign _0955_ = _0954_ | _0940_;
	assign _0956_ = ~(_0948_ ^ _0947_);
	assign _0957_ = _0956_ & ~_0946_;
	assign _0958_ = _0953_ | ~_0957_;
	assign _0959_ = (_0828_ ? _0833_ : _0832_);
	assign _0960_ = (_0883_ ? _0831_ : _0834_);
	assign _0961_ = _0960_ ^ _0959_;
	assign _0962_ = ~_0818_;
	assign _0963_ = (_0828_ ? _0962_ : \mchip.DUT.in_huff_tree [14]);
	assign _0964_ = (_0883_ ? _0854_ : _0933_);
	assign _0965_ = _0964_ ^ _0963_;
	assign _0966_ = (_0828_ ? _0812_ : \mchip.DUT.in_huff_tree [15]);
	assign _0967_ = (_0883_ ? _0848_ : _0934_);
	assign _0968_ = _0967_ ^ _0966_;
	assign _0969_ = ~(_0968_ | _0965_);
	assign _0970_ = (_0828_ ? _0805_ : \mchip.DUT.in_huff_tree [16]);
	assign _0971_ = (_0883_ ? _0841_ : _0842_);
	assign _0972_ = ~(_0971_ ^ _0970_);
	assign _0973_ = (_0828_ ? _0802_ : \mchip.DUT.in_huff_tree [17]);
	assign _0974_ = ~_0836_;
	assign _0975_ = (_0883_ ? _0974_ : _0838_);
	assign _0976_ = ~(_0975_ ^ _0973_);
	assign _0977_ = _0972_ & ~_0976_;
	assign _0978_ = ~(_0977_ & _0969_);
	assign _0979_ = _0978_ | _0961_;
	assign _0980_ = _0975_ | _0973_;
	assign _0981_ = _0971_ & ~_0970_;
	assign _0982_ = _0981_ & ~_0976_;
	assign _0983_ = _0980_ & ~_0982_;
	assign _0984_ = _0966_ | ~_0967_;
	assign _0985_ = _0964_ | ~_0963_;
	assign _0986_ = _0985_ & ~_0968_;
	assign _0987_ = _0984_ & ~_0986_;
	assign _0988_ = _0977_ & ~_0987_;
	assign _0989_ = _0983_ & ~_0988_;
	assign _0990_ = _0989_ | _0961_;
	assign _0991_ = _0959_ & ~_0960_;
	assign _0992_ = _0990_ & ~_0991_;
	assign _0993_ = _0979_ & ~_0992_;
	assign _0994_ = (_0958_ ? _0955_ : _0993_);
	assign _0995_ = _0828_ & _0783_;
	assign _0141_ = (_0994_ ? _0937_ : _0995_);
	assign _0996_ = (_0883_ ? _0889_ : _0888_);
	assign _0997_ = _0828_ & ~_0887_;
	assign _0152_ = (_0994_ ? _0996_ : _0997_);
	assign _0998_ = (_0883_ ? _0894_ : _0893_);
	assign _0999_ = _0828_ & ~_0892_;
	assign _0163_ = (_0994_ ? _0998_ : _0999_);
	assign _1000_ = (_0883_ ? _0899_ : _0898_);
	assign _1001_ = _0828_ & ~_0897_;
	assign _0174_ = (_0994_ ? _1000_ : _1001_);
	assign _1002_ = (_0883_ ? _0904_ : _0903_);
	assign _1003_ = _0828_ & ~_0902_;
	assign _0185_ = (_0994_ ? _1002_ : _1003_);
	assign _1004_ = (_0883_ ? _0909_ : _0908_);
	assign _1005_ = _0828_ & ~_0907_;
	assign _0193_ = (_0994_ ? _1004_ : _1005_);
	assign _1006_ = (_0883_ ? _0914_ : _0913_);
	assign _1007_ = _0828_ & ~_0912_;
	assign _0194_ = (_0994_ ? _1006_ : _1007_);
	assign _1008_ = (_0883_ ? _0919_ : _0918_);
	assign _1009_ = _0828_ & ~_0917_;
	assign _0195_ = (_0994_ ? _1008_ : _1009_);
	assign _1010_ = (_0883_ ? _0924_ : _0923_);
	assign _1011_ = _0828_ & ~_0922_;
	assign _0196_ = (_0994_ ? _1010_ : _1011_);
	assign _1012_ = (_0883_ ? _0929_ : _0928_);
	assign _1013_ = _0828_ & ~_0927_;
	assign _0197_ = (_0994_ ? _1012_ : _1013_);
	assign _1014_ = (_0883_ ? _0932_ : _0931_);
	assign _1015_ = (_0828_ ? _0930_ : \mchip.DUT.in_huff_tree [10]);
	assign _0142_ = (_0994_ ? _1014_ : _1015_);
	assign _0143_ = (_0994_ ? _0947_ : _0948_);
	assign _1016_ = ~_0945_;
	assign _0144_ = (_0994_ ? _1016_ : _0941_);
	assign _0145_ = _0939_ | _0938_;
	assign _0146_ = (_0994_ ? _0964_ : _0963_);
	assign _0147_ = (_0994_ ? _0967_ : _0966_);
	assign _0148_ = (_0994_ ? _0971_ : _0970_);
	assign _1017_ = ~_0975_;
	assign _0149_ = (_0994_ ? _1017_ : _0973_);
	assign _1018_ = ~_0959_;
	assign _1019_ = ~_0960_;
	assign _0150_ = (_0994_ ? _1019_ : _1018_);
	assign _0151_ = (_0994_ ? _0995_ : _0937_);
	assign _0153_ = (_0994_ ? _0997_ : _0996_);
	assign _0154_ = (_0994_ ? _0999_ : _0998_);
	assign _0155_ = (_0994_ ? _1001_ : _1000_);
	assign _0156_ = (_0994_ ? _1003_ : _1002_);
	assign _0157_ = (_0994_ ? _1005_ : _1004_);
	assign _0158_ = (_0994_ ? _1007_ : _1006_);
	assign _0159_ = (_0994_ ? _1009_ : _1008_);
	assign _0160_ = (_0994_ ? _1011_ : _1010_);
	assign _0161_ = (_0994_ ? _1013_ : _1012_);
	assign _0162_ = (_0994_ ? _1015_ : _1014_);
	assign _0164_ = (_0994_ ? _0948_ : _0947_);
	assign _0165_ = (_0994_ ? _0941_ : _1016_);
	assign _0166_ = _0939_ & _0938_;
	assign _0167_ = (_0994_ ? _0963_ : _0964_);
	assign _0168_ = (_0994_ ? _0966_ : _0967_);
	assign _0169_ = (_0994_ ? _0970_ : _0971_);
	assign _0170_ = (_0994_ ? _0973_ : _1017_);
	assign _0171_ = (_0994_ ? _1018_ : _1019_);
	assign _1020_ = ~(_1744_ & _1759_);
	assign _0001_ = \mchip.DUT.state [0] & ~_1020_;
	assign _0000_ = \mchip.DUT.state [5] & ~io_in[13];
	assign _1021_ = ~(_1755_ & _1759_);
	assign _0003_ = \mchip.DUT.state [1] & ~_1021_;
	assign _1022_ = \mchip.DUT.c [1] & ~\mchip.DUT.c [0];
	assign _1023_ = ~(_1022_ ^ _0750_);
	assign _1024_ = ~_1023_;
	assign _1025_ = ~\mchip.DUT.c [0];
	assign _1026_ = ~(\mchip.DUT.c [0] ^ \mchip.DUT.c [1]);
	assign _1027_ = _1026_ | _0750_;
	assign _1028_ = _1025_ & ~_1027_;
	assign _1029_ = _1028_ ^ _0748_;
	assign _1030_ = ~_1029_;
	assign _1031_ = ~_0748_;
	assign _1032_ = _1027_ | _1031_;
	assign _1033_ = _1025_ & ~_1032_;
	assign _1034_ = _1033_ & ~_1031_;
	assign _1035_ = _1034_ ^ _1030_;
	assign _1036_ = ~(_1033_ | _1031_);
	assign _1037_ = _1036_ ^ _1029_;
	assign _1038_ = ~(_1033_ ^ _1031_);
	assign _1039_ = _1038_ ^ _1029_;
	assign _1040_ = _1028_ & ~_0748_;
	assign _1041_ = _1040_ | _1039_;
	assign _1042_ = _1041_ | _1037_;
	assign _1043_ = _1042_ | _1035_;
	assign _1044_ = _1043_ | ~io_in[0];
	assign _1045_ = _1044_ | _1029_;
	assign _1046_ = _1045_ | \mchip.DUT.c [0];
	assign _1047_ = _1026_ ^ \mchip.DUT.c [0];
	assign _1048_ = _1047_ | _1046_;
	assign _1049_ = _1024_ & ~_1048_;
	assign _1050_ = _1043_ | _1029_;
	assign _1051_ = _1050_ | \mchip.DUT.c [0];
	assign _1052_ = _1051_ | _1047_;
	assign _1053_ = _1024_ & ~_1052_;
	assign _1054_ = \mchip.DUT.data_in [0] & ~_1053_;
	assign _0110_ = _1054_ | _1049_;
	assign _1055_ = _1043_ | ~io_in[1];
	assign _1056_ = _1055_ | _1029_;
	assign _1057_ = _1056_ | \mchip.DUT.c [0];
	assign _1058_ = _1057_ | _1047_;
	assign _1059_ = _1024_ & ~_1058_;
	assign _1060_ = \mchip.DUT.data_in [1] & ~_1053_;
	assign _0118_ = _1060_ | _1059_;
	assign _1061_ = _1043_ | ~io_in[2];
	assign _1062_ = _1061_ | _1029_;
	assign _1063_ = _1062_ | \mchip.DUT.c [0];
	assign _1064_ = _1063_ | _1047_;
	assign _1065_ = _1024_ & ~_1064_;
	assign _1066_ = \mchip.DUT.data_in [2] & ~_1053_;
	assign _0120_ = _1066_ | _1065_;
	assign _1067_ = _1043_ | ~io_in[3];
	assign _1068_ = _1067_ | _1029_;
	assign _1069_ = _1068_ | \mchip.DUT.c [0];
	assign _1070_ = _1069_ | _1047_;
	assign _1071_ = _1024_ & ~_1070_;
	assign _1072_ = \mchip.DUT.data_in [3] & ~_1053_;
	assign _0121_ = _1072_ | _1071_;
	assign _1073_ = _1043_ | ~io_in[4];
	assign _1074_ = _1073_ | _1029_;
	assign _1075_ = _1074_ | \mchip.DUT.c [0];
	assign _1076_ = _1075_ | _1047_;
	assign _1077_ = _1024_ & ~_1076_;
	assign _1078_ = \mchip.DUT.data_in [4] & ~_1053_;
	assign _0122_ = _1078_ | _1077_;
	assign _1079_ = ~_1047_;
	assign _1080_ = _1044_ | _1030_;
	assign _1081_ = _1080_ | _1025_;
	assign _1082_ = _1081_ | _1079_;
	assign _1083_ = _1023_ & ~_1082_;
	assign _1084_ = ~(_0748_ & \mchip.DUT.c [0]);
	assign _1085_ = _1084_ | _1079_;
	assign _1086_ = _1023_ & ~_1085_;
	assign _1087_ = \mchip.DUT.data_in [8] & ~_1086_;
	assign _0123_ = _1087_ | _1083_;
	assign _1088_ = _1055_ | _1030_;
	assign _1089_ = _1088_ | _1025_;
	assign _1090_ = _1089_ | _1079_;
	assign _1091_ = _1023_ & ~_1090_;
	assign _1092_ = \mchip.DUT.data_in [9] & ~_1086_;
	assign _0124_ = _1092_ | _1091_;
	assign _1093_ = _1061_ | _1030_;
	assign _1094_ = _1093_ | _1025_;
	assign _1095_ = _1094_ | _1079_;
	assign _1096_ = _1023_ & ~_1095_;
	assign _1097_ = \mchip.DUT.data_in [10] & ~_1086_;
	assign _0111_ = _1097_ | _1096_;
	assign _1098_ = _1067_ | _1030_;
	assign _1099_ = _1098_ | _1025_;
	assign _1100_ = _1099_ | _1079_;
	assign _1101_ = _1023_ & ~_1100_;
	assign _1102_ = \mchip.DUT.data_in [11] & ~_1086_;
	assign _0112_ = _1102_ | _1101_;
	assign _1103_ = _1073_ | _1030_;
	assign _1104_ = _1103_ | _1025_;
	assign _1105_ = _1104_ | _1079_;
	assign _1106_ = _1023_ & ~_1105_;
	assign _1107_ = \mchip.DUT.data_in [12] & ~_1086_;
	assign _0113_ = _1107_ | _1106_;
	assign _1108_ = _1080_ | \mchip.DUT.c [0];
	assign _1109_ = _1108_ | _1079_;
	assign _1110_ = _1023_ & ~_1109_;
	assign _1111_ = _1043_ | _1030_;
	assign _1112_ = _1111_ | \mchip.DUT.c [0];
	assign _1113_ = _1112_ | _1079_;
	assign _1114_ = _1023_ & ~_1113_;
	assign _1115_ = \mchip.DUT.data_in [16] & ~_1114_;
	assign _0114_ = _1115_ | _1110_;
	assign _1116_ = _1088_ | \mchip.DUT.c [0];
	assign _1117_ = _1116_ | _1079_;
	assign _1118_ = _1023_ & ~_1117_;
	assign _1119_ = \mchip.DUT.data_in [17] & ~_1114_;
	assign _0115_ = _1119_ | _1118_;
	assign _1120_ = _1093_ | \mchip.DUT.c [0];
	assign _1121_ = _1120_ | _1079_;
	assign _1122_ = _1023_ & ~_1121_;
	assign _1123_ = \mchip.DUT.data_in [18] & ~_1114_;
	assign _0116_ = _1123_ | _1122_;
	assign _1124_ = _1098_ | \mchip.DUT.c [0];
	assign _1125_ = _1124_ | _1079_;
	assign _1126_ = _1023_ & ~_1125_;
	assign _1127_ = \mchip.DUT.data_in [19] & ~_1114_;
	assign _0117_ = _1127_ | _1126_;
	assign _1128_ = _1103_ | \mchip.DUT.c [0];
	assign _1129_ = _1128_ | _1079_;
	assign _1130_ = _1023_ & ~_1129_;
	assign _1131_ = \mchip.DUT.data_in [20] & ~_1114_;
	assign _0119_ = _1131_ | _1130_;
	assign _1132_ = _1026_ ^ _0750_;
	assign _1133_ = _1132_ ^ _1743_;
	assign _1134_ = (\mchip.DUT.c [2] ? _1026_ : _1743_);
	assign _1135_ = _1134_ ^ _0749_;
	assign _1136_ = _1135_ | _1133_;
	assign _1137_ = _1022_ & ~_1136_;
	assign _1138_ = ~(_1132_ & _0749_);
	assign _1139_ = _1743_ & ~_1138_;
	assign _1140_ = ~(_1139_ | _0750_);
	assign _1141_ = _1140_ ^ _1137_;
	assign _1142_ = ~(_0748_ & io_in[10]);
	assign _1143_ = _1140_ & _1137_;
	assign _1144_ = ~(_1143_ ^ _1031_);
	assign _1145_ = _1144_ | _1142_;
	assign _1146_ = _1145_ | \mchip.DUT.c [0];
	assign _1147_ = ~(_0748_ & io_in[8]);
	assign _1148_ = _1147_ | _1144_;
	assign _1149_ = ~(_0748_ & io_in[9]);
	assign _1150_ = _1149_ | _1144_;
	assign _1151_ = (\mchip.DUT.c [0] ? _1150_ : _1148_);
	assign _1152_ = (_1026_ ? _1146_ : _1151_);
	assign _1153_ = _0750_ ^ \mchip.DUT.c [0];
	assign _1154_ = _1153_ | _1152_;
	assign _1155_ = _1022_ & ~_1133_;
	assign _1156_ = ~(_1155_ ^ _1135_);
	assign _1157_ = _1156_ | _1154_;
	assign _1158_ = ~(_1157_ | _1141_);
	assign _1159_ = ~_1156_;
	assign _1160_ = ~(_1143_ & _0748_);
	assign _1161_ = _1160_ | \mchip.DUT.c [0];
	assign _1162_ = \mchip.DUT.c [0] & ~_1160_;
	assign _1163_ = _1161_ & ~_1162_;
	assign _1164_ = (_1026_ ? _1161_ : _1163_);
	assign _1165_ = _1164_ | _1153_;
	assign _1166_ = _1165_ | ~_1159_;
	assign _1167_ = ~(_1166_ | _1141_);
	assign _1168_ = \mchip.DUT.freq_in [0] & ~_1167_;
	assign _0125_ = _1168_ | _1158_;
	assign _1169_ = ~_1153_;
	assign _1170_ = ~_1026_;
	assign _1171_ = _1147_ | ~_1144_;
	assign _1172_ = _1171_ | _1025_;
	assign _1173_ = _1172_ | _1170_;
	assign _1174_ = _1173_ | _1169_;
	assign _1175_ = _1156_ & ~_1174_;
	assign _1176_ = (\mchip.DUT.c [0] ? _1145_ : _1150_);
	assign _1177_ = _1176_ | _1026_;
	assign _1178_ = _1177_ | _1153_;
	assign _1179_ = _1159_ & ~_1178_;
	assign _1180_ = (_1141_ ? _1175_ : _1179_);
	assign _1181_ = _1084_ | _1170_;
	assign _1182_ = _1153_ & ~_1181_;
	assign _1183_ = _1163_ | _1026_;
	assign _1184_ = _1183_ | _1153_;
	assign _1185_ = (_1141_ ? _1182_ : _1184_);
	assign _1186_ = _1159_ & ~_1185_;
	assign _1187_ = \mchip.DUT.freq_in [1] & ~_1186_;
	assign _0126_ = _1187_ | _1180_;
	assign _1188_ = _1149_ | ~_1144_;
	assign _1189_ = (\mchip.DUT.c [0] ? _1188_ : _1171_);
	assign _1190_ = _1189_ | _1170_;
	assign _1191_ = _1190_ | _1169_;
	assign _1192_ = _1156_ & ~_1191_;
	assign _1193_ = _1146_ | _1026_;
	assign _1194_ = _1193_ | _1153_;
	assign _1195_ = _1159_ & ~_1194_;
	assign _1196_ = (_1141_ ? _1192_ : _1195_);
	assign _1197_ = _1143_ | _1031_;
	assign _1198_ = (\mchip.DUT.c [0] ? _1031_ : _1197_);
	assign _1199_ = _1198_ | ~_1026_;
	assign _1200_ = _1199_ | ~_1153_;
	assign _1201_ = ~(_1200_ | _1159_);
	assign _1202_ = _1161_ | _1026_;
	assign _1203_ = _1202_ | _1153_;
	assign _1204_ = _1159_ & ~_1203_;
	assign _1205_ = (_1141_ ? _1201_ : _1204_);
	assign _1206_ = \mchip.DUT.freq_in [2] & ~_1205_;
	assign _0127_ = _1206_ | _1196_;
	assign _1207_ = _1142_ | ~_1144_;
	assign _1208_ = (\mchip.DUT.c [0] ? _1207_ : _1188_);
	assign _1209_ = (_1026_ ? _1208_ : _1172_);
	assign _1210_ = _1209_ | _1169_;
	assign _1211_ = _1210_ | _1159_;
	assign _1212_ = _1141_ & ~_1211_;
	assign _1213_ = _0748_ & ~_1025_;
	assign _1214_ = ~(_1213_ & _1156_);
	assign _1215_ = _1141_ & ~_1214_;
	assign _1216_ = \mchip.DUT.freq_in [3] & ~_1215_;
	assign _0128_ = _1216_ | _1212_;
	assign _1217_ = _1207_ | \mchip.DUT.c [0];
	assign _1218_ = (_1026_ ? _1217_ : _1189_);
	assign _1219_ = _1218_ | _1169_;
	assign _1220_ = _1219_ | _1159_;
	assign _1221_ = _1141_ & ~_1220_;
	assign _1222_ = _1197_ | \mchip.DUT.c [0];
	assign _1223_ = (_1026_ ? _1222_ : _1198_);
	assign _1224_ = _1223_ | ~_1153_;
	assign _1225_ = _1224_ | _1159_;
	assign _1226_ = _1141_ & ~_1225_;
	assign _1227_ = \mchip.DUT.freq_in [4] & ~_1226_;
	assign _0129_ = _1227_ | _1221_;
	assign _1228_ = _1208_ | _1026_;
	assign _1229_ = (_1153_ ? _1228_ : _1173_);
	assign _1230_ = _1229_ | _1159_;
	assign _1231_ = _1141_ & ~_1230_;
	assign _1232_ = _1198_ | _1026_;
	assign _1233_ = (_1153_ ? _1232_ : _1181_);
	assign _1234_ = _1233_ | _1159_;
	assign _1235_ = _1141_ & ~_1234_;
	assign _1236_ = \mchip.DUT.freq_in [5] & ~_1235_;
	assign _0130_ = _1236_ | _1231_;
	assign _1237_ = _1217_ | _1026_;
	assign _1238_ = (_1153_ ? _1237_ : _1190_);
	assign _1239_ = _1238_ | _1159_;
	assign _1240_ = _1141_ & ~_1239_;
	assign _1241_ = _1222_ | _1026_;
	assign _1242_ = (_1153_ ? _1241_ : _1199_);
	assign _1243_ = _1242_ | _1159_;
	assign _1244_ = _1141_ & ~_1243_;
	assign _1245_ = \mchip.DUT.freq_in [6] & ~_1244_;
	assign _0131_ = _1245_ | _1240_;
	assign _1246_ = _1209_ | _1153_;
	assign _1247_ = _1246_ | _1159_;
	assign _1248_ = _1141_ & ~_1247_;
	assign _1249_ = (_1026_ ? _1198_ : _1084_);
	assign _1250_ = _1249_ | _1153_;
	assign _1251_ = _1250_ | _1159_;
	assign _1252_ = _1141_ & ~_1251_;
	assign _1253_ = \mchip.DUT.freq_in [7] & ~_1252_;
	assign _0132_ = _1253_ | _1248_;
	assign _1254_ = _1218_ | _1153_;
	assign _1255_ = _1254_ | _1159_;
	assign _1256_ = _1141_ & ~_1255_;
	assign _1257_ = _1223_ | _1153_;
	assign _1258_ = _1257_ | _1159_;
	assign _1259_ = _1141_ & ~_1258_;
	assign _1260_ = \mchip.DUT.freq_in [8] & ~_1259_;
	assign _0133_ = _1260_ | _1256_;
	assign _0002_ = \mchip.DUT.state [4] & ~io_in[13];
	assign _1261_ = ~\mchip.DUT.huff_tree[3] [1];
	assign _1262_ = _1723_ | _1261_;
	assign _1263_ = _1715_ | _1261_;
	assign _1264_ = \mchip.DUT.huff_tree[2] [1] & ~_1716_;
	assign _1265_ = _1263_ & ~_1264_;
	assign _1266_ = _1717_ & ~_1265_;
	assign _1767_[1] = _1266_ ^ _1722_;
	assign _1267_ = _1767_[1] & _1724_;
	assign _1268_ = _1262_ & ~_1267_;
	assign _1269_ = _1725_ & ~_1268_;
	assign _1769_[1] = ~(_1269_ ^ _1768_[0]);
	assign _1270_ = _1729_ | ~_1769_[1];
	assign _1271_ = _1767_[1] & _1730_;
	assign _1272_ = _1270_ & ~_1271_;
	assign _1273_ = _1731_ & ~_1272_;
	assign _1773_[1] = _1273_ ^ _1735_;
	assign _1274_ = _1736_ | ~_1769_[1];
	assign _1275_ = _1767_[1] & _1737_;
	assign _1276_ = _1274_ & ~_1275_;
	assign _1277_ = _1738_ & ~_1276_;
	assign _1771_[1] = _1277_ ^ _1742_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[4] [4] <= 1'h0;
		else if (_0007_)
			\mchip.DUT.huff_tree[4] [4] <= \mchip.DUT.node_sorter_ins.output_node [38];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[4] [5] <= 1'h0;
		else if (_0007_)
			\mchip.DUT.huff_tree[4] [5] <= \mchip.DUT.node_sorter_ins.output_node [39];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[4] [6] <= 1'h0;
		else if (_0007_)
			\mchip.DUT.huff_tree[4] [6] <= \mchip.DUT.node_sorter_ins.output_node [40];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[4] [7] <= 1'h0;
		else if (_0007_)
			\mchip.DUT.huff_tree[4] [7] <= \mchip.DUT.node_sorter_ins.output_node [41];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[4] [8] <= 1'h0;
		else if (_0007_)
			\mchip.DUT.huff_tree[4] [8] <= \mchip.DUT.node_sorter_ins.output_node [42];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[4] [9] <= 1'h0;
		else if (_0007_)
			\mchip.DUT.huff_tree[4] [9] <= \mchip.DUT.node_sorter_ins.output_node [43];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[4] [10] <= 1'h0;
		else if (_0007_)
			\mchip.DUT.huff_tree[4] [10] <= \mchip.DUT.node_sorter_ins.output_node [44];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[4] [11] <= 1'h0;
		else if (_0007_)
			\mchip.DUT.huff_tree[4] [11] <= \mchip.DUT.node_sorter_ins.output_node [45];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[4] [12] <= 1'h0;
		else if (_0007_)
			\mchip.DUT.huff_tree[4] [12] <= \mchip.DUT.node_sorter_ins.output_node [46];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[4] [13] <= 1'h0;
		else if (_0007_)
			\mchip.DUT.huff_tree[4] [13] <= \mchip.DUT.node_sorter_ins.output_node [47];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[4] [14] <= 1'h0;
		else if (_0007_)
			\mchip.DUT.huff_tree[4] [14] <= \mchip.DUT.node_sorter_ins.output_node [48];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[4] [15] <= 1'h0;
		else if (_0007_)
			\mchip.DUT.huff_tree[4] [15] <= \mchip.DUT.node_sorter_ins.output_node [52];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[4] [16] <= 1'h0;
		else if (_0007_)
			\mchip.DUT.huff_tree[4] [16] <= \mchip.DUT.node_sorter_ins.output_node [53];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[4] [17] <= 1'h0;
		else if (_0007_)
			\mchip.DUT.huff_tree[4] [17] <= \mchip.DUT.node_sorter_ins.output_node [54];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[4] [18] <= 1'h0;
		else if (_0007_)
			\mchip.DUT.huff_tree[4] [18] <= \mchip.DUT.node_sorter_ins.output_node [55];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[4] [19] <= 1'h0;
		else if (_0007_)
			\mchip.DUT.huff_tree[4] [19] <= \mchip.DUT.node_sorter_ins.output_node [56];
	always @(posedge io_in[12]) \mchip.DUT.state [0] <= _0004_;
	always @(posedge io_in[12]) \mchip.DUT.state [1] <= _0000_;
	always @(posedge io_in[12]) \mchip.DUT.state [2] <= _0001_;
	always @(posedge io_in[12]) \mchip.DUT.state [3] <= _0002_;
	always @(posedge io_in[12]) \mchip.DUT.state [4] <= _0003_;
	always @(posedge io_in[12]) \mchip.DUT.state [5] <= _0005_;
	always @(posedge io_in[12]) \mchip.DUT.state [6] <= _0006_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[5] [0] <= 1'h0;
		else if (\mchip.DUT.state [4])
			\mchip.DUT.huff_tree[5] [0] <= _1772_[0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[5] [1] <= 1'h0;
		else if (\mchip.DUT.state [4])
			\mchip.DUT.huff_tree[5] [1] <= _1773_[1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[5] [2] <= 1'h0;
		else if (\mchip.DUT.state [4])
			\mchip.DUT.huff_tree[5] [2] <= _0020_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[5] [3] <= 1'h0;
		else if (\mchip.DUT.state [4])
			\mchip.DUT.huff_tree[5] [3] <= _0041_;
	reg \mchip.DUT.in_huff_tree_reg[10] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.in_huff_tree_reg[10]  <= 1'h0;
		else if (!_0198_)
			\mchip.DUT.in_huff_tree_reg[10]  <= 1'h1;
	assign \mchip.DUT.in_huff_tree [10] = \mchip.DUT.in_huff_tree_reg[10] ;
	reg \mchip.DUT.in_huff_tree_reg[11] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.in_huff_tree_reg[11]  <= 1'h0;
		else if (!_0198_)
			\mchip.DUT.in_huff_tree_reg[11]  <= \mchip.DUT.freq_in [0];
	assign \mchip.DUT.in_huff_tree [11] = \mchip.DUT.in_huff_tree_reg[11] ;
	reg \mchip.DUT.in_huff_tree_reg[12] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.in_huff_tree_reg[12]  <= 1'h0;
		else if (!_0198_)
			\mchip.DUT.in_huff_tree_reg[12]  <= \mchip.DUT.freq_in [1];
	assign \mchip.DUT.in_huff_tree [12] = \mchip.DUT.in_huff_tree_reg[12] ;
	reg \mchip.DUT.in_huff_tree_reg[13] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.in_huff_tree_reg[13]  <= 1'h0;
		else if (!_0198_)
			\mchip.DUT.in_huff_tree_reg[13]  <= \mchip.DUT.freq_in [2];
	assign \mchip.DUT.in_huff_tree [13] = \mchip.DUT.in_huff_tree_reg[13] ;
	reg \mchip.DUT.in_huff_tree_reg[14] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.in_huff_tree_reg[14]  <= 1'h0;
		else if (!_0198_)
			\mchip.DUT.in_huff_tree_reg[14]  <= \mchip.DUT.data_in [0];
	assign \mchip.DUT.in_huff_tree [14] = \mchip.DUT.in_huff_tree_reg[14] ;
	reg \mchip.DUT.in_huff_tree_reg[15] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.in_huff_tree_reg[15]  <= 1'h0;
		else if (!_0198_)
			\mchip.DUT.in_huff_tree_reg[15]  <= \mchip.DUT.data_in [1];
	assign \mchip.DUT.in_huff_tree [15] = \mchip.DUT.in_huff_tree_reg[15] ;
	reg \mchip.DUT.in_huff_tree_reg[16] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.in_huff_tree_reg[16]  <= 1'h0;
		else if (!_0198_)
			\mchip.DUT.in_huff_tree_reg[16]  <= \mchip.DUT.data_in [2];
	assign \mchip.DUT.in_huff_tree [16] = \mchip.DUT.in_huff_tree_reg[16] ;
	reg \mchip.DUT.in_huff_tree_reg[17] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.in_huff_tree_reg[17]  <= 1'h0;
		else if (!_0198_)
			\mchip.DUT.in_huff_tree_reg[17]  <= \mchip.DUT.data_in [3];
	assign \mchip.DUT.in_huff_tree [17] = \mchip.DUT.in_huff_tree_reg[17] ;
	reg \mchip.DUT.in_huff_tree_reg[18] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.in_huff_tree_reg[18]  <= 1'h0;
		else if (!_0198_)
			\mchip.DUT.in_huff_tree_reg[18]  <= \mchip.DUT.data_in [4];
	assign \mchip.DUT.in_huff_tree [18] = \mchip.DUT.in_huff_tree_reg[18] ;
	reg \mchip.DUT.in_huff_tree_reg[19] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.in_huff_tree_reg[19]  <= 1'h0;
		else if (!_0198_)
			\mchip.DUT.in_huff_tree_reg[19]  <= _0053_;
	assign \mchip.DUT.in_huff_tree [19] = \mchip.DUT.in_huff_tree_reg[19] ;
	reg \mchip.DUT.in_huff_tree_reg[20] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.in_huff_tree_reg[20]  <= 1'h0;
		else if (!_0198_)
			\mchip.DUT.in_huff_tree_reg[20]  <= _0054_;
	assign \mchip.DUT.in_huff_tree [20] = \mchip.DUT.in_huff_tree_reg[20] ;
	reg \mchip.DUT.in_huff_tree_reg[21] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.in_huff_tree_reg[21]  <= 1'h0;
		else if (!_0198_)
			\mchip.DUT.in_huff_tree_reg[21]  <= _0055_;
	assign \mchip.DUT.in_huff_tree [21] = \mchip.DUT.in_huff_tree_reg[21] ;
	reg \mchip.DUT.in_huff_tree_reg[22] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.in_huff_tree_reg[22]  <= 1'h0;
		else if (!_0198_)
			\mchip.DUT.in_huff_tree_reg[22]  <= _0056_;
	assign \mchip.DUT.in_huff_tree [22] = \mchip.DUT.in_huff_tree_reg[22] ;
	reg \mchip.DUT.in_huff_tree_reg[23] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.in_huff_tree_reg[23]  <= 1'h0;
		else if (!_0198_)
			\mchip.DUT.in_huff_tree_reg[23]  <= _0057_;
	assign \mchip.DUT.in_huff_tree [23] = \mchip.DUT.in_huff_tree_reg[23] ;
	reg \mchip.DUT.in_huff_tree_reg[24] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.in_huff_tree_reg[24]  <= 1'h0;
		else if (!_0198_)
			\mchip.DUT.in_huff_tree_reg[24]  <= _0058_;
	assign \mchip.DUT.in_huff_tree [24] = \mchip.DUT.in_huff_tree_reg[24] ;
	reg \mchip.DUT.in_huff_tree_reg[25] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.in_huff_tree_reg[25]  <= 1'h0;
		else if (!_0198_)
			\mchip.DUT.in_huff_tree_reg[25]  <= _0059_;
	assign \mchip.DUT.in_huff_tree [25] = \mchip.DUT.in_huff_tree_reg[25] ;
	reg \mchip.DUT.in_huff_tree_reg[26] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.in_huff_tree_reg[26]  <= 1'h0;
		else if (!_0198_)
			\mchip.DUT.in_huff_tree_reg[26]  <= _0060_;
	assign \mchip.DUT.in_huff_tree [26] = \mchip.DUT.in_huff_tree_reg[26] ;
	reg \mchip.DUT.in_huff_tree_reg[27] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.in_huff_tree_reg[27]  <= 1'h0;
		else if (!_0198_)
			\mchip.DUT.in_huff_tree_reg[27]  <= _0061_;
	assign \mchip.DUT.in_huff_tree [27] = \mchip.DUT.in_huff_tree_reg[27] ;
	reg \mchip.DUT.in_huff_tree_reg[28] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.in_huff_tree_reg[28]  <= 1'h0;
		else if (!_0198_)
			\mchip.DUT.in_huff_tree_reg[28]  <= _0062_;
	assign \mchip.DUT.in_huff_tree [28] = \mchip.DUT.in_huff_tree_reg[28] ;
	reg \mchip.DUT.in_huff_tree_reg[29] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.in_huff_tree_reg[29]  <= 1'h0;
		else if (!_0198_)
			\mchip.DUT.in_huff_tree_reg[29]  <= _0063_;
	assign \mchip.DUT.in_huff_tree [29] = \mchip.DUT.in_huff_tree_reg[29] ;
	reg \mchip.DUT.in_huff_tree_reg[30] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.in_huff_tree_reg[30]  <= 1'h0;
		else if (!_0198_)
			\mchip.DUT.in_huff_tree_reg[30]  <= _0064_;
	assign \mchip.DUT.in_huff_tree [30] = \mchip.DUT.in_huff_tree_reg[30] ;
	reg \mchip.DUT.in_huff_tree_reg[31] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.in_huff_tree_reg[31]  <= 1'h0;
		else if (!_0198_)
			\mchip.DUT.in_huff_tree_reg[31]  <= _0065_;
	assign \mchip.DUT.in_huff_tree [31] = \mchip.DUT.in_huff_tree_reg[31] ;
	reg \mchip.DUT.in_huff_tree_reg[32] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.in_huff_tree_reg[32]  <= 1'h0;
		else if (!_0198_)
			\mchip.DUT.in_huff_tree_reg[32]  <= _0066_;
	assign \mchip.DUT.in_huff_tree [32] = \mchip.DUT.in_huff_tree_reg[32] ;
	reg \mchip.DUT.in_huff_tree_reg[33] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.in_huff_tree_reg[33]  <= 1'h0;
		else if (!_0198_)
			\mchip.DUT.in_huff_tree_reg[33]  <= _0067_;
	assign \mchip.DUT.in_huff_tree [33] = \mchip.DUT.in_huff_tree_reg[33] ;
	reg \mchip.DUT.in_huff_tree_reg[34] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.in_huff_tree_reg[34]  <= 1'h0;
		else if (!_0198_)
			\mchip.DUT.in_huff_tree_reg[34]  <= _0068_;
	assign \mchip.DUT.in_huff_tree [34] = \mchip.DUT.in_huff_tree_reg[34] ;
	reg \mchip.DUT.in_huff_tree_reg[35] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.in_huff_tree_reg[35]  <= 1'h0;
		else if (!_0198_)
			\mchip.DUT.in_huff_tree_reg[35]  <= _0069_;
	assign \mchip.DUT.in_huff_tree [35] = \mchip.DUT.in_huff_tree_reg[35] ;
	reg \mchip.DUT.in_huff_tree_reg[36] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.in_huff_tree_reg[36]  <= 1'h0;
		else if (!_0198_)
			\mchip.DUT.in_huff_tree_reg[36]  <= _0070_;
	assign \mchip.DUT.in_huff_tree [36] = \mchip.DUT.in_huff_tree_reg[36] ;
	reg \mchip.DUT.in_huff_tree_reg[37] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.in_huff_tree_reg[37]  <= 1'h0;
		else if (!_0198_)
			\mchip.DUT.in_huff_tree_reg[37]  <= _0071_;
	assign \mchip.DUT.in_huff_tree [37] = \mchip.DUT.in_huff_tree_reg[37] ;
	reg \mchip.DUT.in_huff_tree_reg[38] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.in_huff_tree_reg[38]  <= 1'h0;
		else if (!_0198_)
			\mchip.DUT.in_huff_tree_reg[38]  <= _0072_;
	assign \mchip.DUT.in_huff_tree [38] = \mchip.DUT.in_huff_tree_reg[38] ;
	reg \mchip.DUT.in_huff_tree_reg[39] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.in_huff_tree_reg[39]  <= 1'h0;
		else if (!_0198_)
			\mchip.DUT.in_huff_tree_reg[39]  <= _0073_;
	assign \mchip.DUT.in_huff_tree [39] = \mchip.DUT.in_huff_tree_reg[39] ;
	reg \mchip.DUT.in_huff_tree_reg[40] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.in_huff_tree_reg[40]  <= 1'h0;
		else if (!_0198_)
			\mchip.DUT.in_huff_tree_reg[40]  <= _0074_;
	assign \mchip.DUT.in_huff_tree [40] = \mchip.DUT.in_huff_tree_reg[40] ;
	reg \mchip.DUT.in_huff_tree_reg[41] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.in_huff_tree_reg[41]  <= 1'h0;
		else if (!_0198_)
			\mchip.DUT.in_huff_tree_reg[41]  <= _0075_;
	assign \mchip.DUT.in_huff_tree [41] = \mchip.DUT.in_huff_tree_reg[41] ;
	reg \mchip.DUT.in_huff_tree_reg[42] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.in_huff_tree_reg[42]  <= 1'h0;
		else if (!_0198_)
			\mchip.DUT.in_huff_tree_reg[42]  <= _0076_;
	assign \mchip.DUT.in_huff_tree [42] = \mchip.DUT.in_huff_tree_reg[42] ;
	reg \mchip.DUT.in_huff_tree_reg[43] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.in_huff_tree_reg[43]  <= 1'h0;
		else if (!_0198_)
			\mchip.DUT.in_huff_tree_reg[43]  <= _0077_;
	assign \mchip.DUT.in_huff_tree [43] = \mchip.DUT.in_huff_tree_reg[43] ;
	reg \mchip.DUT.in_huff_tree_reg[44] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.in_huff_tree_reg[44]  <= 1'h0;
		else if (!_0198_)
			\mchip.DUT.in_huff_tree_reg[44]  <= _0078_;
	assign \mchip.DUT.in_huff_tree [44] = \mchip.DUT.in_huff_tree_reg[44] ;
	reg \mchip.DUT.in_huff_tree_reg[45] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.in_huff_tree_reg[45]  <= 1'h0;
		else if (!_0198_)
			\mchip.DUT.in_huff_tree_reg[45]  <= _0079_;
	assign \mchip.DUT.in_huff_tree [45] = \mchip.DUT.in_huff_tree_reg[45] ;
	reg \mchip.DUT.in_huff_tree_reg[46] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.in_huff_tree_reg[46]  <= 1'h0;
		else if (!_0198_)
			\mchip.DUT.in_huff_tree_reg[46]  <= _0080_;
	assign \mchip.DUT.in_huff_tree [46] = \mchip.DUT.in_huff_tree_reg[46] ;
	reg \mchip.DUT.in_huff_tree_reg[47] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.in_huff_tree_reg[47]  <= 1'h0;
		else if (!_0198_)
			\mchip.DUT.in_huff_tree_reg[47]  <= _0081_;
	assign \mchip.DUT.in_huff_tree [47] = \mchip.DUT.in_huff_tree_reg[47] ;
	reg \mchip.DUT.in_huff_tree_reg[48] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.in_huff_tree_reg[48]  <= 1'h0;
		else if (!_0198_)
			\mchip.DUT.in_huff_tree_reg[48]  <= _0082_;
	assign \mchip.DUT.in_huff_tree [48] = \mchip.DUT.in_huff_tree_reg[48] ;
	reg \mchip.DUT.in_huff_tree_reg[49] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.in_huff_tree_reg[49]  <= 1'h0;
		else if (!_0198_)
			\mchip.DUT.in_huff_tree_reg[49]  <= _0083_;
	assign \mchip.DUT.in_huff_tree [49] = \mchip.DUT.in_huff_tree_reg[49] ;
	reg \mchip.DUT.in_huff_tree_reg[50] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.in_huff_tree_reg[50]  <= 1'h0;
		else if (!_0198_)
			\mchip.DUT.in_huff_tree_reg[50]  <= _0084_;
	assign \mchip.DUT.in_huff_tree [50] = \mchip.DUT.in_huff_tree_reg[50] ;
	reg \mchip.DUT.in_huff_tree_reg[51] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.in_huff_tree_reg[51]  <= 1'h0;
		else if (!_0198_)
			\mchip.DUT.in_huff_tree_reg[51]  <= _0085_;
	assign \mchip.DUT.in_huff_tree [51] = \mchip.DUT.in_huff_tree_reg[51] ;
	reg \mchip.DUT.in_huff_tree_reg[52] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.in_huff_tree_reg[52]  <= 1'h0;
		else if (!_0198_)
			\mchip.DUT.in_huff_tree_reg[52]  <= _0086_;
	assign \mchip.DUT.in_huff_tree [52] = \mchip.DUT.in_huff_tree_reg[52] ;
	reg \mchip.DUT.in_huff_tree_reg[53] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.in_huff_tree_reg[53]  <= 1'h0;
		else if (!_0198_)
			\mchip.DUT.in_huff_tree_reg[53]  <= _0087_;
	assign \mchip.DUT.in_huff_tree [53] = \mchip.DUT.in_huff_tree_reg[53] ;
	reg \mchip.DUT.in_huff_tree_reg[54] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.in_huff_tree_reg[54]  <= 1'h0;
		else if (!_0198_)
			\mchip.DUT.in_huff_tree_reg[54]  <= _0088_;
	assign \mchip.DUT.in_huff_tree [54] = \mchip.DUT.in_huff_tree_reg[54] ;
	reg \mchip.DUT.in_huff_tree_reg[55] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.in_huff_tree_reg[55]  <= 1'h0;
		else if (!_0198_)
			\mchip.DUT.in_huff_tree_reg[55]  <= _0089_;
	assign \mchip.DUT.in_huff_tree [55] = \mchip.DUT.in_huff_tree_reg[55] ;
	reg \mchip.DUT.in_huff_tree_reg[56] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.in_huff_tree_reg[56]  <= 1'h0;
		else if (!_0198_)
			\mchip.DUT.in_huff_tree_reg[56]  <= _0090_;
	assign \mchip.DUT.in_huff_tree [56] = \mchip.DUT.in_huff_tree_reg[56] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[3] [0] <= 1'h0;
		else if (\mchip.DUT.state [4])
			\mchip.DUT.huff_tree[3] [0] <= _1768_[0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[3] [1] <= 1'h0;
		else if (\mchip.DUT.state [4])
			\mchip.DUT.huff_tree[3] [1] <= _1769_[1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[3] [2] <= 1'h0;
		else if (\mchip.DUT.state [4])
			\mchip.DUT.huff_tree[3] [2] <= _0018_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[3] [3] <= 1'h0;
		else if (\mchip.DUT.state [4])
			\mchip.DUT.huff_tree[3] [3] <= _0039_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[2] [4] <= 1'h0;
		else if (_0008_)
			\mchip.DUT.huff_tree[2] [4] <= \mchip.DUT.node_sorter_ins.output_node [38];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[2] [5] <= 1'h0;
		else if (_0008_)
			\mchip.DUT.huff_tree[2] [5] <= \mchip.DUT.node_sorter_ins.output_node [39];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[2] [6] <= 1'h0;
		else if (_0008_)
			\mchip.DUT.huff_tree[2] [6] <= \mchip.DUT.node_sorter_ins.output_node [40];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[2] [7] <= 1'h0;
		else if (_0008_)
			\mchip.DUT.huff_tree[2] [7] <= \mchip.DUT.node_sorter_ins.output_node [41];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[2] [8] <= 1'h0;
		else if (_0008_)
			\mchip.DUT.huff_tree[2] [8] <= \mchip.DUT.node_sorter_ins.output_node [42];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[2] [9] <= 1'h0;
		else if (_0008_)
			\mchip.DUT.huff_tree[2] [9] <= \mchip.DUT.node_sorter_ins.output_node [43];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[2] [10] <= 1'h0;
		else if (_0008_)
			\mchip.DUT.huff_tree[2] [10] <= \mchip.DUT.node_sorter_ins.output_node [44];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[2] [11] <= 1'h0;
		else if (_0008_)
			\mchip.DUT.huff_tree[2] [11] <= \mchip.DUT.node_sorter_ins.output_node [45];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[2] [12] <= 1'h0;
		else if (_0008_)
			\mchip.DUT.huff_tree[2] [12] <= \mchip.DUT.node_sorter_ins.output_node [46];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[2] [13] <= 1'h0;
		else if (_0008_)
			\mchip.DUT.huff_tree[2] [13] <= \mchip.DUT.node_sorter_ins.output_node [47];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[2] [14] <= 1'h0;
		else if (_0008_)
			\mchip.DUT.huff_tree[2] [14] <= \mchip.DUT.node_sorter_ins.output_node [48];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[2] [15] <= 1'h0;
		else if (_0008_)
			\mchip.DUT.huff_tree[2] [15] <= \mchip.DUT.node_sorter_ins.output_node [52];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[2] [16] <= 1'h0;
		else if (_0008_)
			\mchip.DUT.huff_tree[2] [16] <= \mchip.DUT.node_sorter_ins.output_node [53];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[2] [17] <= 1'h0;
		else if (_0008_)
			\mchip.DUT.huff_tree[2] [17] <= \mchip.DUT.node_sorter_ins.output_node [54];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[2] [18] <= 1'h0;
		else if (_0008_)
			\mchip.DUT.huff_tree[2] [18] <= \mchip.DUT.node_sorter_ins.output_node [55];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[2] [19] <= 1'h0;
		else if (_0008_)
			\mchip.DUT.huff_tree[2] [19] <= \mchip.DUT.node_sorter_ins.output_node [56];
	reg \mchip.DUT.huff_tree_reg[1][4] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree_reg[1][4]  <= 1'h0;
		else if (\mchip.DUT.state [1])
			\mchip.DUT.huff_tree_reg[1][4]  <= \mchip.DUT.node_sorter_ins.output_node [38];
	assign \mchip.DUT.huff_tree[1] [4] = \mchip.DUT.huff_tree_reg[1][4] ;
	reg \mchip.DUT.huff_tree_reg[1][5] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree_reg[1][5]  <= 1'h0;
		else if (\mchip.DUT.state [1])
			\mchip.DUT.huff_tree_reg[1][5]  <= \mchip.DUT.node_sorter_ins.output_node [39];
	assign \mchip.DUT.huff_tree[1] [5] = \mchip.DUT.huff_tree_reg[1][5] ;
	reg \mchip.DUT.huff_tree_reg[1][6] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree_reg[1][6]  <= 1'h0;
		else if (\mchip.DUT.state [1])
			\mchip.DUT.huff_tree_reg[1][6]  <= \mchip.DUT.node_sorter_ins.output_node [40];
	assign \mchip.DUT.huff_tree[1] [6] = \mchip.DUT.huff_tree_reg[1][6] ;
	reg \mchip.DUT.huff_tree_reg[1][7] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree_reg[1][7]  <= 1'h0;
		else if (\mchip.DUT.state [1])
			\mchip.DUT.huff_tree_reg[1][7]  <= \mchip.DUT.node_sorter_ins.output_node [41];
	assign \mchip.DUT.huff_tree[1] [7] = \mchip.DUT.huff_tree_reg[1][7] ;
	reg \mchip.DUT.huff_tree_reg[1][8] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree_reg[1][8]  <= 1'h0;
		else if (\mchip.DUT.state [1])
			\mchip.DUT.huff_tree_reg[1][8]  <= \mchip.DUT.node_sorter_ins.output_node [42];
	assign \mchip.DUT.huff_tree[1] [8] = \mchip.DUT.huff_tree_reg[1][8] ;
	reg \mchip.DUT.huff_tree_reg[1][9] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree_reg[1][9]  <= 1'h0;
		else if (\mchip.DUT.state [1])
			\mchip.DUT.huff_tree_reg[1][9]  <= \mchip.DUT.node_sorter_ins.output_node [43];
	assign \mchip.DUT.huff_tree[1] [9] = \mchip.DUT.huff_tree_reg[1][9] ;
	reg \mchip.DUT.huff_tree_reg[1][10] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree_reg[1][10]  <= 1'h0;
		else if (\mchip.DUT.state [1])
			\mchip.DUT.huff_tree_reg[1][10]  <= \mchip.DUT.node_sorter_ins.output_node [44];
	assign \mchip.DUT.huff_tree[1] [10] = \mchip.DUT.huff_tree_reg[1][10] ;
	reg \mchip.DUT.huff_tree_reg[1][11] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree_reg[1][11]  <= 1'h0;
		else if (\mchip.DUT.state [1])
			\mchip.DUT.huff_tree_reg[1][11]  <= \mchip.DUT.node_sorter_ins.output_node [45];
	assign \mchip.DUT.huff_tree[1] [11] = \mchip.DUT.huff_tree_reg[1][11] ;
	reg \mchip.DUT.huff_tree_reg[1][12] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree_reg[1][12]  <= 1'h0;
		else if (\mchip.DUT.state [1])
			\mchip.DUT.huff_tree_reg[1][12]  <= \mchip.DUT.node_sorter_ins.output_node [46];
	assign \mchip.DUT.huff_tree[1] [12] = \mchip.DUT.huff_tree_reg[1][12] ;
	reg \mchip.DUT.huff_tree_reg[1][13] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree_reg[1][13]  <= 1'h0;
		else if (\mchip.DUT.state [1])
			\mchip.DUT.huff_tree_reg[1][13]  <= \mchip.DUT.node_sorter_ins.output_node [47];
	assign \mchip.DUT.huff_tree[1] [13] = \mchip.DUT.huff_tree_reg[1][13] ;
	reg \mchip.DUT.huff_tree_reg[1][14] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree_reg[1][14]  <= 1'h0;
		else if (\mchip.DUT.state [1])
			\mchip.DUT.huff_tree_reg[1][14]  <= \mchip.DUT.node_sorter_ins.output_node [48];
	assign \mchip.DUT.huff_tree[1] [14] = \mchip.DUT.huff_tree_reg[1][14] ;
	reg \mchip.DUT.huff_tree_reg[1][15] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree_reg[1][15]  <= 1'h0;
		else if (\mchip.DUT.state [1])
			\mchip.DUT.huff_tree_reg[1][15]  <= \mchip.DUT.node_sorter_ins.output_node [52];
	assign \mchip.DUT.huff_tree[1] [15] = \mchip.DUT.huff_tree_reg[1][15] ;
	reg \mchip.DUT.huff_tree_reg[1][16] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree_reg[1][16]  <= 1'h0;
		else if (\mchip.DUT.state [1])
			\mchip.DUT.huff_tree_reg[1][16]  <= \mchip.DUT.node_sorter_ins.output_node [53];
	assign \mchip.DUT.huff_tree[1] [16] = \mchip.DUT.huff_tree_reg[1][16] ;
	reg \mchip.DUT.huff_tree_reg[1][17] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree_reg[1][17]  <= 1'h0;
		else if (\mchip.DUT.state [1])
			\mchip.DUT.huff_tree_reg[1][17]  <= \mchip.DUT.node_sorter_ins.output_node [54];
	assign \mchip.DUT.huff_tree[1] [17] = \mchip.DUT.huff_tree_reg[1][17] ;
	reg \mchip.DUT.huff_tree_reg[1][18] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree_reg[1][18]  <= 1'h0;
		else if (\mchip.DUT.state [1])
			\mchip.DUT.huff_tree_reg[1][18]  <= \mchip.DUT.node_sorter_ins.output_node [55];
	assign \mchip.DUT.huff_tree[1] [18] = \mchip.DUT.huff_tree_reg[1][18] ;
	reg \mchip.DUT.huff_tree_reg[1][19] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree_reg[1][19]  <= 1'h0;
		else if (\mchip.DUT.state [1])
			\mchip.DUT.huff_tree_reg[1][19]  <= \mchip.DUT.node_sorter_ins.output_node [56];
	assign \mchip.DUT.huff_tree[1] [19] = \mchip.DUT.huff_tree_reg[1][19] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.character [5] <= 1'h0;
		else if (_0012_)
			\mchip.DUT.character [5] <= _0027_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.character [6] <= 1'h0;
		else if (_0012_)
			\mchip.DUT.character [6] <= _0028_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.character [7] <= 1'h0;
		else if (_0012_)
			\mchip.DUT.character [7] <= _0029_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.character [8] <= 1'h0;
		else if (_0012_)
			\mchip.DUT.character [8] <= _0030_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.character [9] <= 1'h0;
		else if (_0012_)
			\mchip.DUT.character [9] <= _0031_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.character [0] <= 1'h0;
		else if (_0013_)
			\mchip.DUT.character [0] <= _0042_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.character [1] <= 1'h0;
		else if (_0013_)
			\mchip.DUT.character [1] <= _0043_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.character [2] <= 1'h0;
		else if (_0013_)
			\mchip.DUT.character [2] <= _0044_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.character [3] <= 1'h0;
		else if (_0013_)
			\mchip.DUT.character [3] <= _0045_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.character [4] <= 1'h0;
		else if (_0013_)
			\mchip.DUT.character [4] <= _0046_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.encoded_mask [3] <= 1'h0;
		else if (_0012_)
			\mchip.DUT.encoded_mask [3] <= _0032_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.encoded_mask [4] <= 1'h0;
		else if (_0012_)
			\mchip.DUT.encoded_mask [4] <= _0033_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.encoded_mask [5] <= 1'h0;
		else if (_0012_)
			\mchip.DUT.encoded_mask [5] <= _0034_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.encoded_mask [0] <= 1'h0;
		else if (_0013_)
			\mchip.DUT.encoded_mask [0] <= _0047_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.encoded_mask [1] <= 1'h0;
		else if (_0013_)
			\mchip.DUT.encoded_mask [1] <= _0048_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.encoded_mask [2] <= 1'h0;
		else if (_0013_)
			\mchip.DUT.encoded_mask [2] <= _0049_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.encoded_value [3] <= 1'h0;
		else if (_0012_)
			\mchip.DUT.encoded_value [3] <= _0035_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.encoded_value [4] <= 1'h0;
		else if (_0012_)
			\mchip.DUT.encoded_value [4] <= _0036_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.encoded_value [5] <= 1'h0;
		else if (_0012_)
			\mchip.DUT.encoded_value [5] <= _0037_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.encoded_value [0] <= 1'h0;
		else if (_0013_)
			\mchip.DUT.encoded_value [0] <= _0050_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.encoded_value [1] <= 1'h0;
		else if (_0013_)
			\mchip.DUT.encoded_value [1] <= _0051_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.encoded_value [2] <= 1'h0;
		else if (_0013_)
			\mchip.DUT.encoded_value [2] <= _0052_;
	always @(posedge io_in[12])
		if (_0014_)
			if (!\mchip.DUT.state [1])
				\mchip.DUT.count [0] <= 1'h1;
			else
				\mchip.DUT.count [0] <= _1775_[0];
	always @(posedge io_in[12])
		if (_0014_)
			if (!\mchip.DUT.state [1])
				\mchip.DUT.count [1] <= 1'h1;
			else
				\mchip.DUT.count [1] <= _1775_[1];
	reg \mchip.DUT.io_out_reg[0] ;
	always @(posedge io_in[12])
		if (_0016_)
			if (!\mchip.DUT.state [6])
				\mchip.DUT.io_out_reg[0]  <= 1'h0;
			else
				\mchip.DUT.io_out_reg[0]  <= _0021_;
	assign \mchip.DUT.io_out [0] = \mchip.DUT.io_out_reg[0] ;
	reg \mchip.DUT.io_out_reg[1] ;
	always @(posedge io_in[12])
		if (_0016_)
			if (!\mchip.DUT.state [6])
				\mchip.DUT.io_out_reg[1]  <= 1'h0;
			else
				\mchip.DUT.io_out_reg[1]  <= _0022_;
	assign \mchip.DUT.io_out [1] = \mchip.DUT.io_out_reg[1] ;
	reg \mchip.DUT.io_out_reg[2] ;
	always @(posedge io_in[12])
		if (_0016_)
			if (!\mchip.DUT.state [6])
				\mchip.DUT.io_out_reg[2]  <= 1'h0;
			else
				\mchip.DUT.io_out_reg[2]  <= _0023_;
	assign \mchip.DUT.io_out [2] = \mchip.DUT.io_out_reg[2] ;
	reg \mchip.DUT.io_out_reg[3] ;
	always @(posedge io_in[12])
		if (_0016_)
			if (!\mchip.DUT.state [6])
				\mchip.DUT.io_out_reg[3]  <= 1'h0;
			else
				\mchip.DUT.io_out_reg[3]  <= _0024_;
	assign \mchip.DUT.io_out [3] = \mchip.DUT.io_out_reg[3] ;
	reg \mchip.DUT.io_out_reg[4] ;
	always @(posedge io_in[12])
		if (_0016_)
			if (!\mchip.DUT.state [6])
				\mchip.DUT.io_out_reg[4]  <= 1'h0;
			else
				\mchip.DUT.io_out_reg[4]  <= _0025_;
	assign \mchip.DUT.io_out [4] = \mchip.DUT.io_out_reg[4] ;
	reg \mchip.DUT.io_out_reg[5] ;
	always @(posedge io_in[12])
		if (_0016_)
			if (!\mchip.DUT.state [6])
				\mchip.DUT.io_out_reg[5]  <= 1'h0;
			else
				\mchip.DUT.io_out_reg[5]  <= _0026_;
	assign \mchip.DUT.io_out [5] = \mchip.DUT.io_out_reg[5] ;
	reg \mchip.DUT.io_out_reg[6] ;
	always @(posedge io_in[12])
		if (_0016_)
			if (!\mchip.DUT.state [6])
				\mchip.DUT.io_out_reg[6]  <= 1'h0;
			else
				\mchip.DUT.io_out_reg[6]  <= _1774_[0];
	assign \mchip.DUT.io_out [6] = \mchip.DUT.io_out_reg[6] ;
	reg \mchip.DUT.data_in_reg[0] ;
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.DUT.data_in_reg[0]  <= _0110_;
	assign \mchip.DUT.data_in [0] = \mchip.DUT.data_in_reg[0] ;
	reg \mchip.DUT.data_in_reg[1] ;
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.DUT.data_in_reg[1]  <= _0118_;
	assign \mchip.DUT.data_in [1] = \mchip.DUT.data_in_reg[1] ;
	reg \mchip.DUT.data_in_reg[2] ;
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.DUT.data_in_reg[2]  <= _0120_;
	assign \mchip.DUT.data_in [2] = \mchip.DUT.data_in_reg[2] ;
	reg \mchip.DUT.data_in_reg[3] ;
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.DUT.data_in_reg[3]  <= _0121_;
	assign \mchip.DUT.data_in [3] = \mchip.DUT.data_in_reg[3] ;
	reg \mchip.DUT.data_in_reg[4] ;
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.DUT.data_in_reg[4]  <= _0122_;
	assign \mchip.DUT.data_in [4] = \mchip.DUT.data_in_reg[4] ;
	reg \mchip.DUT.data_in_reg[8] ;
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.DUT.data_in_reg[8]  <= _0123_;
	assign \mchip.DUT.data_in [8] = \mchip.DUT.data_in_reg[8] ;
	reg \mchip.DUT.data_in_reg[9] ;
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.DUT.data_in_reg[9]  <= _0124_;
	assign \mchip.DUT.data_in [9] = \mchip.DUT.data_in_reg[9] ;
	reg \mchip.DUT.data_in_reg[10] ;
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.DUT.data_in_reg[10]  <= _0111_;
	assign \mchip.DUT.data_in [10] = \mchip.DUT.data_in_reg[10] ;
	reg \mchip.DUT.data_in_reg[11] ;
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.DUT.data_in_reg[11]  <= _0112_;
	assign \mchip.DUT.data_in [11] = \mchip.DUT.data_in_reg[11] ;
	reg \mchip.DUT.data_in_reg[12] ;
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.DUT.data_in_reg[12]  <= _0113_;
	assign \mchip.DUT.data_in [12] = \mchip.DUT.data_in_reg[12] ;
	reg \mchip.DUT.data_in_reg[16] ;
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.DUT.data_in_reg[16]  <= _0114_;
	assign \mchip.DUT.data_in [16] = \mchip.DUT.data_in_reg[16] ;
	reg \mchip.DUT.data_in_reg[17] ;
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.DUT.data_in_reg[17]  <= _0115_;
	assign \mchip.DUT.data_in [17] = \mchip.DUT.data_in_reg[17] ;
	reg \mchip.DUT.data_in_reg[18] ;
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.DUT.data_in_reg[18]  <= _0116_;
	assign \mchip.DUT.data_in [18] = \mchip.DUT.data_in_reg[18] ;
	reg \mchip.DUT.data_in_reg[19] ;
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.DUT.data_in_reg[19]  <= _0117_;
	assign \mchip.DUT.data_in [19] = \mchip.DUT.data_in_reg[19] ;
	reg \mchip.DUT.data_in_reg[20] ;
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.DUT.data_in_reg[20]  <= _0119_;
	assign \mchip.DUT.data_in [20] = \mchip.DUT.data_in_reg[20] ;
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.DUT.freq_in [0] <= _0125_;
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.DUT.freq_in [1] <= _0126_;
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.DUT.freq_in [2] <= _0127_;
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.DUT.freq_in [3] <= _0128_;
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.DUT.freq_in [4] <= _0129_;
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.DUT.freq_in [5] <= _0130_;
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.DUT.freq_in [6] <= _0131_;
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.DUT.freq_in [7] <= _0132_;
	always @(posedge io_in[12])
		if (_0015_)
			\mchip.DUT.freq_in [8] <= _0133_;
	reg \mchip.DUT.io_out_reg[8] ;
	always @(posedge io_in[12])
		if (_0016_)
			\mchip.DUT.io_out_reg[8]  <= \mchip.DUT.state [6];
	assign \mchip.DUT.io_out [8] = \mchip.DUT.io_out_reg[8] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.encoded_value [6] <= 1'h0;
		else if (_0011_)
			\mchip.DUT.encoded_value [6] <= _0107_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.encoded_value [7] <= 1'h0;
		else if (_0011_)
			\mchip.DUT.encoded_value [7] <= _0108_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.encoded_value [8] <= 1'h0;
		else if (_0011_)
			\mchip.DUT.encoded_value [8] <= _0109_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.encoded_mask [6] <= 1'h0;
		else if (_0011_)
			\mchip.DUT.encoded_mask [6] <= _0104_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.encoded_mask [7] <= 1'h0;
		else if (_0011_)
			\mchip.DUT.encoded_mask [7] <= _0105_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.encoded_mask [8] <= 1'h0;
		else if (_0011_)
			\mchip.DUT.encoded_mask [8] <= _0106_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.character [10] <= 1'h0;
		else if (_0011_)
			\mchip.DUT.character [10] <= _0099_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.character [11] <= 1'h0;
		else if (_0011_)
			\mchip.DUT.character [11] <= _0100_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.character [12] <= 1'h0;
		else if (_0011_)
			\mchip.DUT.character [12] <= _0101_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.character [13] <= 1'h0;
		else if (_0011_)
			\mchip.DUT.character [13] <= _0102_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.character [14] <= 1'h0;
		else if (_0011_)
			\mchip.DUT.character [14] <= _0103_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.a [0] <= 1'h0;
		else if (_0010_)
			\mchip.DUT.a [0] <= _0138_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.a [1] <= 1'h0;
		else if (_0010_)
			\mchip.DUT.a [1] <= _0139_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.a [2] <= 1'h0;
		else if (_0010_)
			\mchip.DUT.a [2] <= _0140_;
	reg \mchip.DUT.b_reg[0] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.b_reg[0]  <= 1'h0;
		else if (!_0199_)
			\mchip.DUT.b_reg[0]  <= _0137_;
	assign \mchip.DUT.b [0] = \mchip.DUT.b_reg[0] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.c [0] <= 1'h0;
		else if (_0009_)
			\mchip.DUT.c [0] <= _0134_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.c [1] <= 1'h0;
		else if (_0009_)
			\mchip.DUT.c [1] <= _0135_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.c [2] <= 1'h0;
		else if (_0009_)
			\mchip.DUT.c [2] <= _0136_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.encoded_value_h[2] [0] <= 1'h0;
		else if (\mchip.DUT.state [3])
			\mchip.DUT.encoded_value_h[2] [0] <= _1776_[2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.encoded_value_h[2] [1] <= 1'h0;
		else if (\mchip.DUT.state [3])
			\mchip.DUT.encoded_value_h[2] [1] <= _1776_[3];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.encoded_value_h[2] [2] <= 1'h0;
		else if (\mchip.DUT.state [3])
			\mchip.DUT.encoded_value_h[2] [2] <= _0091_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.encoded_value_h[3] [0] <= 1'h0;
		else if (\mchip.DUT.state [3])
			\mchip.DUT.encoded_value_h[3] [0] <= _1776_[0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.encoded_value_h[3] [1] <= 1'h0;
		else if (\mchip.DUT.state [3])
			\mchip.DUT.encoded_value_h[3] [1] <= _1776_[1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.encoded_value_h[3] [2] <= 1'h0;
		else if (\mchip.DUT.state [3])
			\mchip.DUT.encoded_value_h[3] [2] <= _0092_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.encoded_value_h[4] [0] <= 1'h0;
		else if (\mchip.DUT.state [3])
			\mchip.DUT.encoded_value_h[4] [0] <= _0093_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.encoded_value_h[4] [1] <= 1'h0;
		else if (\mchip.DUT.state [3])
			\mchip.DUT.encoded_value_h[4] [1] <= _0094_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.encoded_value_h[4] [2] <= 1'h0;
		else if (\mchip.DUT.state [3])
			\mchip.DUT.encoded_value_h[4] [2] <= _0095_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.encoded_value_h[5] [0] <= 1'h0;
		else if (\mchip.DUT.state [3])
			\mchip.DUT.encoded_value_h[5] [0] <= _0096_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.encoded_value_h[5] [1] <= 1'h0;
		else if (\mchip.DUT.state [3])
			\mchip.DUT.encoded_value_h[5] [1] <= _0097_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.encoded_value_h[5] [2] <= 1'h0;
		else if (\mchip.DUT.state [3])
			\mchip.DUT.encoded_value_h[5] [2] <= _0098_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[2] [0] <= 1'h0;
		else if (\mchip.DUT.state [4])
			\mchip.DUT.huff_tree[2] [0] <= _1766_[0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[2] [1] <= 1'h0;
		else if (\mchip.DUT.state [4])
			\mchip.DUT.huff_tree[2] [1] <= _1767_[1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[2] [2] <= 1'h0;
		else if (\mchip.DUT.state [4])
			\mchip.DUT.huff_tree[2] [2] <= _0019_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[2] [3] <= 1'h0;
		else if (\mchip.DUT.state [4])
			\mchip.DUT.huff_tree[2] [3] <= _0038_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[3] [4] <= 1'h0;
		else if (_0008_)
			\mchip.DUT.huff_tree[3] [4] <= \mchip.DUT.node_sorter_ins.output_node [19];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[3] [5] <= 1'h0;
		else if (_0008_)
			\mchip.DUT.huff_tree[3] [5] <= \mchip.DUT.node_sorter_ins.output_node [20];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[3] [6] <= 1'h0;
		else if (_0008_)
			\mchip.DUT.huff_tree[3] [6] <= \mchip.DUT.node_sorter_ins.output_node [21];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[3] [7] <= 1'h0;
		else if (_0008_)
			\mchip.DUT.huff_tree[3] [7] <= \mchip.DUT.node_sorter_ins.output_node [22];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[3] [8] <= 1'h0;
		else if (_0008_)
			\mchip.DUT.huff_tree[3] [8] <= \mchip.DUT.node_sorter_ins.output_node [23];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[3] [9] <= 1'h0;
		else if (_0008_)
			\mchip.DUT.huff_tree[3] [9] <= \mchip.DUT.node_sorter_ins.output_node [24];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[3] [10] <= 1'h0;
		else if (_0008_)
			\mchip.DUT.huff_tree[3] [10] <= \mchip.DUT.node_sorter_ins.output_node [25];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[3] [11] <= 1'h0;
		else if (_0008_)
			\mchip.DUT.huff_tree[3] [11] <= \mchip.DUT.node_sorter_ins.output_node [26];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[3] [12] <= 1'h0;
		else if (_0008_)
			\mchip.DUT.huff_tree[3] [12] <= \mchip.DUT.node_sorter_ins.output_node [27];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[3] [13] <= 1'h0;
		else if (_0008_)
			\mchip.DUT.huff_tree[3] [13] <= \mchip.DUT.node_sorter_ins.output_node [28];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[3] [14] <= 1'h0;
		else if (_0008_)
			\mchip.DUT.huff_tree[3] [14] <= \mchip.DUT.node_sorter_ins.output_node [29];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[3] [15] <= 1'h0;
		else if (_0008_)
			\mchip.DUT.huff_tree[3] [15] <= \mchip.DUT.node_sorter_ins.output_node [33];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[3] [16] <= 1'h0;
		else if (_0008_)
			\mchip.DUT.huff_tree[3] [16] <= \mchip.DUT.node_sorter_ins.output_node [34];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[3] [17] <= 1'h0;
		else if (_0008_)
			\mchip.DUT.huff_tree[3] [17] <= \mchip.DUT.node_sorter_ins.output_node [35];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[3] [18] <= 1'h0;
		else if (_0008_)
			\mchip.DUT.huff_tree[3] [18] <= \mchip.DUT.node_sorter_ins.output_node [36];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[3] [19] <= 1'h0;
		else if (_0008_)
			\mchip.DUT.huff_tree[3] [19] <= \mchip.DUT.node_sorter_ins.output_node [37];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[4] [0] <= 1'h0;
		else if (\mchip.DUT.state [4])
			\mchip.DUT.huff_tree[4] [0] <= _1770_[0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[4] [1] <= 1'h0;
		else if (\mchip.DUT.state [4])
			\mchip.DUT.huff_tree[4] [1] <= _1771_[1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[4] [2] <= 1'h0;
		else if (\mchip.DUT.state [4])
			\mchip.DUT.huff_tree[4] [2] <= _0017_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[4] [3] <= 1'h0;
		else if (\mchip.DUT.state [4])
			\mchip.DUT.huff_tree[4] [3] <= _0040_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[5] [4] <= 1'h0;
		else if (_0007_)
			\mchip.DUT.huff_tree[5] [4] <= \mchip.DUT.node_sorter_ins.output_node [19];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[5] [5] <= 1'h0;
		else if (_0007_)
			\mchip.DUT.huff_tree[5] [5] <= \mchip.DUT.node_sorter_ins.output_node [20];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[5] [6] <= 1'h0;
		else if (_0007_)
			\mchip.DUT.huff_tree[5] [6] <= \mchip.DUT.node_sorter_ins.output_node [21];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[5] [7] <= 1'h0;
		else if (_0007_)
			\mchip.DUT.huff_tree[5] [7] <= \mchip.DUT.node_sorter_ins.output_node [22];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[5] [8] <= 1'h0;
		else if (_0007_)
			\mchip.DUT.huff_tree[5] [8] <= \mchip.DUT.node_sorter_ins.output_node [23];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[5] [9] <= 1'h0;
		else if (_0007_)
			\mchip.DUT.huff_tree[5] [9] <= \mchip.DUT.node_sorter_ins.output_node [24];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[5] [10] <= 1'h0;
		else if (_0007_)
			\mchip.DUT.huff_tree[5] [10] <= \mchip.DUT.node_sorter_ins.output_node [25];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[5] [11] <= 1'h0;
		else if (_0007_)
			\mchip.DUT.huff_tree[5] [11] <= \mchip.DUT.node_sorter_ins.output_node [26];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[5] [12] <= 1'h0;
		else if (_0007_)
			\mchip.DUT.huff_tree[5] [12] <= \mchip.DUT.node_sorter_ins.output_node [27];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[5] [13] <= 1'h0;
		else if (_0007_)
			\mchip.DUT.huff_tree[5] [13] <= \mchip.DUT.node_sorter_ins.output_node [28];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[5] [14] <= 1'h0;
		else if (_0007_)
			\mchip.DUT.huff_tree[5] [14] <= \mchip.DUT.node_sorter_ins.output_node [29];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[5] [15] <= 1'h0;
		else if (_0007_)
			\mchip.DUT.huff_tree[5] [15] <= \mchip.DUT.node_sorter_ins.output_node [33];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[5] [16] <= 1'h0;
		else if (_0007_)
			\mchip.DUT.huff_tree[5] [16] <= \mchip.DUT.node_sorter_ins.output_node [34];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[5] [17] <= 1'h0;
		else if (_0007_)
			\mchip.DUT.huff_tree[5] [17] <= \mchip.DUT.node_sorter_ins.output_node [35];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[5] [18] <= 1'h0;
		else if (_0007_)
			\mchip.DUT.huff_tree[5] [18] <= \mchip.DUT.node_sorter_ins.output_node [36];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.DUT.huff_tree[5] [19] <= 1'h0;
		else if (_0007_)
			\mchip.DUT.huff_tree[5] [19] <= \mchip.DUT.node_sorter_ins.output_node [37];
	always @(posedge io_in[12]) \mchip.DUT.node_sorter_ins.output_node [0] <= _0141_;
	always @(posedge io_in[12]) \mchip.DUT.node_sorter_ins.output_node [1] <= _0152_;
	always @(posedge io_in[12]) \mchip.DUT.node_sorter_ins.output_node [2] <= _0163_;
	always @(posedge io_in[12]) \mchip.DUT.node_sorter_ins.output_node [3] <= _0174_;
	always @(posedge io_in[12]) \mchip.DUT.node_sorter_ins.output_node [4] <= _0185_;
	always @(posedge io_in[12]) \mchip.DUT.node_sorter_ins.output_node [5] <= _0193_;
	always @(posedge io_in[12]) \mchip.DUT.node_sorter_ins.output_node [6] <= _0194_;
	always @(posedge io_in[12]) \mchip.DUT.node_sorter_ins.output_node [7] <= _0195_;
	always @(posedge io_in[12]) \mchip.DUT.node_sorter_ins.output_node [8] <= _0196_;
	always @(posedge io_in[12]) \mchip.DUT.node_sorter_ins.output_node [9] <= _0197_;
	always @(posedge io_in[12]) \mchip.DUT.node_sorter_ins.output_node [10] <= _0142_;
	always @(posedge io_in[12]) \mchip.DUT.node_sorter_ins.output_node [11] <= _0143_;
	always @(posedge io_in[12]) \mchip.DUT.node_sorter_ins.output_node [12] <= _0144_;
	always @(posedge io_in[12]) \mchip.DUT.node_sorter_ins.output_node [13] <= _0145_;
	always @(posedge io_in[12]) \mchip.DUT.node_sorter_ins.output_node [14] <= _0146_;
	always @(posedge io_in[12]) \mchip.DUT.node_sorter_ins.output_node [15] <= _0147_;
	always @(posedge io_in[12]) \mchip.DUT.node_sorter_ins.output_node [16] <= _0148_;
	always @(posedge io_in[12]) \mchip.DUT.node_sorter_ins.output_node [17] <= _0149_;
	always @(posedge io_in[12]) \mchip.DUT.node_sorter_ins.output_node [18] <= _0150_;
	always @(posedge io_in[12]) \mchip.DUT.node_sorter_ins.output_node [19] <= _0151_;
	always @(posedge io_in[12]) \mchip.DUT.node_sorter_ins.output_node [20] <= _0153_;
	always @(posedge io_in[12]) \mchip.DUT.node_sorter_ins.output_node [21] <= _0154_;
	always @(posedge io_in[12]) \mchip.DUT.node_sorter_ins.output_node [22] <= _0155_;
	always @(posedge io_in[12]) \mchip.DUT.node_sorter_ins.output_node [23] <= _0156_;
	always @(posedge io_in[12]) \mchip.DUT.node_sorter_ins.output_node [24] <= _0157_;
	always @(posedge io_in[12]) \mchip.DUT.node_sorter_ins.output_node [25] <= _0158_;
	always @(posedge io_in[12]) \mchip.DUT.node_sorter_ins.output_node [26] <= _0159_;
	always @(posedge io_in[12]) \mchip.DUT.node_sorter_ins.output_node [27] <= _0160_;
	always @(posedge io_in[12]) \mchip.DUT.node_sorter_ins.output_node [28] <= _0161_;
	always @(posedge io_in[12]) \mchip.DUT.node_sorter_ins.output_node [29] <= _0162_;
	always @(posedge io_in[12]) \mchip.DUT.node_sorter_ins.output_node [30] <= _0164_;
	always @(posedge io_in[12]) \mchip.DUT.node_sorter_ins.output_node [31] <= _0165_;
	always @(posedge io_in[12]) \mchip.DUT.node_sorter_ins.output_node [32] <= _0166_;
	always @(posedge io_in[12]) \mchip.DUT.node_sorter_ins.output_node [33] <= _0167_;
	always @(posedge io_in[12]) \mchip.DUT.node_sorter_ins.output_node [34] <= _0168_;
	always @(posedge io_in[12]) \mchip.DUT.node_sorter_ins.output_node [35] <= _0169_;
	always @(posedge io_in[12]) \mchip.DUT.node_sorter_ins.output_node [36] <= _0170_;
	always @(posedge io_in[12]) \mchip.DUT.node_sorter_ins.output_node [37] <= _0171_;
	always @(posedge io_in[12]) \mchip.DUT.node_sorter_ins.output_node [38] <= _0172_;
	always @(posedge io_in[12]) \mchip.DUT.node_sorter_ins.output_node [39] <= _0173_;
	always @(posedge io_in[12]) \mchip.DUT.node_sorter_ins.output_node [40] <= _0175_;
	always @(posedge io_in[12]) \mchip.DUT.node_sorter_ins.output_node [41] <= _0176_;
	always @(posedge io_in[12]) \mchip.DUT.node_sorter_ins.output_node [42] <= _0177_;
	always @(posedge io_in[12]) \mchip.DUT.node_sorter_ins.output_node [43] <= _0178_;
	always @(posedge io_in[12]) \mchip.DUT.node_sorter_ins.output_node [44] <= _0179_;
	always @(posedge io_in[12]) \mchip.DUT.node_sorter_ins.output_node [45] <= _0180_;
	always @(posedge io_in[12]) \mchip.DUT.node_sorter_ins.output_node [46] <= _0181_;
	always @(posedge io_in[12]) \mchip.DUT.node_sorter_ins.output_node [47] <= _0182_;
	always @(posedge io_in[12]) \mchip.DUT.node_sorter_ins.output_node [48] <= _0183_;
	always @(posedge io_in[12]) \mchip.DUT.node_sorter_ins.output_node [49] <= _0184_;
	always @(posedge io_in[12]) \mchip.DUT.node_sorter_ins.output_node [50] <= _0186_;
	always @(posedge io_in[12]) \mchip.DUT.node_sorter_ins.output_node [51] <= _0187_;
	always @(posedge io_in[12]) \mchip.DUT.node_sorter_ins.output_node [52] <= _0188_;
	always @(posedge io_in[12]) \mchip.DUT.node_sorter_ins.output_node [53] <= _0189_;
	always @(posedge io_in[12]) \mchip.DUT.node_sorter_ins.output_node [54] <= _0190_;
	always @(posedge io_in[12]) \mchip.DUT.node_sorter_ins.output_node [55] <= _0191_;
	always @(posedge io_in[12]) \mchip.DUT.node_sorter_ins.output_node [56] <= _0192_;
	assign _1766_[1] = 1'h0;
	assign _1767_[0] = _1766_[0];
	assign _1768_[1] = 1'h0;
	assign _1769_[0] = _1768_[0];
	assign _1770_[1] = 1'h0;
	assign _1771_[0] = _1770_[0];
	assign _1772_[1] = 1'h0;
	assign _1773_[0] = _1772_[0];
	assign _1774_[2:1] = 2'h0;
	assign io_out = {5'h00, \mchip.DUT.io_out [8], 1'h0, \mchip.DUT.io_out [6:0]};
	assign \mchip.DUT.b [2:1] = 2'h0;
	assign \mchip.DUT.clk  = io_in[12];
	assign {\mchip.DUT.data_in [23:21], \mchip.DUT.data_in [15:13], \mchip.DUT.data_in [7:5]} = 9'h000;
	assign \mchip.DUT.encoded_value_h[0]  = 3'h0;
	assign \mchip.DUT.encoded_value_h[1]  = 3'h0;
	assign \mchip.DUT.freq_calc_ins.data_in  = {3'h0, \mchip.DUT.data_in [20:16], 3'h0, \mchip.DUT.data_in [12:8], 3'h0, \mchip.DUT.data_in [4:0]};
	assign \mchip.DUT.freq_calc_ins.freq_in  = \mchip.DUT.freq_in ;
	assign \mchip.DUT.freq_calc_ins.node  = {\mchip.DUT.data_in [20:16], \mchip.DUT.freq_in [8:6], 11'h400, \mchip.DUT.data_in [12:8], \mchip.DUT.freq_in [5:3], 11'h400, \mchip.DUT.data_in [4:0], \mchip.DUT.freq_in [2:0], 11'h400};
	assign \mchip.DUT.freq_calc_ins.sv2v_autoblock_1.i  = 32'd3;
	assign \mchip.DUT.huff_tree[0]  = 20'h00000;
	assign \mchip.DUT.huff_tree[1] [3:0] = 4'h0;
	assign \mchip.DUT.in_huff_tree [9:0] = 10'h000;
	assign \mchip.DUT.initial_node  = {\mchip.DUT.data_in [20:16], \mchip.DUT.freq_in [8:6], 11'h400, \mchip.DUT.data_in [12:8], \mchip.DUT.freq_in [5:3], 11'h400, \mchip.DUT.data_in [4:0], \mchip.DUT.freq_in [2:0], 11'h400};
	assign \mchip.DUT.io_in  = io_in[11:0];
	assign {\mchip.DUT.io_out [11:9], \mchip.DUT.io_out [7]} = 4'h0;
	assign \mchip.DUT.merge_nodes_ins.merged_node  = {9'h000, \mchip.DUT.node_sorter_ins.output_node [56:52], \mchip.DUT.node_sorter_ins.output_node [37:33]};
	assign \mchip.DUT.merge_nodes_ins.min_node  = \mchip.DUT.node_sorter_ins.output_node [56:38];
	assign \mchip.DUT.merge_nodes_ins.second_min_node  = \mchip.DUT.node_sorter_ins.output_node [37:19];
	assign \mchip.DUT.merged_node  = {9'h000, \mchip.DUT.node_sorter_ins.output_node [56:52], \mchip.DUT.node_sorter_ins.output_node [37:33]};
	assign \mchip.DUT.node_sorter_ins.clk  = io_in[12];
	assign \mchip.DUT.node_sorter_ins.input_node  = {\mchip.DUT.in_huff_tree [56:10], 10'h000};
	assign \mchip.DUT.out_huff_tree  = {\mchip.DUT.node_sorter_ins.output_node , 19'h00000};
	assign \mchip.DUT.reset  = io_in[13];
	assign \mchip.clock  = io_in[12];
	assign \mchip.io_in  = io_in[11:0];
	assign \mchip.io_out  = {3'h0, \mchip.DUT.io_out [8], 1'h0, \mchip.DUT.io_out [6:0]};
	assign \mchip.reset  = io_in[13];
endmodule
module d26_cjstange_perceptron (
	io_in,
	io_out
);
	wire _0000_;
	wire _0001_;
	wire _0002_;
	wire _0003_;
	wire _0004_;
	wire _0005_;
	wire _0006_;
	wire _0007_;
	wire _0008_;
	wire _0009_;
	wire _0010_;
	wire _0011_;
	wire _0012_;
	wire _0013_;
	wire _0014_;
	wire _0015_;
	wire _0016_;
	wire _0017_;
	wire _0018_;
	wire _0019_;
	wire _0020_;
	wire _0021_;
	wire _0022_;
	wire _0023_;
	wire _0024_;
	wire _0025_;
	wire _0026_;
	wire _0027_;
	wire _0028_;
	wire _0029_;
	wire _0030_;
	wire _0031_;
	wire _0032_;
	wire _0033_;
	wire _0034_;
	wire _0035_;
	wire _0036_;
	wire _0037_;
	wire _0038_;
	wire _0039_;
	wire _0040_;
	wire _0041_;
	wire _0042_;
	wire _0043_;
	wire _0044_;
	wire _0045_;
	wire _0046_;
	wire _0047_;
	wire _0048_;
	wire _0049_;
	wire _0050_;
	wire _0051_;
	wire _0052_;
	wire _0053_;
	wire _0054_;
	wire _0055_;
	wire _0056_;
	wire _0057_;
	wire _0058_;
	wire _0059_;
	wire _0060_;
	wire _0061_;
	wire _0062_;
	wire _0063_;
	wire _0064_;
	wire _0065_;
	wire _0066_;
	wire _0067_;
	wire _0068_;
	wire _0069_;
	wire _0070_;
	wire _0071_;
	wire _0072_;
	wire _0073_;
	wire _0074_;
	wire _0075_;
	wire _0076_;
	wire _0077_;
	wire _0078_;
	wire _0079_;
	wire _0080_;
	wire _0081_;
	wire _0082_;
	wire _0083_;
	wire _0084_;
	wire _0085_;
	wire _0086_;
	wire _0087_;
	wire _0088_;
	wire _0089_;
	wire _0090_;
	wire _0091_;
	wire _0092_;
	wire _0093_;
	wire _0094_;
	wire _0095_;
	wire _0096_;
	wire _0097_;
	wire _0098_;
	wire _0099_;
	wire _0100_;
	wire _0101_;
	wire _0102_;
	wire _0103_;
	wire _0104_;
	wire _0105_;
	wire _0106_;
	wire _0107_;
	wire _0108_;
	wire _0109_;
	wire _0110_;
	wire _0111_;
	wire _0112_;
	wire _0113_;
	wire _0114_;
	wire _0115_;
	wire _0116_;
	wire _0117_;
	wire _0118_;
	wire _0119_;
	wire _0120_;
	wire _0121_;
	wire _0122_;
	wire _0123_;
	wire _0124_;
	wire _0125_;
	wire _0126_;
	wire _0127_;
	wire _0128_;
	wire _0129_;
	wire _0130_;
	wire _0131_;
	wire _0132_;
	wire _0133_;
	wire _0134_;
	wire _0135_;
	wire _0136_;
	wire _0137_;
	wire _0138_;
	wire _0139_;
	wire _0140_;
	wire _0141_;
	wire _0142_;
	wire _0143_;
	wire _0144_;
	wire _0145_;
	wire _0146_;
	wire _0147_;
	wire _0148_;
	wire _0149_;
	wire _0150_;
	wire _0151_;
	wire _0152_;
	wire _0153_;
	wire _0154_;
	wire _0155_;
	wire _0156_;
	wire _0157_;
	wire _0158_;
	wire _0159_;
	wire _0160_;
	wire _0161_;
	wire _0162_;
	wire _0163_;
	wire _0164_;
	wire _0165_;
	wire _0166_;
	wire _0167_;
	wire _0168_;
	wire _0169_;
	wire _0170_;
	wire _0171_;
	wire _0172_;
	wire _0173_;
	wire _0174_;
	wire _0175_;
	wire _0176_;
	wire _0177_;
	wire _0178_;
	wire _0179_;
	wire _0180_;
	wire _0181_;
	wire _0182_;
	wire _0183_;
	wire _0184_;
	wire _0185_;
	wire _0186_;
	wire _0187_;
	wire _0188_;
	wire _0189_;
	wire _0190_;
	wire _0191_;
	wire _0192_;
	wire _0193_;
	wire _0194_;
	wire _0195_;
	wire _0196_;
	wire _0197_;
	wire _0198_;
	wire _0199_;
	wire _0200_;
	wire _0201_;
	wire _0202_;
	wire _0203_;
	wire _0204_;
	wire _0205_;
	wire _0206_;
	wire _0207_;
	wire _0208_;
	wire _0209_;
	wire _0210_;
	wire _0211_;
	wire _0212_;
	wire _0213_;
	wire _0214_;
	wire _0215_;
	wire _0216_;
	wire _0217_;
	wire _0218_;
	wire _0219_;
	wire _0220_;
	wire _0221_;
	wire _0222_;
	wire _0223_;
	wire _0224_;
	wire _0225_;
	wire _0226_;
	wire _0227_;
	wire _0228_;
	wire _0229_;
	wire _0230_;
	wire _0231_;
	wire _0232_;
	wire _0233_;
	wire _0234_;
	wire _0235_;
	wire _0236_;
	wire _0237_;
	wire _0238_;
	wire _0239_;
	wire _0240_;
	wire _0241_;
	wire _0242_;
	wire _0243_;
	wire _0244_;
	wire _0245_;
	wire _0246_;
	wire _0247_;
	wire _0248_;
	wire _0249_;
	wire _0250_;
	wire _0251_;
	wire _0252_;
	wire _0253_;
	wire _0254_;
	wire _0255_;
	wire _0256_;
	wire _0257_;
	wire _0258_;
	wire _0259_;
	wire _0260_;
	wire _0261_;
	wire _0262_;
	wire _0263_;
	wire _0264_;
	wire _0265_;
	wire _0266_;
	wire _0267_;
	wire _0268_;
	wire _0269_;
	wire _0270_;
	wire _0271_;
	wire _0272_;
	wire _0273_;
	wire _0274_;
	wire _0275_;
	wire _0276_;
	wire _0277_;
	wire _0278_;
	wire _0279_;
	wire _0280_;
	wire _0281_;
	wire _0282_;
	wire _0283_;
	wire _0284_;
	wire _0285_;
	wire _0286_;
	wire _0287_;
	wire _0288_;
	wire _0289_;
	wire _0290_;
	wire _0291_;
	wire _0292_;
	wire _0293_;
	wire _0294_;
	wire _0295_;
	wire _0296_;
	wire _0297_;
	wire _0298_;
	wire _0299_;
	wire _0300_;
	wire _0301_;
	wire _0302_;
	wire _0303_;
	wire _0304_;
	wire _0305_;
	wire _0306_;
	wire _0307_;
	wire _0308_;
	wire _0309_;
	wire _0310_;
	wire _0311_;
	wire _0312_;
	wire _0313_;
	wire _0314_;
	wire _0315_;
	wire _0316_;
	wire _0317_;
	wire _0318_;
	wire _0319_;
	wire _0320_;
	wire _0321_;
	wire _0322_;
	wire _0323_;
	wire _0324_;
	wire _0325_;
	wire _0326_;
	wire _0327_;
	wire _0328_;
	wire _0329_;
	wire _0330_;
	wire _0331_;
	wire _0332_;
	wire _0333_;
	wire _0334_;
	wire _0335_;
	wire _0336_;
	wire _0337_;
	wire _0338_;
	wire _0339_;
	wire _0340_;
	wire _0341_;
	wire _0342_;
	wire _0343_;
	wire _0344_;
	wire _0345_;
	wire _0346_;
	wire _0347_;
	wire _0348_;
	wire _0349_;
	wire _0350_;
	wire _0351_;
	wire _0352_;
	wire _0353_;
	wire _0354_;
	wire _0355_;
	wire _0356_;
	wire _0357_;
	wire _0358_;
	wire _0359_;
	wire _0360_;
	wire _0361_;
	wire _0362_;
	wire _0363_;
	wire _0364_;
	wire _0365_;
	wire _0366_;
	wire _0367_;
	wire _0368_;
	wire _0369_;
	wire _0370_;
	wire _0371_;
	wire _0372_;
	wire _0373_;
	wire _0374_;
	wire _0375_;
	wire _0376_;
	wire _0377_;
	wire _0378_;
	wire _0379_;
	wire _0380_;
	wire _0381_;
	wire _0382_;
	wire _0383_;
	wire _0384_;
	wire _0385_;
	wire _0386_;
	wire _0387_;
	wire _0388_;
	wire _0389_;
	wire _0390_;
	wire _0391_;
	wire _0392_;
	wire _0393_;
	wire _0394_;
	wire _0395_;
	wire _0396_;
	wire _0397_;
	wire _0398_;
	wire _0399_;
	wire _0400_;
	wire _0401_;
	wire _0402_;
	wire _0403_;
	wire _0404_;
	wire _0405_;
	wire _0406_;
	wire _0407_;
	wire _0408_;
	wire _0409_;
	wire _0410_;
	wire _0411_;
	wire _0412_;
	wire _0413_;
	wire _0414_;
	wire _0415_;
	wire _0416_;
	wire _0417_;
	wire _0418_;
	wire _0419_;
	wire _0420_;
	wire _0421_;
	wire _0422_;
	wire _0423_;
	wire _0424_;
	wire _0425_;
	wire _0426_;
	wire _0427_;
	wire _0428_;
	wire _0429_;
	wire _0430_;
	wire _0431_;
	wire _0432_;
	wire _0433_;
	wire _0434_;
	wire _0435_;
	wire _0436_;
	wire _0437_;
	wire _0438_;
	wire _0439_;
	wire _0440_;
	wire _0441_;
	wire _0442_;
	wire _0443_;
	wire _0444_;
	wire _0445_;
	wire _0446_;
	wire _0447_;
	wire _0448_;
	wire _0449_;
	wire _0450_;
	wire _0451_;
	wire _0452_;
	wire _0453_;
	wire _0454_;
	wire _0455_;
	wire _0456_;
	wire _0457_;
	wire _0458_;
	wire _0459_;
	wire _0460_;
	wire _0461_;
	wire _0462_;
	wire _0463_;
	wire _0464_;
	wire _0465_;
	wire _0466_;
	wire _0467_;
	wire _0468_;
	wire _0469_;
	wire _0470_;
	wire _0471_;
	wire _0472_;
	wire _0473_;
	wire _0474_;
	wire _0475_;
	wire _0476_;
	wire _0477_;
	wire _0478_;
	wire _0479_;
	wire _0480_;
	wire _0481_;
	wire _0482_;
	wire _0483_;
	wire _0484_;
	wire _0485_;
	wire _0486_;
	wire _0487_;
	wire _0488_;
	wire _0489_;
	wire _0490_;
	wire _0491_;
	wire _0492_;
	wire _0493_;
	wire _0494_;
	wire _0495_;
	wire _0496_;
	wire _0497_;
	wire _0498_;
	wire _0499_;
	wire _0500_;
	wire _0501_;
	wire _0502_;
	wire _0503_;
	wire _0504_;
	wire _0505_;
	wire _0506_;
	wire _0507_;
	wire _0508_;
	wire _0509_;
	wire _0510_;
	wire _0511_;
	wire _0512_;
	wire _0513_;
	wire _0514_;
	wire _0515_;
	wire _0516_;
	wire _0517_;
	wire _0518_;
	wire _0519_;
	wire _0520_;
	wire _0521_;
	wire _0522_;
	wire _0523_;
	wire _0524_;
	wire _0525_;
	wire _0526_;
	wire _0527_;
	wire _0528_;
	wire _0529_;
	wire _0530_;
	wire _0531_;
	wire _0532_;
	wire _0533_;
	wire _0534_;
	wire _0535_;
	wire _0536_;
	wire _0537_;
	wire _0538_;
	wire _0539_;
	wire _0540_;
	wire _0541_;
	wire _0542_;
	wire _0543_;
	wire _0544_;
	wire _0545_;
	wire _0546_;
	wire _0547_;
	wire _0548_;
	wire _0549_;
	wire _0550_;
	wire _0551_;
	wire _0552_;
	wire [1:0] _0553_;
	wire [1:0] _0554_;
	input wire [13:0] io_in;
	output wire [13:0] io_out;
	wire \mchip.clock ;
	wire [11:0] \mchip.io_in ;
	wire [11:0] \mchip.io_out ;
	wire \mchip.learning.classification ;
	wire \mchip.learning.clk ;
	wire \mchip.learning.control.classification ;
	wire \mchip.learning.control.clk ;
	wire \mchip.learning.control.correct ;
	wire [1:0] \mchip.learning.control.count ;
	wire \mchip.learning.control.done ;
	wire \mchip.learning.control.en_add ;
	wire \mchip.learning.control.en_count ;
	wire \mchip.learning.control.en_mult ;
	wire \mchip.learning.control.en_n ;
	wire \mchip.learning.control.en_w0 ;
	wire \mchip.learning.control.en_w1 ;
	wire \mchip.learning.control.en_w2 ;
	wire \mchip.learning.control.en_x1 ;
	wire \mchip.learning.control.en_x2 ;
	wire \mchip.learning.control.go ;
	wire \mchip.learning.control.sel_add_A ;
	reg [10:0] \mchip.learning.control.state ;
	wire \mchip.learning.control.sync ;
	wire \mchip.learning.control.update ;
	wire \mchip.learning.correct ;
	wire [1:0] \mchip.learning.count ;
	wire \mchip.learning.data.add.cin ;
	wire [5:0] \mchip.learning.data.add.sum ;
	wire [11:0] \mchip.learning.data.add_A_mux.in ;
	wire \mchip.learning.data.add_A_mux.sel ;
	wire [23:0] \mchip.learning.data.add_B_mux.in ;
	wire [5:0] \mchip.learning.data.add_out ;
	wire [5:0] \mchip.learning.data.add_out_reg ;
	wire [5:0] \mchip.learning.data.add_reg.D ;
	reg [5:0] \mchip.learning.data.add_reg.Q ;
	wire \mchip.learning.data.add_reg.clk ;
	wire \mchip.learning.data.add_reg.en ;
	wire \mchip.learning.data.classification ;
	wire \mchip.learning.data.clk ;
	wire \mchip.learning.data.correct ;
	wire [1:0] \mchip.learning.data.count ;
	wire \mchip.learning.data.counter.clk ;
	reg [1:0] \mchip.learning.data.counter.count ;
	wire \mchip.learning.data.counter.en ;
	wire [5:0] \mchip.learning.data.d ;
	wire \mchip.learning.data.en_add ;
	wire \mchip.learning.data.en_count ;
	wire \mchip.learning.data.en_mult ;
	wire \mchip.learning.data.en_n ;
	wire \mchip.learning.data.en_w0 ;
	wire \mchip.learning.data.en_w1 ;
	wire \mchip.learning.data.en_w2 ;
	wire \mchip.learning.data.en_x1 ;
	wire \mchip.learning.data.en_x2 ;
	wire [5:0] \mchip.learning.data.in_val ;
	wire [23:0] \mchip.learning.data.input_mux.in ;
	wire [5:0] \mchip.learning.data.input_mux.out ;
	wire [1:0] \mchip.learning.data.input_mux.sel ;
	wire [5:0] \mchip.learning.data.mult.M ;
	wire [11:0] \mchip.learning.data.mult.tmp ;
	wire [23:0] \mchip.learning.data.mult_A_mux.in ;
	wire [23:0] \mchip.learning.data.mult_B_mux.in ;
	wire [5:0] \mchip.learning.data.mult_out ;
	wire [5:0] \mchip.learning.data.mult_out_reg ;
	wire [5:0] \mchip.learning.data.mult_reg.D ;
	reg [5:0] \mchip.learning.data.mult_reg.Q ;
	wire \mchip.learning.data.mult_reg.clk ;
	wire \mchip.learning.data.mult_reg.en ;
	wire [5:0] \mchip.learning.data.n ;
	wire [5:0] \mchip.learning.data.n_reg.D ;
	reg [5:0] \mchip.learning.data.n_reg.Q ;
	wire \mchip.learning.data.n_reg.clk ;
	wire \mchip.learning.data.n_reg.en ;
	wire [5:0] \mchip.learning.data.out_val ;
	wire \mchip.learning.data.sel_add_A ;
	wire [1:0] \mchip.learning.data.sel_out ;
	wire [5:0] \mchip.learning.data.w0 ;
	wire [5:0] \mchip.learning.data.w0_reg.D ;
	reg [5:0] \mchip.learning.data.w0_reg.Q ;
	wire \mchip.learning.data.w0_reg.clk ;
	wire \mchip.learning.data.w0_reg.en ;
	wire [5:0] \mchip.learning.data.w1 ;
	wire [5:0] \mchip.learning.data.w1_reg.D ;
	reg [5:0] \mchip.learning.data.w1_reg.Q ;
	wire \mchip.learning.data.w1_reg.clk ;
	wire \mchip.learning.data.w1_reg.en ;
	wire [5:0] \mchip.learning.data.w2 ;
	wire [5:0] \mchip.learning.data.w2_reg.D ;
	reg [5:0] \mchip.learning.data.w2_reg.Q ;
	wire \mchip.learning.data.w2_reg.clk ;
	wire \mchip.learning.data.w2_reg.en ;
	wire [5:0] \mchip.learning.data.x1 ;
	wire [5:0] \mchip.learning.data.x1_reg.D ;
	reg [5:0] \mchip.learning.data.x1_reg.Q ;
	wire \mchip.learning.data.x1_reg.clk ;
	wire \mchip.learning.data.x1_reg.en ;
	wire [5:0] \mchip.learning.data.x2 ;
	wire [5:0] \mchip.learning.data.x2_reg.D ;
	reg [5:0] \mchip.learning.data.x2_reg.Q ;
	wire \mchip.learning.data.x2_reg.clk ;
	wire \mchip.learning.data.x2_reg.en ;
	wire \mchip.learning.done ;
	wire \mchip.learning.en_add ;
	wire \mchip.learning.en_count ;
	wire \mchip.learning.en_mult ;
	wire \mchip.learning.en_n ;
	wire \mchip.learning.en_w0 ;
	wire \mchip.learning.en_w1 ;
	wire \mchip.learning.en_w2 ;
	wire \mchip.learning.en_x1 ;
	wire \mchip.learning.en_x2 ;
	wire \mchip.learning.go ;
	wire [5:0] \mchip.learning.in_val ;
	wire [5:0] \mchip.learning.out_val ;
	wire \mchip.learning.sel_add_A ;
	wire [1:0] \mchip.learning.sel_out ;
	wire \mchip.learning.sync ;
	wire \mchip.learning.update ;
	wire \mchip.reset ;
	assign _0553_[0] = ~\mchip.learning.data.counter.count [0];
	assign _0012_ = io_in[9] | io_in[13];
	assign _0013_ = \mchip.learning.control.state [10] & ~_0012_;
	assign _0014_ = io_in[10] | io_in[13];
	assign _0015_ = \mchip.learning.control.state [2] & ~_0014_;
	assign _0016_ = _0015_ | _0013_;
	assign _0017_ = io_in[13] | ~io_in[10];
	assign _0018_ = \mchip.learning.control.state [9] & ~_0017_;
	assign _0019_ = \mchip.learning.data.counter.count [1] & \mchip.learning.data.counter.count [0];
	assign _0020_ = ~io_in[8];
	assign _0021_ = \mchip.learning.data.add_reg.Q [3] | \mchip.learning.data.add_reg.Q [4];
	assign \mchip.learning.classification  = _0021_ & ~\mchip.learning.data.add_reg.Q [5];
	assign _0022_ = \mchip.learning.classification  ^ _0020_;
	assign _0023_ = _0022_ | _0019_;
	assign _0024_ = io_in[13] | ~_0023_;
	assign _0025_ = \mchip.learning.control.state [1] & ~_0024_;
	assign _0026_ = _0025_ | _0018_;
	assign _0006_ = _0026_ | _0016_;
	assign \mchip.learning.control.en_x2  = \mchip.learning.control.state [8] & io_in[10];
	assign \mchip.learning.control.en_x1  = \mchip.learning.control.state [2] & io_in[10];
	assign _0027_ = \mchip.learning.control.state [9] & ~_0014_;
	assign _0028_ = \mchip.learning.control.state [3] & ~_0017_;
	assign _0010_ = _0028_ | _0027_;
	assign _0029_ = \mchip.learning.control.state [8] & ~_0014_;
	assign _0030_ = \mchip.learning.control.state [2] & ~_0017_;
	assign _0009_ = _0030_ | _0029_;
	assign _0031_ = \mchip.learning.control.state [6] & ~_0014_;
	assign _0032_ = \mchip.learning.control.state [0] & ~_0017_;
	assign _0008_ = _0032_ | _0031_;
	assign _0033_ = \mchip.learning.control.state [3] & ~_0014_;
	assign _0034_ = \mchip.learning.control.state [6] & ~_0017_;
	assign _0007_ = _0034_ | _0033_;
	assign _0035_ = io_in[13] | ~io_in[9];
	assign _0036_ = \mchip.learning.control.state [10] & ~_0035_;
	assign _0037_ = \mchip.learning.control.state [4] & ~io_in[13];
	assign _0005_ = _0037_ | _0036_;
	assign _0038_ = \mchip.learning.control.state [10] & io_in[9];
	assign _0011_ = _0038_ | io_in[13];
	assign _0039_ = \mchip.learning.control.state [0] & ~_0014_;
	assign _0004_ = _0039_ | io_in[13];
	assign _0040_ = ~\mchip.learning.control.state [2];
	assign _0041_ = \mchip.learning.control.state [5] | \mchip.learning.control.state [10];
	assign _0042_ = _0041_ | \mchip.learning.control.state [4];
	assign _0043_ = _0040_ & ~_0042_;
	assign _0044_ = ~\mchip.learning.control.en_x1 ;
	assign _0045_ = \mchip.learning.data.counter.count [1] | ~\mchip.learning.data.counter.count [0];
	assign _0046_ = ~(\mchip.learning.data.counter.count [1] | \mchip.learning.data.counter.count [0]);
	assign _0047_ = _0045_ & ~_0046_;
	assign _0048_ = \mchip.learning.control.state [4] & ~_0047_;
	assign _0049_ = _0044_ & ~_0048_;
	assign _0050_ = _0049_ | _0043_;
	assign _0051_ = _0046_ & \mchip.learning.control.state [4];
	assign _0052_ = _0051_ | _0041_;
	assign _0053_ = _0044_ & ~_0052_;
	assign _0054_ = _0053_ | _0043_;
	assign _0055_ = ~(_0054_ | _0050_);
	assign _0056_ = ~\mchip.learning.data.w0_reg.Q [2];
	assign _0057_ = ~\mchip.learning.data.w0_reg.Q [4];
	assign _0058_ = (_0050_ ? _0056_ : _0057_);
	assign _0059_ = _0054_ ^ _0050_;
	assign _0060_ = (_0050_ ? \mchip.learning.data.add_reg.Q [4] : \mchip.learning.data.w0_reg.Q [0]);
	assign _0061_ = ~_0060_;
	assign _0062_ = (_0059_ ? _0058_ : _0061_);
	assign _0063_ = _0050_ & ~_0054_;
	assign _0064_ = ~(_0063_ | _0062_);
	assign _0065_ = (_0050_ ? \mchip.learning.data.add_reg.Q [0] : \mchip.learning.data.add_reg.Q [2]);
	assign _0066_ = (_0050_ ? \mchip.learning.data.w1_reg.Q [2] : \mchip.learning.data.w1_reg.Q [4]);
	assign _0067_ = (_0059_ ? _0065_ : _0066_);
	assign _0068_ = (_0050_ ? \mchip.learning.data.w2_reg.Q [4] : \mchip.learning.data.w1_reg.Q [0]);
	assign _0069_ = (_0050_ ? \mchip.learning.data.w2_reg.Q [0] : \mchip.learning.data.w2_reg.Q [2]);
	assign _0070_ = (_0059_ ? _0068_ : _0069_);
	assign _0071_ = (_0063_ ? _0067_ : _0070_);
	assign _0072_ = (_0055_ ? _0064_ : _0071_);
	assign _0073_ = ~\mchip.learning.data.mult_reg.Q [0];
	assign _0074_ = ~\mchip.learning.data.mult_reg.Q [2];
	assign _0075_ = (\mchip.learning.control.en_x1  ? _0074_ : _0073_);
	assign _0076_ = \mchip.learning.data.mult_reg.Q [4] & ~\mchip.learning.control.en_x1 ;
	assign _0077_ = ~_0076_;
	assign _0078_ = (\mchip.learning.control.en_x1  ? _0077_ : _0075_);
	assign \mchip.learning.data.add_out [0] = ~(_0078_ ^ _0072_);
	assign _0079_ = \mchip.learning.control.state [3] & io_in[10];
	assign \mchip.learning.data.w2_reg.D [0] = (_0079_ ? io_in[0] : \mchip.learning.data.add_out [0]);
	assign _0080_ = _0072_ & ~_0078_;
	assign _0081_ = ~\mchip.learning.data.w0_reg.Q [3];
	assign _0082_ = ~\mchip.learning.data.w0_reg.Q [5];
	assign _0083_ = (_0050_ ? _0081_ : _0082_);
	assign _0084_ = (_0050_ ? \mchip.learning.data.add_reg.Q [5] : \mchip.learning.data.w0_reg.Q [1]);
	assign _0085_ = ~_0084_;
	assign _0086_ = (_0059_ ? _0083_ : _0085_);
	assign _0087_ = ~(_0086_ | _0063_);
	assign _0088_ = (_0050_ ? \mchip.learning.data.add_reg.Q [1] : \mchip.learning.data.add_reg.Q [3]);
	assign _0089_ = (_0050_ ? \mchip.learning.data.w1_reg.Q [3] : \mchip.learning.data.w1_reg.Q [5]);
	assign _0090_ = (_0059_ ? _0088_ : _0089_);
	assign _0091_ = (_0050_ ? \mchip.learning.data.w2_reg.Q [5] : \mchip.learning.data.w1_reg.Q [1]);
	assign _0092_ = (_0050_ ? \mchip.learning.data.w2_reg.Q [1] : \mchip.learning.data.w2_reg.Q [3]);
	assign _0093_ = (_0059_ ? _0091_ : _0092_);
	assign _0094_ = (_0063_ ? _0090_ : _0093_);
	assign _0095_ = (_0055_ ? _0087_ : _0094_);
	assign _0096_ = (\mchip.learning.control.en_x1  ? \mchip.learning.data.mult_reg.Q [3] : \mchip.learning.data.mult_reg.Q [1]);
	assign _0097_ = \mchip.learning.data.mult_reg.Q [5] & ~\mchip.learning.control.en_x1 ;
	assign _0098_ = (\mchip.learning.control.en_x1  ? _0097_ : _0096_);
	assign _0099_ = ~_0098_;
	assign _0100_ = _0099_ ^ _0095_;
	assign \mchip.learning.data.add_out [1] = ~(_0100_ ^ _0080_);
	assign \mchip.learning.data.w2_reg.D [1] = (_0079_ ? io_in[1] : \mchip.learning.data.add_out [1]);
	assign _0101_ = _0080_ & ~_0100_;
	assign _0102_ = _0095_ & ~_0099_;
	assign _0103_ = _0102_ | _0101_;
	assign _0104_ = _0050_ & ~_0057_;
	assign _0105_ = (_0050_ ? \mchip.learning.data.w0_reg.Q [0] : \mchip.learning.data.w0_reg.Q [2]);
	assign _0106_ = (_0059_ ? _0104_ : _0105_);
	assign _0107_ = _0106_ & ~_0063_;
	assign _0108_ = (_0050_ ? \mchip.learning.data.add_reg.Q [2] : \mchip.learning.data.add_reg.Q [4]);
	assign _0109_ = (_0050_ ? \mchip.learning.data.w1_reg.Q [4] : \mchip.learning.data.add_reg.Q [0]);
	assign _0110_ = (_0059_ ? _0108_ : _0109_);
	assign _0111_ = (_0050_ ? \mchip.learning.data.w1_reg.Q [0] : \mchip.learning.data.w1_reg.Q [2]);
	assign _0112_ = (_0050_ ? \mchip.learning.data.w2_reg.Q [2] : \mchip.learning.data.w2_reg.Q [4]);
	assign _0113_ = (_0059_ ? _0111_ : _0112_);
	assign _0114_ = (_0063_ ? _0110_ : _0113_);
	assign _0115_ = (_0055_ ? _0107_ : _0114_);
	assign _0116_ = ~\mchip.learning.data.mult_reg.Q [4];
	assign _0117_ = (\mchip.learning.control.en_x1  ? _0116_ : _0074_);
	assign _0118_ = _0044_ & ~_0117_;
	assign _0119_ = _0118_ ^ _0115_;
	assign \mchip.learning.data.add_out [2] = _0119_ ^ _0103_;
	assign \mchip.learning.data.w2_reg.D [2] = (_0079_ ? io_in[2] : \mchip.learning.data.add_out [2]);
	assign _0120_ = _0118_ & _0115_;
	assign _0121_ = _0119_ & _0103_;
	assign _0122_ = _0121_ | _0120_;
	assign _0123_ = _0050_ & ~_0082_;
	assign _0124_ = (_0050_ ? \mchip.learning.data.w0_reg.Q [1] : \mchip.learning.data.w0_reg.Q [3]);
	assign _0125_ = (_0059_ ? _0123_ : _0124_);
	assign _0126_ = _0125_ & ~_0063_;
	assign _0127_ = (_0050_ ? \mchip.learning.data.add_reg.Q [3] : \mchip.learning.data.add_reg.Q [5]);
	assign _0128_ = (_0050_ ? \mchip.learning.data.w1_reg.Q [5] : \mchip.learning.data.add_reg.Q [1]);
	assign _0129_ = (_0059_ ? _0127_ : _0128_);
	assign _0130_ = (_0050_ ? \mchip.learning.data.w1_reg.Q [1] : \mchip.learning.data.w1_reg.Q [3]);
	assign _0131_ = (_0050_ ? \mchip.learning.data.w2_reg.Q [3] : \mchip.learning.data.w2_reg.Q [5]);
	assign _0132_ = (_0059_ ? _0130_ : _0131_);
	assign _0133_ = (_0063_ ? _0129_ : _0132_);
	assign _0134_ = (_0055_ ? _0126_ : _0133_);
	assign _0135_ = ~\mchip.learning.data.mult_reg.Q [3];
	assign _0136_ = ~\mchip.learning.data.mult_reg.Q [5];
	assign _0137_ = (\mchip.learning.control.en_x1  ? _0136_ : _0135_);
	assign _0138_ = _0044_ & ~_0137_;
	assign _0139_ = _0138_ ^ _0134_;
	assign \mchip.learning.data.add_out [3] = _0139_ ^ _0122_;
	assign \mchip.learning.data.w2_reg.D [3] = (_0079_ ? io_in[3] : \mchip.learning.data.add_out [3]);
	assign _0140_ = _0138_ & _0134_;
	assign _0141_ = _0139_ & _0120_;
	assign _0142_ = _0141_ | _0140_;
	assign _0143_ = ~(_0139_ & _0119_);
	assign _0144_ = _0103_ & ~_0143_;
	assign _0145_ = _0144_ | _0142_;
	assign _0146_ = _0059_ | _0058_;
	assign _0147_ = ~(_0146_ | _0063_);
	assign _0148_ = (_0059_ ? _0060_ : _0065_);
	assign _0149_ = (_0059_ ? _0066_ : _0068_);
	assign _0150_ = (_0063_ ? _0148_ : _0149_);
	assign _0151_ = (_0055_ ? _0147_ : _0150_);
	assign _0152_ = _0151_ ^ _0076_;
	assign \mchip.learning.data.add_out [4] = _0152_ ^ _0145_;
	assign \mchip.learning.data.w2_reg.D [4] = (_0079_ ? io_in[4] : \mchip.learning.data.add_out [4]);
	assign _0153_ = _0151_ & ~_0077_;
	assign _0154_ = _0152_ & _0145_;
	assign _0155_ = _0154_ | _0153_;
	assign _0156_ = _0083_ | _0059_;
	assign _0157_ = ~(_0156_ | _0063_);
	assign _0158_ = (_0059_ ? _0084_ : _0088_);
	assign _0159_ = (_0059_ ? _0089_ : _0091_);
	assign _0160_ = (_0063_ ? _0158_ : _0159_);
	assign _0161_ = (_0055_ ? _0157_ : _0160_);
	assign _0162_ = _0161_ ^ _0097_;
	assign \mchip.learning.data.add_out [5] = _0162_ ^ _0155_;
	assign \mchip.learning.data.w2_reg.D [5] = (_0079_ ? io_in[5] : \mchip.learning.data.add_out [5]);
	assign _0163_ = \mchip.learning.control.state [6] & io_in[10];
	assign \mchip.learning.data.w1_reg.D [0] = (_0163_ ? io_in[0] : \mchip.learning.data.add_out [0]);
	assign \mchip.learning.data.w1_reg.D [1] = (_0163_ ? io_in[1] : \mchip.learning.data.add_out [1]);
	assign \mchip.learning.data.w1_reg.D [2] = (_0163_ ? io_in[2] : \mchip.learning.data.add_out [2]);
	assign \mchip.learning.data.w1_reg.D [3] = (_0163_ ? io_in[3] : \mchip.learning.data.add_out [3]);
	assign \mchip.learning.data.w1_reg.D [4] = (_0163_ ? io_in[4] : \mchip.learning.data.add_out [4]);
	assign \mchip.learning.data.w1_reg.D [5] = (_0163_ ? io_in[5] : \mchip.learning.data.add_out [5]);
	assign _0164_ = \mchip.learning.control.state [0] & io_in[10];
	assign \mchip.learning.data.w0_reg.D [0] = (_0164_ ? io_in[0] : \mchip.learning.data.add_out [0]);
	assign \mchip.learning.data.w0_reg.D [1] = (_0164_ ? io_in[1] : \mchip.learning.data.add_out [1]);
	assign \mchip.learning.data.w0_reg.D [2] = (_0164_ ? io_in[2] : \mchip.learning.data.add_out [2]);
	assign \mchip.learning.data.w0_reg.D [3] = (_0164_ ? io_in[3] : \mchip.learning.data.add_out [3]);
	assign \mchip.learning.data.w0_reg.D [4] = (_0164_ ? io_in[4] : \mchip.learning.data.add_out [4]);
	assign \mchip.learning.data.w0_reg.D [5] = (_0164_ ? io_in[5] : \mchip.learning.data.add_out [5]);
	assign _0165_ = _0164_ | _0051_;
	assign _0166_ = ~(\mchip.learning.control.state [4] | \mchip.learning.control.state [0]);
	assign \mchip.learning.control.en_w0  = _0165_ & ~_0166_;
	assign _0167_ = io_in[7] & io_in[6];
	assign _0168_ = (io_in[6] ? \mchip.learning.data.w0_reg.Q [4] : \mchip.learning.data.w0_reg.Q [2]);
	assign _0169_ = io_in[7] ^ io_in[6];
	assign _0170_ = (io_in[6] ? \mchip.learning.data.w0_reg.Q [0] : \mchip.learning.data.w1_reg.Q [4]);
	assign _0171_ = (_0169_ ? _0168_ : _0170_);
	assign _0172_ = io_in[7] & ~io_in[6];
	assign _0173_ = _0171_ & ~_0172_;
	assign _0174_ = (io_in[6] ? \mchip.learning.data.w1_reg.Q [2] : \mchip.learning.data.w1_reg.Q [0]);
	assign _0175_ = (io_in[6] ? \mchip.learning.data.w2_reg.Q [4] : \mchip.learning.data.w2_reg.Q [2]);
	assign _0176_ = (_0169_ ? _0174_ : _0175_);
	assign _0177_ = (io_in[6] ? \mchip.learning.data.w2_reg.Q [0] : \mchip.learning.data.add_reg.Q [4]);
	assign _0178_ = (io_in[6] ? \mchip.learning.data.add_reg.Q [2] : \mchip.learning.data.add_reg.Q [0]);
	assign _0179_ = (_0169_ ? _0177_ : _0178_);
	assign _0180_ = (_0172_ ? _0176_ : _0179_);
	assign io_out[0] = (_0167_ ? _0173_ : _0180_);
	assign _0181_ = (io_in[6] ? \mchip.learning.data.w0_reg.Q [5] : \mchip.learning.data.w0_reg.Q [3]);
	assign _0182_ = (io_in[6] ? \mchip.learning.data.w0_reg.Q [1] : \mchip.learning.data.w1_reg.Q [5]);
	assign _0183_ = (_0169_ ? _0181_ : _0182_);
	assign _0184_ = _0183_ & ~_0172_;
	assign _0185_ = (io_in[6] ? \mchip.learning.data.w1_reg.Q [3] : \mchip.learning.data.w1_reg.Q [1]);
	assign _0186_ = (io_in[6] ? \mchip.learning.data.w2_reg.Q [5] : \mchip.learning.data.w2_reg.Q [3]);
	assign _0187_ = (_0169_ ? _0185_ : _0186_);
	assign _0188_ = (io_in[6] ? \mchip.learning.data.w2_reg.Q [1] : \mchip.learning.data.add_reg.Q [5]);
	assign _0189_ = (io_in[6] ? \mchip.learning.data.add_reg.Q [3] : \mchip.learning.data.add_reg.Q [1]);
	assign _0190_ = (_0169_ ? _0188_ : _0189_);
	assign _0191_ = (_0172_ ? _0187_ : _0190_);
	assign io_out[1] = (_0167_ ? _0184_ : _0191_);
	assign _0192_ = \mchip.learning.data.w0_reg.Q [4] & ~io_in[6];
	assign _0193_ = (io_in[6] ? \mchip.learning.data.w0_reg.Q [2] : \mchip.learning.data.w0_reg.Q [0]);
	assign _0194_ = (_0169_ ? _0192_ : _0193_);
	assign _0195_ = _0194_ & ~_0172_;
	assign _0196_ = (io_in[6] ? \mchip.learning.data.w1_reg.Q [4] : \mchip.learning.data.w1_reg.Q [2]);
	assign _0197_ = (io_in[6] ? \mchip.learning.data.w1_reg.Q [0] : \mchip.learning.data.w2_reg.Q [4]);
	assign _0198_ = (_0169_ ? _0196_ : _0197_);
	assign _0199_ = (io_in[6] ? \mchip.learning.data.w2_reg.Q [2] : \mchip.learning.data.w2_reg.Q [0]);
	assign _0200_ = (io_in[6] ? \mchip.learning.data.add_reg.Q [4] : \mchip.learning.data.add_reg.Q [2]);
	assign _0201_ = (_0169_ ? _0199_ : _0200_);
	assign _0202_ = (_0172_ ? _0198_ : _0201_);
	assign io_out[2] = (_0167_ ? _0195_ : _0202_);
	assign _0203_ = \mchip.learning.data.w0_reg.Q [5] & ~io_in[6];
	assign _0204_ = (io_in[6] ? \mchip.learning.data.w0_reg.Q [3] : \mchip.learning.data.w0_reg.Q [1]);
	assign _0205_ = (_0169_ ? _0203_ : _0204_);
	assign _0206_ = _0205_ & ~_0172_;
	assign _0207_ = (io_in[6] ? \mchip.learning.data.w1_reg.Q [5] : \mchip.learning.data.w1_reg.Q [3]);
	assign _0208_ = (io_in[6] ? \mchip.learning.data.w1_reg.Q [1] : \mchip.learning.data.w2_reg.Q [5]);
	assign _0209_ = (_0169_ ? _0207_ : _0208_);
	assign _0210_ = (io_in[6] ? \mchip.learning.data.w2_reg.Q [3] : \mchip.learning.data.w2_reg.Q [1]);
	assign _0211_ = (io_in[6] ? \mchip.learning.data.add_reg.Q [5] : \mchip.learning.data.add_reg.Q [3]);
	assign _0212_ = (_0169_ ? _0210_ : _0211_);
	assign _0213_ = (_0172_ ? _0209_ : _0212_);
	assign io_out[3] = (_0167_ ? _0206_ : _0213_);
	assign _0214_ = ~_0172_;
	assign _0215_ = _0169_ | ~_0168_;
	assign _0216_ = _0214_ & ~_0215_;
	assign _0217_ = (_0169_ ? _0170_ : _0174_);
	assign _0218_ = (_0169_ ? _0175_ : _0177_);
	assign _0219_ = (_0172_ ? _0217_ : _0218_);
	assign io_out[4] = (_0167_ ? _0216_ : _0219_);
	assign _0220_ = _0169_ | ~_0181_;
	assign _0221_ = _0214_ & ~_0220_;
	assign _0222_ = (_0169_ ? _0182_ : _0185_);
	assign _0223_ = (_0169_ ? _0186_ : _0188_);
	assign _0224_ = (_0172_ ? _0222_ : _0223_);
	assign io_out[5] = (_0167_ ? _0221_ : _0224_);
	assign _0225_ = \mchip.learning.control.state [1] & ~_0023_;
	assign _0226_ = \mchip.learning.control.state [7] | \mchip.learning.control.state [5];
	assign _0227_ = _0226_ | _0225_;
	assign _0228_ = _0227_ | \mchip.learning.control.en_x2 ;
	assign _0229_ = ~\mchip.learning.control.state [8];
	assign _0230_ = _0226_ | \mchip.learning.control.state [1];
	assign _0231_ = _0229_ & ~_0230_;
	assign \mchip.learning.control.en_mult  = _0228_ & ~_0231_;
	assign _0232_ = _0041_ | \mchip.learning.control.en_x1 ;
	assign _0233_ = _0040_ & ~_0041_;
	assign \mchip.learning.control.en_add  = _0232_ & ~_0233_;
	assign _0234_ = _0047_ & \mchip.learning.control.state [4];
	assign _0235_ = _0234_ | _0079_;
	assign _0236_ = ~(\mchip.learning.control.state [4] | \mchip.learning.control.state [3]);
	assign \mchip.learning.control.en_w2  = _0235_ & ~_0236_;
	assign _0237_ = \mchip.learning.control.state [4] & ~_0045_;
	assign _0238_ = _0237_ | _0163_;
	assign _0239_ = ~(\mchip.learning.control.state [4] | \mchip.learning.control.state [6]);
	assign \mchip.learning.control.en_w1  = _0238_ & ~_0239_;
	assign _0240_ = \mchip.learning.control.state [10] & ~io_in[9];
	assign _0241_ = _0023_ & \mchip.learning.control.state [1];
	assign _0242_ = _0241_ | _0240_;
	assign _0243_ = ~(\mchip.learning.control.state [10] | \mchip.learning.control.state [1]);
	assign \mchip.learning.control.done  = _0242_ & ~_0243_;
	assign \mchip.learning.control.en_n  = \mchip.learning.control.state [9] & io_in[10];
	assign _0244_ = \mchip.learning.control.state [6] | \mchip.learning.control.state [3];
	assign _0245_ = \mchip.learning.control.state [0] | \mchip.learning.control.state [2];
	assign _0246_ = ~(_0245_ | _0244_);
	assign _0247_ = _0246_ & ~\mchip.learning.control.state [9];
	assign \mchip.learning.control.sync  = io_in[10] & ~_0247_;
	assign _0554_[1] = \mchip.learning.data.counter.count [1] ^ \mchip.learning.data.counter.count [0];
	assign _0248_ = _0225_ | \mchip.learning.control.en_x2 ;
	assign _0249_ = \mchip.learning.control.state [5] | \mchip.learning.control.state [1];
	assign _0250_ = _0229_ & ~_0249_;
	assign _0251_ = _0248_ & ~_0250_;
	assign _0252_ = ~(\mchip.learning.control.en_x2  | \mchip.learning.control.state [5]);
	assign _0253_ = _0252_ | _0250_;
	assign _0254_ = _0251_ & ~_0253_;
	assign _0255_ = \mchip.learning.data.w1_reg.Q [4] & ~_0251_;
	assign _0256_ = ~(_0253_ ^ _0251_);
	assign _0257_ = (_0251_ ? \mchip.learning.data.w1_reg.Q [2] : \mchip.learning.data.w1_reg.Q [0]);
	assign _0258_ = (_0256_ ? _0255_ : _0257_);
	assign _0259_ = ~(_0253_ | _0251_);
	assign _0260_ = _0258_ & ~_0259_;
	assign _0261_ = (_0251_ ? \mchip.learning.data.w2_reg.Q [4] : \mchip.learning.data.w2_reg.Q [2]);
	assign _0262_ = (_0251_ ? \mchip.learning.data.w2_reg.Q [0] : \mchip.learning.data.n_reg.Q [4]);
	assign _0263_ = (_0256_ ? _0261_ : _0262_);
	assign _0264_ = (_0251_ ? \mchip.learning.data.n_reg.Q [2] : \mchip.learning.data.n_reg.Q [0]);
	assign _0265_ = (_0251_ ? \mchip.learning.data.mult_reg.Q [4] : \mchip.learning.data.mult_reg.Q [2]);
	assign _0266_ = (_0256_ ? _0264_ : _0265_);
	assign _0267_ = (_0259_ ? _0263_ : _0266_);
	assign _0268_ = (_0254_ ? _0260_ : _0267_);
	assign _0269_ = ~_0268_;
	assign _0270_ = _0047_ | _0023_;
	assign _0271_ = _0270_ | ~\mchip.learning.control.state [1];
	assign _0272_ = _0271_ & ~\mchip.learning.control.en_x2 ;
	assign _0273_ = _0272_ | _0250_;
	assign _0274_ = _0046_ | _0023_;
	assign _0275_ = \mchip.learning.control.state [1] & ~_0274_;
	assign _0276_ = _0275_ | \mchip.learning.control.state [5];
	assign _0277_ = ~(_0276_ | \mchip.learning.control.en_x2 );
	assign _0278_ = ~(_0277_ | _0250_);
	assign _0279_ = _0278_ & ~_0273_;
	assign _0280_ = ~\mchip.learning.data.x1_reg.Q [2];
	assign _0281_ = ~\mchip.learning.data.x1_reg.Q [4];
	assign _0282_ = (_0273_ ? _0280_ : _0281_);
	assign _0283_ = _0277_ | _0250_;
	assign _0284_ = _0283_ ^ _0273_;
	assign _0285_ = ~\mchip.learning.data.x2_reg.Q [4];
	assign _0286_ = ~\mchip.learning.data.x1_reg.Q [0];
	assign _0287_ = (_0273_ ? _0285_ : _0286_);
	assign _0288_ = (_0284_ ? _0282_ : _0287_);
	assign _0289_ = _0273_ & ~_0283_;
	assign _0290_ = _0289_ | _0288_;
	assign _0291_ = ~\mchip.learning.data.x2_reg.Q [0];
	assign _0292_ = ~\mchip.learning.data.x2_reg.Q [2];
	assign _0293_ = (_0273_ ? _0291_ : _0292_);
	assign _0294_ = _0293_ | ~_0284_;
	assign _0295_ = _0278_ | _0273_;
	assign _0296_ = (_0289_ ? _0294_ : _0295_);
	assign _0297_ = (_0279_ ? _0290_ : _0296_);
	assign _0298_ = _0297_ | _0269_;
	assign _0299_ = ~\mchip.learning.data.w1_reg.Q [3];
	assign _0300_ = ~\mchip.learning.data.w1_reg.Q [5];
	assign _0301_ = (_0251_ ? _0300_ : _0299_);
	assign _0302_ = ~\mchip.learning.data.w2_reg.Q [5];
	assign _0303_ = ~\mchip.learning.data.w1_reg.Q [1];
	assign _0304_ = (_0251_ ? _0303_ : _0302_);
	assign _0305_ = (_0256_ ? _0301_ : _0304_);
	assign _0306_ = _0305_ | _0259_;
	assign _0307_ = ~\mchip.learning.data.w2_reg.Q [1];
	assign _0308_ = ~\mchip.learning.data.w2_reg.Q [3];
	assign _0309_ = (_0251_ ? _0308_ : _0307_);
	assign _0310_ = ~\mchip.learning.data.n_reg.Q [3];
	assign _0311_ = ~\mchip.learning.data.n_reg.Q [5];
	assign _0312_ = (_0251_ ? _0311_ : _0310_);
	assign _0313_ = (_0256_ ? _0309_ : _0312_);
	assign _0314_ = ~\mchip.learning.data.n_reg.Q [1];
	assign _0315_ = (_0251_ ? _0314_ : _0136_);
	assign _0316_ = ~\mchip.learning.data.mult_reg.Q [1];
	assign _0317_ = (_0251_ ? _0135_ : _0316_);
	assign _0318_ = (_0256_ ? _0315_ : _0317_);
	assign _0319_ = (_0259_ ? _0313_ : _0318_);
	assign _0320_ = (_0254_ ? _0306_ : _0319_);
	assign _0321_ = ~\mchip.learning.data.x1_reg.Q [3];
	assign _0322_ = ~\mchip.learning.data.x1_reg.Q [5];
	assign _0323_ = (_0273_ ? _0321_ : _0322_);
	assign _0324_ = ~\mchip.learning.data.x2_reg.Q [5];
	assign _0325_ = ~\mchip.learning.data.x1_reg.Q [1];
	assign _0326_ = (_0273_ ? _0324_ : _0325_);
	assign _0327_ = (_0284_ ? _0323_ : _0326_);
	assign _0328_ = _0327_ | _0289_;
	assign _0329_ = ~\mchip.learning.data.x2_reg.Q [1];
	assign _0330_ = ~\mchip.learning.data.x2_reg.Q [3];
	assign _0331_ = (_0273_ ? _0329_ : _0330_);
	assign _0332_ = _0331_ | ~_0284_;
	assign _0333_ = ~(_0273_ & _0020_);
	assign _0334_ = _0273_ | _0020_;
	assign _0335_ = (_0284_ ? _0333_ : _0334_);
	assign _0336_ = (_0289_ ? _0332_ : _0335_);
	assign _0337_ = (_0279_ ? _0328_ : _0336_);
	assign _0338_ = ~(_0337_ | _0320_);
	assign _0339_ = _0338_ ^ _0298_;
	assign _0340_ = ~\mchip.learning.data.w1_reg.Q [2];
	assign _0341_ = ~\mchip.learning.data.w1_reg.Q [4];
	assign _0342_ = (_0251_ ? _0341_ : _0340_);
	assign _0343_ = ~\mchip.learning.data.w2_reg.Q [4];
	assign _0344_ = ~\mchip.learning.data.w1_reg.Q [0];
	assign _0345_ = (_0251_ ? _0344_ : _0343_);
	assign _0346_ = (_0256_ ? _0342_ : _0345_);
	assign _0347_ = _0346_ | _0259_;
	assign _0348_ = ~\mchip.learning.data.w2_reg.Q [0];
	assign _0349_ = ~\mchip.learning.data.w2_reg.Q [2];
	assign _0350_ = (_0251_ ? _0349_ : _0348_);
	assign _0351_ = ~\mchip.learning.data.n_reg.Q [2];
	assign _0352_ = ~\mchip.learning.data.n_reg.Q [4];
	assign _0353_ = (_0251_ ? _0352_ : _0351_);
	assign _0354_ = (_0256_ ? _0350_ : _0353_);
	assign _0355_ = ~\mchip.learning.data.n_reg.Q [0];
	assign _0356_ = (_0251_ ? _0355_ : _0116_);
	assign _0357_ = (_0251_ ? _0074_ : _0073_);
	assign _0358_ = (_0256_ ? _0356_ : _0357_);
	assign _0359_ = (_0259_ ? _0354_ : _0358_);
	assign _0360_ = (_0254_ ? _0347_ : _0359_);
	assign _0361_ = _0360_ | _0337_;
	assign _0362_ = _0320_ | _0297_;
	assign _0363_ = _0362_ | _0361_;
	assign _0364_ = ~(_0363_ | _0339_);
	assign _0365_ = ~(_0273_ & \mchip.learning.data.x1_reg.Q [4]);
	assign _0366_ = (_0273_ ? _0286_ : _0280_);
	assign _0367_ = (_0284_ ? _0365_ : _0366_);
	assign _0368_ = _0367_ | _0289_;
	assign _0369_ = (_0273_ ? _0292_ : _0285_);
	assign _0370_ = _0273_ | _0291_;
	assign _0371_ = (_0284_ ? _0369_ : _0370_);
	assign _0372_ = _0371_ | ~_0289_;
	assign _0373_ = (_0279_ ? _0368_ : _0372_);
	assign _0374_ = ~(_0373_ | _0360_);
	assign _0375_ = ~(_0363_ ^ _0339_);
	assign _0376_ = _0374_ & ~_0375_;
	assign _0377_ = _0376_ | _0364_;
	assign _0378_ = ~(_0373_ | _0320_);
	assign _0379_ = _0338_ & ~_0298_;
	assign _0380_ = _0337_ | _0269_;
	assign _0381_ = _0251_ | _0300_;
	assign _0382_ = (_0251_ ? _0299_ : _0303_);
	assign _0383_ = (_0256_ ? _0381_ : _0382_);
	assign _0384_ = _0383_ | _0259_;
	assign _0385_ = (_0251_ ? _0302_ : _0308_);
	assign _0386_ = (_0251_ ? _0307_ : _0311_);
	assign _0387_ = (_0256_ ? _0385_ : _0386_);
	assign _0388_ = (_0251_ ? _0310_ : _0314_);
	assign _0389_ = (_0251_ ? _0136_ : _0135_);
	assign _0390_ = (_0256_ ? _0388_ : _0389_);
	assign _0391_ = (_0259_ ? _0387_ : _0390_);
	assign _0392_ = (_0254_ ? _0384_ : _0391_);
	assign _0393_ = ~(_0392_ | _0297_);
	assign _0394_ = ~(_0273_ & \mchip.learning.data.x1_reg.Q [5]);
	assign _0395_ = (_0273_ ? _0325_ : _0321_);
	assign _0396_ = (_0284_ ? _0394_ : _0395_);
	assign _0397_ = _0396_ | _0289_;
	assign _0398_ = (_0273_ ? _0330_ : _0324_);
	assign _0399_ = _0273_ | _0329_;
	assign _0400_ = (_0284_ ? _0398_ : _0399_);
	assign _0401_ = _0273_ ^ io_in[8];
	assign _0402_ = _0401_ | _0284_;
	assign _0403_ = (_0289_ ? _0400_ : _0402_);
	assign _0404_ = (_0279_ ? _0397_ : _0403_);
	assign _0405_ = _0404_ | _0360_;
	assign _0406_ = _0405_ ^ _0393_;
	assign _0407_ = ~(_0406_ ^ _0380_);
	assign _0408_ = _0407_ ^ _0379_;
	assign _0409_ = _0408_ ^ _0378_;
	assign \mchip.learning.data.mult.tmp [3] = ~(_0409_ ^ _0377_);
	assign _0410_ = _0377_ & ~_0409_;
	assign _0411_ = _0408_ | ~_0378_;
	assign _0412_ = _0379_ & ~_0407_;
	assign _0413_ = _0411_ & ~_0412_;
	assign _0414_ = _0406_ | _0380_;
	assign _0415_ = _0393_ & ~_0405_;
	assign _0416_ = _0414_ & ~_0415_;
	assign _0417_ = _0342_ | _0256_;
	assign _0418_ = _0417_ | _0259_;
	assign _0419_ = (_0256_ ? _0345_ : _0350_);
	assign _0420_ = (_0256_ ? _0353_ : _0356_);
	assign _0421_ = (_0259_ ? _0419_ : _0420_);
	assign _0422_ = (_0254_ ? _0418_ : _0421_);
	assign _0423_ = ~(_0422_ | _0297_);
	assign _0424_ = ~(_0404_ | _0320_);
	assign _0425_ = _0424_ ^ _0423_;
	assign _0426_ = _0392_ | _0337_;
	assign _0427_ = _0426_ ^ _0425_;
	assign _0428_ = _0427_ ^ _0416_;
	assign _0429_ = _0284_ | _0282_;
	assign _0430_ = _0429_ | _0289_;
	assign _0431_ = ~_0279_;
	assign _0432_ = (_0284_ ? _0287_ : _0293_);
	assign _0433_ = (_0289_ ? _0432_ : _0431_);
	assign _0434_ = (_0279_ ? _0430_ : _0433_);
	assign _0435_ = _0434_ | _0360_;
	assign _0436_ = _0268_ & ~_0373_;
	assign _0437_ = _0436_ ^ _0435_;
	assign _0438_ = ~(_0437_ ^ _0428_);
	assign _0439_ = _0438_ ^ _0413_;
	assign _0440_ = _0410_ & ~_0439_;
	assign _0441_ = _0438_ & ~_0413_;
	assign _0442_ = _0436_ & ~_0435_;
	assign _0443_ = _0427_ | _0416_;
	assign _0444_ = _0428_ & ~_0437_;
	assign _0445_ = _0444_ | ~_0443_;
	assign _0446_ = _0323_ | _0284_;
	assign _0447_ = _0446_ | _0289_;
	assign _0448_ = (_0284_ ? _0326_ : _0331_);
	assign _0449_ = _0333_ | _0284_;
	assign _0450_ = (_0289_ ? _0448_ : _0449_);
	assign _0451_ = (_0279_ ? _0447_ : _0450_);
	assign _0452_ = ~(_0451_ | _0360_);
	assign _0453_ = _0434_ | _0320_;
	assign _0454_ = ~(_0392_ | _0373_);
	assign _0455_ = _0454_ ^ _0453_;
	assign _0456_ = ~(_0455_ ^ _0452_);
	assign _0457_ = ~(_0424_ & _0423_);
	assign _0458_ = _0425_ & ~_0426_;
	assign _0459_ = _0458_ | ~_0457_;
	assign _0460_ = ~(_0422_ | _0337_);
	assign _0461_ = _0301_ | _0256_;
	assign _0462_ = _0461_ | _0259_;
	assign _0463_ = (_0256_ ? _0304_ : _0309_);
	assign _0464_ = (_0256_ ? _0312_ : _0315_);
	assign _0465_ = (_0259_ ? _0463_ : _0464_);
	assign _0466_ = (_0254_ ? _0462_ : _0465_);
	assign _0467_ = ~(_0466_ | _0297_);
	assign _0468_ = _0404_ | _0269_;
	assign _0469_ = _0468_ ^ _0467_;
	assign _0470_ = _0469_ ^ _0460_;
	assign _0471_ = _0470_ ^ _0459_;
	assign _0472_ = _0471_ ^ _0456_;
	assign _0473_ = _0472_ ^ _0445_;
	assign _0474_ = _0473_ ^ _0442_;
	assign _0475_ = _0474_ ^ _0441_;
	assign \mchip.learning.data.mult.tmp [5] = ~(_0475_ ^ _0440_);
	assign _0476_ = _0440_ & ~_0475_;
	assign _0477_ = _0441_ & ~_0474_;
	assign _0478_ = _0477_ | _0476_;
	assign _0479_ = _0442_ & ~_0473_;
	assign _0480_ = _0445_ & ~_0472_;
	assign _0481_ = _0480_ | _0479_;
	assign _0482_ = _0452_ & ~_0455_;
	assign _0483_ = _0454_ & ~_0453_;
	assign _0484_ = _0483_ | _0482_;
	assign _0485_ = _0471_ | ~_0456_;
	assign _0486_ = _0459_ & ~_0470_;
	assign _0487_ = _0486_ | ~_0485_;
	assign _0488_ = ~(_0451_ | _0320_);
	assign _0489_ = _0268_ & ~_0434_;
	assign _0490_ = ~(_0422_ | _0373_);
	assign _0491_ = _0490_ ^ _0489_;
	assign _0492_ = _0491_ ^ _0488_;
	assign _0493_ = _0469_ | ~_0460_;
	assign _0494_ = _0467_ & ~_0468_;
	assign _0495_ = _0494_ | ~_0493_;
	assign _0496_ = _0466_ | _0337_;
	assign _0497_ = ~(_0404_ | _0392_);
	assign _0498_ = _0497_ ^ _0496_;
	assign _0499_ = _0498_ ^ _0495_;
	assign _0500_ = _0499_ ^ _0492_;
	assign _0501_ = _0500_ ^ _0487_;
	assign _0502_ = ~(_0501_ ^ _0484_);
	assign _0503_ = ~(_0502_ ^ _0481_);
	assign \mchip.learning.data.mult.tmp [6] = ~(_0503_ ^ _0478_);
	assign _0504_ = _0502_ & _0481_;
	assign _0505_ = _0478_ & ~_0503_;
	assign _0506_ = ~(_0505_ | _0504_);
	assign _0507_ = _0484_ & ~_0501_;
	assign _0508_ = _0487_ & ~_0500_;
	assign _0509_ = _0508_ | _0507_;
	assign _0510_ = ~(_0490_ & _0489_);
	assign _0511_ = _0491_ & _0488_;
	assign _0512_ = _0510_ & ~_0511_;
	assign _0513_ = _0499_ | ~_0492_;
	assign _0514_ = _0495_ & ~_0498_;
	assign _0515_ = _0514_ | ~_0513_;
	assign _0516_ = _0268_ & ~_0451_;
	assign _0517_ = _0434_ | _0392_;
	assign _0518_ = ~(_0466_ | _0373_);
	assign _0519_ = ~(_0518_ ^ _0517_);
	assign _0520_ = ~(_0519_ ^ _0516_);
	assign _0521_ = _0496_ | ~_0497_;
	assign _0522_ = ~(_0422_ | _0404_);
	assign _0523_ = _0522_ ^ _0521_;
	assign _0524_ = _0523_ ^ _0520_;
	assign _0525_ = ~_0524_;
	assign _0526_ = _0525_ ^ _0515_;
	assign _0527_ = _0526_ ^ _0512_;
	assign _0528_ = ~(_0527_ ^ _0509_);
	assign \mchip.learning.data.mult.tmp [7] = _0528_ ^ _0506_;
	assign _0529_ = _0527_ & _0509_;
	assign _0530_ = _0504_ & ~_0528_;
	assign _0531_ = _0530_ | _0529_;
	assign _0532_ = _0528_ | _0503_;
	assign _0533_ = _0478_ & ~_0532_;
	assign _0534_ = _0533_ | _0531_;
	assign _0535_ = _0526_ | _0512_;
	assign _0536_ = _0515_ & ~_0525_;
	assign _0537_ = _0535_ & ~_0536_;
	assign _0538_ = _0517_ | ~_0518_;
	assign _0539_ = _0519_ & _0516_;
	assign _0540_ = _0538_ & ~_0539_;
	assign _0541_ = _0523_ | _0520_;
	assign _0542_ = _0522_ & ~_0521_;
	assign _0543_ = _0541_ & ~_0542_;
	assign _0544_ = _0451_ | _0392_;
	assign _0545_ = ~(_0434_ | _0422_);
	assign _0546_ = _0545_ ^ _0544_;
	assign _0547_ = ~(_0466_ | _0404_);
	assign _0548_ = _0547_ ^ _0546_;
	assign _0549_ = _0548_ ^ _0543_;
	assign _0550_ = _0549_ ^ _0540_;
	assign _0551_ = _0550_ ^ _0537_;
	assign \mchip.learning.data.mult.tmp [8] = _0551_ ^ _0534_;
	assign \mchip.learning.data.mult.tmp [4] = ~(_0439_ ^ _0410_);
	assign _0003_ = \mchip.learning.control.state [5] & ~io_in[13];
	assign _0552_ = _0023_ | io_in[13];
	assign _0002_ = \mchip.learning.control.state [1] & ~_0552_;
	assign _0001_ = \mchip.learning.control.state [8] & ~_0017_;
	assign _0000_ = \mchip.learning.control.state [7] & ~io_in[13];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.learning.data.add_reg.Q [0] <= 1'h0;
		else if (\mchip.learning.control.en_add )
			\mchip.learning.data.add_reg.Q [0] <= \mchip.learning.data.add_out [0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.learning.data.add_reg.Q [1] <= 1'h0;
		else if (\mchip.learning.control.en_add )
			\mchip.learning.data.add_reg.Q [1] <= \mchip.learning.data.add_out [1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.learning.data.add_reg.Q [2] <= 1'h0;
		else if (\mchip.learning.control.en_add )
			\mchip.learning.data.add_reg.Q [2] <= \mchip.learning.data.add_out [2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.learning.data.add_reg.Q [3] <= 1'h0;
		else if (\mchip.learning.control.en_add )
			\mchip.learning.data.add_reg.Q [3] <= \mchip.learning.data.add_out [3];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.learning.data.add_reg.Q [4] <= 1'h0;
		else if (\mchip.learning.control.en_add )
			\mchip.learning.data.add_reg.Q [4] <= \mchip.learning.data.add_out [4];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.learning.data.add_reg.Q [5] <= 1'h0;
		else if (\mchip.learning.control.en_add )
			\mchip.learning.data.add_reg.Q [5] <= \mchip.learning.data.add_out [5];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.learning.data.mult_reg.Q [0] <= 1'h0;
		else if (\mchip.learning.control.en_mult )
			\mchip.learning.data.mult_reg.Q [0] <= \mchip.learning.data.mult.tmp [3];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.learning.data.mult_reg.Q [1] <= 1'h0;
		else if (\mchip.learning.control.en_mult )
			\mchip.learning.data.mult_reg.Q [1] <= \mchip.learning.data.mult.tmp [4];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.learning.data.mult_reg.Q [2] <= 1'h0;
		else if (\mchip.learning.control.en_mult )
			\mchip.learning.data.mult_reg.Q [2] <= \mchip.learning.data.mult.tmp [5];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.learning.data.mult_reg.Q [3] <= 1'h0;
		else if (\mchip.learning.control.en_mult )
			\mchip.learning.data.mult_reg.Q [3] <= \mchip.learning.data.mult.tmp [6];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.learning.data.mult_reg.Q [4] <= 1'h0;
		else if (\mchip.learning.control.en_mult )
			\mchip.learning.data.mult_reg.Q [4] <= \mchip.learning.data.mult.tmp [7];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.learning.data.mult_reg.Q [5] <= 1'h0;
		else if (\mchip.learning.control.en_mult )
			\mchip.learning.data.mult_reg.Q [5] <= \mchip.learning.data.mult.tmp [8];
	always @(posedge io_in[12])
		if (_0011_)
			\mchip.learning.data.counter.count [0] <= 1'h0;
		else if (\mchip.learning.control.state [4])
			\mchip.learning.data.counter.count [0] <= _0553_[0];
	always @(posedge io_in[12])
		if (_0011_)
			\mchip.learning.data.counter.count [1] <= 1'h0;
		else if (\mchip.learning.control.state [4])
			\mchip.learning.data.counter.count [1] <= _0554_[1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.learning.data.x2_reg.Q [0] <= 1'h0;
		else if (\mchip.learning.control.en_x2 )
			\mchip.learning.data.x2_reg.Q [0] <= io_in[0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.learning.data.x2_reg.Q [1] <= 1'h0;
		else if (\mchip.learning.control.en_x2 )
			\mchip.learning.data.x2_reg.Q [1] <= io_in[1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.learning.data.x2_reg.Q [2] <= 1'h0;
		else if (\mchip.learning.control.en_x2 )
			\mchip.learning.data.x2_reg.Q [2] <= io_in[2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.learning.data.x2_reg.Q [3] <= 1'h0;
		else if (\mchip.learning.control.en_x2 )
			\mchip.learning.data.x2_reg.Q [3] <= io_in[3];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.learning.data.x2_reg.Q [4] <= 1'h0;
		else if (\mchip.learning.control.en_x2 )
			\mchip.learning.data.x2_reg.Q [4] <= io_in[4];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.learning.data.x2_reg.Q [5] <= 1'h0;
		else if (\mchip.learning.control.en_x2 )
			\mchip.learning.data.x2_reg.Q [5] <= io_in[5];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.learning.data.x1_reg.Q [0] <= 1'h0;
		else if (\mchip.learning.control.en_x1 )
			\mchip.learning.data.x1_reg.Q [0] <= io_in[0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.learning.data.x1_reg.Q [1] <= 1'h0;
		else if (\mchip.learning.control.en_x1 )
			\mchip.learning.data.x1_reg.Q [1] <= io_in[1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.learning.data.x1_reg.Q [2] <= 1'h0;
		else if (\mchip.learning.control.en_x1 )
			\mchip.learning.data.x1_reg.Q [2] <= io_in[2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.learning.data.x1_reg.Q [3] <= 1'h0;
		else if (\mchip.learning.control.en_x1 )
			\mchip.learning.data.x1_reg.Q [3] <= io_in[3];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.learning.data.x1_reg.Q [4] <= 1'h0;
		else if (\mchip.learning.control.en_x1 )
			\mchip.learning.data.x1_reg.Q [4] <= io_in[4];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.learning.data.x1_reg.Q [5] <= 1'h0;
		else if (\mchip.learning.control.en_x1 )
			\mchip.learning.data.x1_reg.Q [5] <= io_in[5];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.learning.data.n_reg.Q [0] <= 1'h0;
		else if (\mchip.learning.control.en_n )
			\mchip.learning.data.n_reg.Q [0] <= io_in[0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.learning.data.n_reg.Q [1] <= 1'h0;
		else if (\mchip.learning.control.en_n )
			\mchip.learning.data.n_reg.Q [1] <= io_in[1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.learning.data.n_reg.Q [2] <= 1'h0;
		else if (\mchip.learning.control.en_n )
			\mchip.learning.data.n_reg.Q [2] <= io_in[2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.learning.data.n_reg.Q [3] <= 1'h0;
		else if (\mchip.learning.control.en_n )
			\mchip.learning.data.n_reg.Q [3] <= io_in[3];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.learning.data.n_reg.Q [4] <= 1'h0;
		else if (\mchip.learning.control.en_n )
			\mchip.learning.data.n_reg.Q [4] <= io_in[4];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.learning.data.n_reg.Q [5] <= 1'h0;
		else if (\mchip.learning.control.en_n )
			\mchip.learning.data.n_reg.Q [5] <= io_in[5];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.learning.data.w2_reg.Q [0] <= 1'h0;
		else if (\mchip.learning.control.en_w2 )
			\mchip.learning.data.w2_reg.Q [0] <= \mchip.learning.data.w2_reg.D [0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.learning.data.w2_reg.Q [1] <= 1'h0;
		else if (\mchip.learning.control.en_w2 )
			\mchip.learning.data.w2_reg.Q [1] <= \mchip.learning.data.w2_reg.D [1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.learning.data.w2_reg.Q [2] <= 1'h0;
		else if (\mchip.learning.control.en_w2 )
			\mchip.learning.data.w2_reg.Q [2] <= \mchip.learning.data.w2_reg.D [2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.learning.data.w2_reg.Q [3] <= 1'h0;
		else if (\mchip.learning.control.en_w2 )
			\mchip.learning.data.w2_reg.Q [3] <= \mchip.learning.data.w2_reg.D [3];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.learning.data.w2_reg.Q [4] <= 1'h0;
		else if (\mchip.learning.control.en_w2 )
			\mchip.learning.data.w2_reg.Q [4] <= \mchip.learning.data.w2_reg.D [4];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.learning.data.w2_reg.Q [5] <= 1'h0;
		else if (\mchip.learning.control.en_w2 )
			\mchip.learning.data.w2_reg.Q [5] <= \mchip.learning.data.w2_reg.D [5];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.learning.data.w1_reg.Q [0] <= 1'h0;
		else if (\mchip.learning.control.en_w1 )
			\mchip.learning.data.w1_reg.Q [0] <= \mchip.learning.data.w1_reg.D [0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.learning.data.w1_reg.Q [1] <= 1'h0;
		else if (\mchip.learning.control.en_w1 )
			\mchip.learning.data.w1_reg.Q [1] <= \mchip.learning.data.w1_reg.D [1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.learning.data.w1_reg.Q [2] <= 1'h0;
		else if (\mchip.learning.control.en_w1 )
			\mchip.learning.data.w1_reg.Q [2] <= \mchip.learning.data.w1_reg.D [2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.learning.data.w1_reg.Q [3] <= 1'h0;
		else if (\mchip.learning.control.en_w1 )
			\mchip.learning.data.w1_reg.Q [3] <= \mchip.learning.data.w1_reg.D [3];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.learning.data.w1_reg.Q [4] <= 1'h0;
		else if (\mchip.learning.control.en_w1 )
			\mchip.learning.data.w1_reg.Q [4] <= \mchip.learning.data.w1_reg.D [4];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.learning.data.w1_reg.Q [5] <= 1'h0;
		else if (\mchip.learning.control.en_w1 )
			\mchip.learning.data.w1_reg.Q [5] <= \mchip.learning.data.w1_reg.D [5];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.learning.data.w0_reg.Q [0] <= 1'h0;
		else if (\mchip.learning.control.en_w0 )
			\mchip.learning.data.w0_reg.Q [0] <= \mchip.learning.data.w0_reg.D [0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.learning.data.w0_reg.Q [1] <= 1'h0;
		else if (\mchip.learning.control.en_w0 )
			\mchip.learning.data.w0_reg.Q [1] <= \mchip.learning.data.w0_reg.D [1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.learning.data.w0_reg.Q [2] <= 1'h0;
		else if (\mchip.learning.control.en_w0 )
			\mchip.learning.data.w0_reg.Q [2] <= \mchip.learning.data.w0_reg.D [2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.learning.data.w0_reg.Q [3] <= 1'h0;
		else if (\mchip.learning.control.en_w0 )
			\mchip.learning.data.w0_reg.Q [3] <= \mchip.learning.data.w0_reg.D [3];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.learning.data.w0_reg.Q [4] <= 1'h0;
		else if (\mchip.learning.control.en_w0 )
			\mchip.learning.data.w0_reg.Q [4] <= \mchip.learning.data.w0_reg.D [4];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.learning.data.w0_reg.Q [5] <= 1'h0;
		else if (\mchip.learning.control.en_w0 )
			\mchip.learning.data.w0_reg.Q [5] <= \mchip.learning.data.w0_reg.D [5];
	always @(posedge io_in[12]) \mchip.learning.control.state [0] <= _0004_;
	always @(posedge io_in[12]) \mchip.learning.control.state [1] <= _0005_;
	always @(posedge io_in[12]) \mchip.learning.control.state [2] <= _0006_;
	always @(posedge io_in[12]) \mchip.learning.control.state [3] <= _0007_;
	always @(posedge io_in[12]) \mchip.learning.control.state [4] <= _0000_;
	always @(posedge io_in[12]) \mchip.learning.control.state [5] <= _0001_;
	always @(posedge io_in[12]) \mchip.learning.control.state [6] <= _0008_;
	always @(posedge io_in[12]) \mchip.learning.control.state [7] <= _0002_;
	always @(posedge io_in[12]) \mchip.learning.control.state [8] <= _0009_;
	always @(posedge io_in[12]) \mchip.learning.control.state [9] <= _0010_;
	always @(posedge io_in[12]) \mchip.learning.control.state [10] <= _0003_;
	assign _0553_[1] = 1'h0;
	assign _0554_[0] = _0553_[0];
	assign io_out[13:6] = {5'h00, \mchip.learning.control.done , \mchip.learning.classification , \mchip.learning.control.sync };
	assign \mchip.clock  = io_in[12];
	assign \mchip.io_in  = io_in[11:0];
	assign \mchip.io_out  = {3'h0, \mchip.learning.control.done , \mchip.learning.classification , \mchip.learning.control.sync , io_out[5:0]};
	assign \mchip.learning.clk  = io_in[12];
	assign \mchip.learning.control.classification  = \mchip.learning.classification ;
	assign \mchip.learning.control.clk  = io_in[12];
	assign \mchip.learning.control.correct  = io_in[8];
	assign \mchip.learning.control.count  = \mchip.learning.data.counter.count ;
	assign \mchip.learning.control.en_count  = \mchip.learning.control.state [4];
	assign \mchip.learning.control.go  = io_in[10];
	assign \mchip.learning.control.sel_add_A  = \mchip.learning.control.en_x1 ;
	assign \mchip.learning.control.update  = io_in[9];
	assign \mchip.learning.correct  = io_in[8];
	assign \mchip.learning.count  = \mchip.learning.data.counter.count ;
	assign \mchip.learning.data.add.cin  = 1'h0;
	assign \mchip.learning.data.add.sum  = \mchip.learning.data.add_out ;
	assign \mchip.learning.data.add_A_mux.in  = {6'h00, \mchip.learning.data.mult_reg.Q };
	assign \mchip.learning.data.add_A_mux.sel  = \mchip.learning.control.en_x1 ;
	assign \mchip.learning.data.add_B_mux.in  = {\mchip.learning.data.w0_reg.Q , \mchip.learning.data.add_reg.Q , \mchip.learning.data.w1_reg.Q , \mchip.learning.data.w2_reg.Q };
	assign \mchip.learning.data.add_out_reg  = \mchip.learning.data.add_reg.Q ;
	assign \mchip.learning.data.add_reg.D  = \mchip.learning.data.add_out ;
	assign \mchip.learning.data.add_reg.clk  = io_in[12];
	assign \mchip.learning.data.add_reg.en  = \mchip.learning.control.en_add ;
	assign \mchip.learning.data.classification  = \mchip.learning.classification ;
	assign \mchip.learning.data.clk  = io_in[12];
	assign \mchip.learning.data.correct  = io_in[8];
	assign \mchip.learning.data.count  = \mchip.learning.data.counter.count ;
	assign \mchip.learning.data.counter.clk  = io_in[12];
	assign \mchip.learning.data.counter.en  = \mchip.learning.control.state [4];
	assign \mchip.learning.data.d  = {2'h0, io_in[8], 3'h0};
	assign \mchip.learning.data.en_add  = \mchip.learning.control.en_add ;
	assign \mchip.learning.data.en_count  = \mchip.learning.control.state [4];
	assign \mchip.learning.data.en_mult  = \mchip.learning.control.en_mult ;
	assign \mchip.learning.data.en_n  = \mchip.learning.control.en_n ;
	assign \mchip.learning.data.en_w0  = \mchip.learning.control.en_w0 ;
	assign \mchip.learning.data.en_w1  = \mchip.learning.control.en_w1 ;
	assign \mchip.learning.data.en_w2  = \mchip.learning.control.en_w2 ;
	assign \mchip.learning.data.en_x1  = \mchip.learning.control.en_x1 ;
	assign \mchip.learning.data.en_x2  = \mchip.learning.control.en_x2 ;
	assign \mchip.learning.data.in_val  = io_in[5:0];
	assign \mchip.learning.data.input_mux.in  = {\mchip.learning.data.w0_reg.Q , \mchip.learning.data.w1_reg.Q , \mchip.learning.data.w2_reg.Q , \mchip.learning.data.add_reg.Q };
	assign \mchip.learning.data.input_mux.out  = io_out[5:0];
	assign \mchip.learning.data.input_mux.sel  = io_in[7:6];
	assign \mchip.learning.data.mult.M  = \mchip.learning.data.mult.tmp [8:3];
	assign {\mchip.learning.data.mult.tmp [11:9], \mchip.learning.data.mult.tmp [2:0]} = 6'h00;
	assign \mchip.learning.data.mult_A_mux.in  = {\mchip.learning.data.w1_reg.Q , \mchip.learning.data.w2_reg.Q , \mchip.learning.data.n_reg.Q , \mchip.learning.data.mult_reg.Q };
	assign \mchip.learning.data.mult_B_mux.in  = {\mchip.learning.data.x1_reg.Q , \mchip.learning.data.x2_reg.Q , 8'h04, io_in[8], 3'h0};
	assign \mchip.learning.data.mult_out  = \mchip.learning.data.mult.tmp [8:3];
	assign \mchip.learning.data.mult_out_reg  = \mchip.learning.data.mult_reg.Q ;
	assign \mchip.learning.data.mult_reg.D  = \mchip.learning.data.mult.tmp [8:3];
	assign \mchip.learning.data.mult_reg.clk  = io_in[12];
	assign \mchip.learning.data.mult_reg.en  = \mchip.learning.control.en_mult ;
	assign \mchip.learning.data.n  = \mchip.learning.data.n_reg.Q ;
	assign \mchip.learning.data.n_reg.D  = io_in[5:0];
	assign \mchip.learning.data.n_reg.clk  = io_in[12];
	assign \mchip.learning.data.n_reg.en  = \mchip.learning.control.en_n ;
	assign \mchip.learning.data.out_val  = io_out[5:0];
	assign \mchip.learning.data.sel_add_A  = \mchip.learning.control.en_x1 ;
	assign \mchip.learning.data.sel_out  = io_in[7:6];
	assign \mchip.learning.data.w0  = \mchip.learning.data.w0_reg.Q ;
	assign \mchip.learning.data.w0_reg.clk  = io_in[12];
	assign \mchip.learning.data.w0_reg.en  = \mchip.learning.control.en_w0 ;
	assign \mchip.learning.data.w1  = \mchip.learning.data.w1_reg.Q ;
	assign \mchip.learning.data.w1_reg.clk  = io_in[12];
	assign \mchip.learning.data.w1_reg.en  = \mchip.learning.control.en_w1 ;
	assign \mchip.learning.data.w2  = \mchip.learning.data.w2_reg.Q ;
	assign \mchip.learning.data.w2_reg.clk  = io_in[12];
	assign \mchip.learning.data.w2_reg.en  = \mchip.learning.control.en_w2 ;
	assign \mchip.learning.data.x1  = \mchip.learning.data.x1_reg.Q ;
	assign \mchip.learning.data.x1_reg.D  = io_in[5:0];
	assign \mchip.learning.data.x1_reg.clk  = io_in[12];
	assign \mchip.learning.data.x1_reg.en  = \mchip.learning.control.en_x1 ;
	assign \mchip.learning.data.x2  = \mchip.learning.data.x2_reg.Q ;
	assign \mchip.learning.data.x2_reg.D  = io_in[5:0];
	assign \mchip.learning.data.x2_reg.clk  = io_in[12];
	assign \mchip.learning.data.x2_reg.en  = \mchip.learning.control.en_x2 ;
	assign \mchip.learning.done  = \mchip.learning.control.done ;
	assign \mchip.learning.en_add  = \mchip.learning.control.en_add ;
	assign \mchip.learning.en_count  = \mchip.learning.control.state [4];
	assign \mchip.learning.en_mult  = \mchip.learning.control.en_mult ;
	assign \mchip.learning.en_n  = \mchip.learning.control.en_n ;
	assign \mchip.learning.en_w0  = \mchip.learning.control.en_w0 ;
	assign \mchip.learning.en_w1  = \mchip.learning.control.en_w1 ;
	assign \mchip.learning.en_w2  = \mchip.learning.control.en_w2 ;
	assign \mchip.learning.en_x1  = \mchip.learning.control.en_x1 ;
	assign \mchip.learning.en_x2  = \mchip.learning.control.en_x2 ;
	assign \mchip.learning.go  = io_in[10];
	assign \mchip.learning.in_val  = io_in[5:0];
	assign \mchip.learning.out_val  = io_out[5:0];
	assign \mchip.learning.sel_add_A  = \mchip.learning.control.en_x1 ;
	assign \mchip.learning.sel_out  = io_in[7:6];
	assign \mchip.learning.sync  = \mchip.learning.control.sync ;
	assign \mchip.learning.update  = io_in[9];
	assign \mchip.reset  = io_in[13];
endmodule
module d27_svemulap_fpu (
	io_in,
	io_out
);
	wire _0000_;
	wire _0001_;
	wire _0002_;
	wire _0003_;
	wire _0004_;
	wire _0005_;
	wire _0006_;
	wire _0007_;
	wire _0008_;
	wire _0009_;
	wire _0010_;
	wire _0011_;
	wire _0012_;
	wire _0013_;
	wire _0014_;
	wire _0015_;
	wire _0016_;
	wire _0017_;
	wire _0018_;
	wire _0019_;
	wire _0020_;
	wire _0021_;
	wire _0022_;
	wire _0023_;
	wire _0024_;
	wire _0025_;
	wire _0026_;
	wire _0027_;
	wire _0028_;
	wire _0029_;
	wire _0030_;
	wire _0031_;
	wire _0032_;
	wire _0033_;
	wire _0034_;
	wire _0035_;
	wire _0036_;
	wire _0037_;
	wire _0038_;
	wire _0039_;
	wire _0040_;
	wire _0041_;
	wire _0042_;
	wire _0043_;
	wire _0044_;
	wire _0045_;
	wire _0046_;
	wire _0047_;
	wire _0048_;
	wire _0049_;
	wire _0050_;
	wire _0051_;
	wire _0052_;
	wire _0053_;
	wire _0054_;
	wire _0055_;
	wire _0056_;
	wire _0057_;
	wire _0058_;
	wire _0059_;
	wire _0060_;
	wire _0061_;
	wire _0062_;
	wire _0063_;
	wire _0064_;
	wire _0065_;
	wire _0066_;
	wire _0067_;
	wire _0068_;
	wire _0069_;
	wire _0070_;
	wire _0071_;
	wire _0072_;
	wire _0073_;
	wire _0074_;
	wire _0075_;
	wire _0076_;
	wire _0077_;
	wire _0078_;
	wire _0079_;
	wire _0080_;
	wire _0081_;
	wire _0082_;
	wire _0083_;
	wire _0084_;
	wire _0085_;
	wire _0086_;
	wire _0087_;
	wire _0088_;
	wire _0089_;
	wire _0090_;
	wire _0091_;
	wire _0092_;
	wire _0093_;
	wire _0094_;
	wire _0095_;
	wire _0096_;
	wire _0097_;
	wire _0098_;
	wire _0099_;
	wire _0100_;
	wire _0101_;
	wire _0102_;
	wire _0103_;
	wire _0104_;
	wire _0105_;
	wire _0106_;
	wire _0107_;
	wire _0108_;
	wire _0109_;
	wire _0110_;
	wire _0111_;
	wire _0112_;
	wire _0113_;
	wire _0114_;
	wire _0115_;
	wire _0116_;
	wire _0117_;
	wire _0118_;
	wire _0119_;
	wire _0120_;
	wire _0121_;
	wire _0122_;
	wire _0123_;
	wire _0124_;
	wire _0125_;
	wire _0126_;
	wire _0127_;
	wire _0128_;
	wire _0129_;
	wire _0130_;
	wire _0131_;
	wire _0132_;
	wire _0133_;
	wire _0134_;
	wire _0135_;
	wire _0136_;
	wire _0137_;
	wire _0138_;
	wire _0139_;
	wire _0140_;
	wire _0141_;
	wire _0142_;
	wire _0143_;
	wire _0144_;
	wire _0145_;
	wire _0146_;
	wire _0147_;
	wire _0148_;
	wire _0149_;
	wire _0150_;
	wire _0151_;
	wire _0152_;
	wire _0153_;
	wire _0154_;
	wire _0155_;
	wire _0156_;
	wire _0157_;
	wire _0158_;
	wire _0159_;
	wire _0160_;
	wire _0161_;
	wire _0162_;
	wire _0163_;
	wire _0164_;
	wire _0165_;
	wire _0166_;
	wire _0167_;
	wire _0168_;
	wire _0169_;
	wire _0170_;
	wire _0171_;
	wire _0172_;
	wire _0173_;
	wire _0174_;
	wire _0175_;
	wire _0176_;
	wire _0177_;
	wire _0178_;
	wire _0179_;
	wire _0180_;
	wire _0181_;
	wire _0182_;
	wire _0183_;
	wire _0184_;
	wire _0185_;
	wire _0186_;
	wire _0187_;
	wire _0188_;
	wire _0189_;
	wire _0190_;
	wire _0191_;
	wire _0192_;
	wire _0193_;
	wire _0194_;
	wire _0195_;
	wire _0196_;
	wire _0197_;
	wire _0198_;
	wire _0199_;
	wire _0200_;
	wire _0201_;
	wire _0202_;
	wire _0203_;
	wire _0204_;
	wire _0205_;
	wire _0206_;
	wire _0207_;
	wire _0208_;
	wire _0209_;
	wire _0210_;
	wire _0211_;
	wire _0212_;
	wire _0213_;
	wire _0214_;
	wire _0215_;
	wire _0216_;
	wire _0217_;
	wire _0218_;
	wire _0219_;
	wire _0220_;
	wire _0221_;
	wire _0222_;
	wire _0223_;
	wire _0224_;
	wire _0225_;
	wire _0226_;
	wire _0227_;
	wire _0228_;
	wire _0229_;
	wire _0230_;
	wire _0231_;
	wire _0232_;
	wire _0233_;
	wire _0234_;
	wire _0235_;
	wire _0236_;
	wire _0237_;
	wire _0238_;
	wire _0239_;
	wire _0240_;
	wire _0241_;
	wire _0242_;
	wire _0243_;
	wire _0244_;
	wire _0245_;
	wire _0246_;
	wire _0247_;
	wire _0248_;
	wire _0249_;
	wire _0250_;
	wire _0251_;
	wire _0252_;
	wire _0253_;
	wire _0254_;
	wire _0255_;
	wire _0256_;
	wire _0257_;
	wire _0258_;
	wire _0259_;
	wire _0260_;
	wire _0261_;
	wire _0262_;
	wire _0263_;
	wire _0264_;
	wire _0265_;
	wire _0266_;
	wire _0267_;
	wire _0268_;
	wire _0269_;
	wire _0270_;
	wire _0271_;
	wire _0272_;
	wire _0273_;
	wire _0274_;
	wire _0275_;
	wire _0276_;
	wire _0277_;
	wire _0278_;
	wire _0279_;
	wire _0280_;
	wire _0281_;
	wire _0282_;
	wire _0283_;
	wire _0284_;
	wire _0285_;
	wire _0286_;
	wire _0287_;
	wire _0288_;
	wire _0289_;
	wire _0290_;
	wire _0291_;
	wire _0292_;
	wire _0293_;
	wire _0294_;
	wire _0295_;
	wire _0296_;
	wire _0297_;
	wire _0298_;
	wire _0299_;
	wire _0300_;
	wire _0301_;
	wire _0302_;
	wire _0303_;
	wire _0304_;
	wire _0305_;
	wire _0306_;
	wire _0307_;
	wire _0308_;
	wire _0309_;
	wire _0310_;
	wire _0311_;
	wire _0312_;
	wire _0313_;
	wire _0314_;
	wire _0315_;
	wire _0316_;
	wire _0317_;
	wire _0318_;
	wire _0319_;
	wire _0320_;
	wire _0321_;
	wire _0322_;
	wire _0323_;
	wire _0324_;
	wire _0325_;
	wire _0326_;
	wire _0327_;
	wire _0328_;
	wire _0329_;
	wire _0330_;
	wire _0331_;
	wire _0332_;
	wire _0333_;
	wire _0334_;
	wire _0335_;
	wire _0336_;
	wire _0337_;
	wire _0338_;
	wire _0339_;
	wire _0340_;
	wire _0341_;
	wire _0342_;
	wire _0343_;
	wire _0344_;
	wire _0345_;
	wire _0346_;
	wire _0347_;
	wire _0348_;
	wire _0349_;
	wire _0350_;
	wire _0351_;
	wire _0352_;
	wire _0353_;
	wire _0354_;
	wire _0355_;
	wire _0356_;
	wire _0357_;
	wire _0358_;
	wire _0359_;
	wire _0360_;
	wire _0361_;
	wire _0362_;
	wire _0363_;
	wire _0364_;
	wire _0365_;
	wire _0366_;
	wire _0367_;
	wire _0368_;
	wire _0369_;
	wire _0370_;
	wire _0371_;
	wire _0372_;
	wire _0373_;
	wire _0374_;
	wire _0375_;
	wire _0376_;
	wire _0377_;
	wire _0378_;
	wire _0379_;
	wire _0380_;
	wire _0381_;
	wire _0382_;
	wire _0383_;
	wire _0384_;
	wire _0385_;
	wire _0386_;
	wire _0387_;
	wire _0388_;
	wire _0389_;
	wire _0390_;
	wire _0391_;
	wire _0392_;
	wire _0393_;
	wire _0394_;
	wire _0395_;
	wire _0396_;
	wire _0397_;
	wire _0398_;
	wire _0399_;
	wire _0400_;
	wire _0401_;
	wire _0402_;
	wire _0403_;
	wire _0404_;
	wire _0405_;
	wire _0406_;
	wire _0407_;
	wire _0408_;
	wire _0409_;
	wire _0410_;
	wire _0411_;
	wire _0412_;
	wire _0413_;
	wire _0414_;
	wire _0415_;
	wire _0416_;
	wire _0417_;
	wire _0418_;
	wire _0419_;
	wire _0420_;
	wire _0421_;
	wire _0422_;
	wire _0423_;
	wire _0424_;
	wire _0425_;
	wire _0426_;
	wire _0427_;
	wire _0428_;
	wire _0429_;
	wire _0430_;
	wire _0431_;
	wire _0432_;
	wire _0433_;
	wire _0434_;
	wire _0435_;
	wire _0436_;
	wire _0437_;
	wire _0438_;
	wire _0439_;
	wire _0440_;
	wire _0441_;
	wire _0442_;
	wire _0443_;
	wire _0444_;
	wire _0445_;
	wire _0446_;
	wire _0447_;
	wire _0448_;
	wire _0449_;
	wire _0450_;
	wire _0451_;
	wire _0452_;
	wire _0453_;
	wire _0454_;
	wire _0455_;
	wire _0456_;
	wire _0457_;
	wire _0458_;
	wire _0459_;
	wire _0460_;
	wire _0461_;
	wire _0462_;
	wire _0463_;
	wire _0464_;
	wire _0465_;
	wire _0466_;
	wire _0467_;
	wire _0468_;
	wire _0469_;
	wire _0470_;
	wire _0471_;
	wire _0472_;
	wire _0473_;
	wire _0474_;
	wire _0475_;
	wire _0476_;
	wire _0477_;
	wire _0478_;
	wire _0479_;
	wire _0480_;
	wire _0481_;
	wire _0482_;
	wire _0483_;
	wire _0484_;
	wire _0485_;
	wire _0486_;
	wire _0487_;
	wire _0488_;
	wire _0489_;
	wire _0490_;
	wire _0491_;
	wire _0492_;
	wire _0493_;
	wire _0494_;
	wire _0495_;
	wire _0496_;
	wire _0497_;
	wire _0498_;
	wire _0499_;
	wire _0500_;
	wire _0501_;
	wire _0502_;
	wire _0503_;
	wire _0504_;
	wire _0505_;
	wire _0506_;
	wire _0507_;
	wire _0508_;
	wire _0509_;
	wire _0510_;
	wire _0511_;
	wire _0512_;
	wire _0513_;
	wire _0514_;
	wire _0515_;
	wire _0516_;
	wire _0517_;
	wire _0518_;
	wire _0519_;
	wire _0520_;
	wire _0521_;
	wire _0522_;
	wire _0523_;
	wire _0524_;
	wire _0525_;
	wire _0526_;
	wire _0527_;
	wire _0528_;
	wire _0529_;
	wire _0530_;
	wire _0531_;
	wire _0532_;
	wire _0533_;
	wire _0534_;
	wire _0535_;
	wire _0536_;
	wire _0537_;
	wire _0538_;
	wire _0539_;
	wire _0540_;
	wire _0541_;
	wire _0542_;
	wire _0543_;
	wire _0544_;
	wire _0545_;
	wire _0546_;
	wire _0547_;
	wire _0548_;
	wire _0549_;
	wire _0550_;
	wire _0551_;
	wire _0552_;
	wire _0553_;
	wire _0554_;
	wire _0555_;
	wire _0556_;
	wire _0557_;
	wire _0558_;
	wire _0559_;
	wire _0560_;
	wire _0561_;
	wire _0562_;
	wire _0563_;
	wire _0564_;
	wire _0565_;
	wire _0566_;
	wire _0567_;
	wire _0568_;
	wire _0569_;
	wire _0570_;
	wire _0571_;
	wire _0572_;
	wire _0573_;
	wire _0574_;
	wire _0575_;
	wire _0576_;
	wire _0577_;
	wire _0578_;
	wire _0579_;
	wire _0580_;
	wire _0581_;
	wire _0582_;
	wire _0583_;
	wire _0584_;
	wire _0585_;
	wire _0586_;
	wire _0587_;
	wire _0588_;
	wire _0589_;
	wire _0590_;
	wire _0591_;
	wire _0592_;
	wire _0593_;
	wire _0594_;
	wire _0595_;
	wire _0596_;
	wire _0597_;
	wire _0598_;
	wire _0599_;
	wire _0600_;
	wire _0601_;
	wire _0602_;
	wire _0603_;
	wire _0604_;
	wire _0605_;
	wire _0606_;
	wire _0607_;
	wire _0608_;
	wire _0609_;
	wire _0610_;
	wire _0611_;
	wire _0612_;
	wire _0613_;
	wire _0614_;
	wire _0615_;
	wire _0616_;
	wire _0617_;
	wire _0618_;
	wire _0619_;
	wire _0620_;
	wire _0621_;
	wire _0622_;
	wire _0623_;
	wire _0624_;
	wire _0625_;
	wire _0626_;
	wire _0627_;
	wire _0628_;
	wire _0629_;
	wire _0630_;
	wire _0631_;
	wire _0632_;
	wire _0633_;
	wire _0634_;
	wire _0635_;
	wire _0636_;
	wire _0637_;
	wire _0638_;
	wire _0639_;
	wire _0640_;
	wire _0641_;
	wire _0642_;
	wire _0643_;
	wire _0644_;
	wire _0645_;
	wire _0646_;
	wire _0647_;
	wire _0648_;
	wire _0649_;
	wire _0650_;
	wire _0651_;
	wire _0652_;
	wire _0653_;
	wire _0654_;
	wire _0655_;
	wire _0656_;
	wire _0657_;
	wire _0658_;
	wire _0659_;
	wire _0660_;
	wire _0661_;
	wire _0662_;
	wire _0663_;
	wire _0664_;
	wire _0665_;
	wire _0666_;
	wire _0667_;
	wire _0668_;
	wire _0669_;
	wire _0670_;
	wire _0671_;
	wire _0672_;
	wire _0673_;
	wire _0674_;
	wire _0675_;
	wire _0676_;
	wire _0677_;
	wire _0678_;
	wire _0679_;
	wire _0680_;
	wire _0681_;
	wire _0682_;
	wire _0683_;
	wire _0684_;
	wire _0685_;
	wire _0686_;
	wire _0687_;
	wire _0688_;
	wire _0689_;
	wire _0690_;
	wire _0691_;
	wire _0692_;
	wire _0693_;
	wire _0694_;
	wire _0695_;
	wire _0696_;
	wire _0697_;
	wire _0698_;
	wire _0699_;
	wire _0700_;
	wire _0701_;
	wire _0702_;
	wire _0703_;
	wire _0704_;
	wire _0705_;
	wire _0706_;
	wire _0707_;
	wire _0708_;
	wire _0709_;
	wire _0710_;
	wire _0711_;
	wire _0712_;
	wire _0713_;
	wire _0714_;
	wire _0715_;
	wire _0716_;
	wire _0717_;
	wire _0718_;
	wire _0719_;
	wire _0720_;
	wire _0721_;
	wire _0722_;
	wire _0723_;
	wire _0724_;
	wire _0725_;
	wire _0726_;
	wire _0727_;
	wire _0728_;
	wire _0729_;
	wire _0730_;
	wire _0731_;
	wire _0732_;
	wire _0733_;
	wire _0734_;
	wire _0735_;
	wire _0736_;
	wire _0737_;
	wire _0738_;
	wire _0739_;
	wire _0740_;
	wire _0741_;
	wire _0742_;
	wire _0743_;
	wire _0744_;
	wire _0745_;
	wire _0746_;
	wire _0747_;
	wire _0748_;
	wire _0749_;
	wire _0750_;
	wire _0751_;
	wire _0752_;
	wire _0753_;
	wire _0754_;
	wire _0755_;
	wire _0756_;
	wire _0757_;
	wire _0758_;
	wire _0759_;
	wire _0760_;
	wire _0761_;
	wire _0762_;
	wire _0763_;
	wire _0764_;
	wire _0765_;
	wire _0766_;
	wire _0767_;
	wire _0768_;
	wire _0769_;
	wire _0770_;
	wire _0771_;
	wire _0772_;
	wire _0773_;
	wire _0774_;
	wire _0775_;
	wire _0776_;
	wire _0777_;
	wire _0778_;
	wire _0779_;
	wire _0780_;
	wire _0781_;
	wire _0782_;
	wire _0783_;
	wire _0784_;
	wire _0785_;
	wire _0786_;
	wire _0787_;
	wire _0788_;
	wire _0789_;
	wire _0790_;
	wire _0791_;
	wire _0792_;
	wire _0793_;
	wire _0794_;
	wire _0795_;
	wire _0796_;
	wire _0797_;
	wire _0798_;
	wire _0799_;
	wire _0800_;
	wire _0801_;
	wire _0802_;
	wire _0803_;
	wire _0804_;
	wire _0805_;
	wire _0806_;
	wire _0807_;
	wire _0808_;
	wire _0809_;
	wire _0810_;
	wire _0811_;
	wire _0812_;
	wire _0813_;
	wire _0814_;
	wire _0815_;
	wire _0816_;
	wire _0817_;
	wire _0818_;
	wire _0819_;
	wire _0820_;
	wire _0821_;
	wire _0822_;
	wire _0823_;
	wire _0824_;
	wire _0825_;
	wire _0826_;
	wire _0827_;
	wire _0828_;
	wire _0829_;
	wire _0830_;
	wire _0831_;
	wire _0832_;
	wire _0833_;
	wire _0834_;
	wire _0835_;
	wire _0836_;
	wire _0837_;
	wire _0838_;
	wire _0839_;
	wire _0840_;
	wire _0841_;
	wire _0842_;
	wire _0843_;
	wire _0844_;
	wire _0845_;
	wire _0846_;
	wire _0847_;
	wire _0848_;
	wire _0849_;
	wire _0850_;
	wire _0851_;
	wire _0852_;
	wire _0853_;
	wire _0854_;
	wire _0855_;
	wire _0856_;
	wire _0857_;
	wire _0858_;
	wire _0859_;
	wire _0860_;
	wire _0861_;
	wire _0862_;
	wire _0863_;
	wire _0864_;
	wire _0865_;
	wire _0866_;
	wire _0867_;
	wire _0868_;
	wire _0869_;
	wire _0870_;
	wire _0871_;
	wire _0872_;
	wire _0873_;
	wire _0874_;
	wire _0875_;
	wire _0876_;
	wire _0877_;
	wire _0878_;
	wire _0879_;
	wire _0880_;
	wire _0881_;
	wire _0882_;
	wire _0883_;
	wire _0884_;
	wire _0885_;
	wire _0886_;
	wire _0887_;
	wire _0888_;
	wire _0889_;
	wire _0890_;
	wire _0891_;
	wire _0892_;
	wire _0893_;
	wire _0894_;
	wire _0895_;
	wire _0896_;
	wire _0897_;
	wire _0898_;
	wire _0899_;
	wire _0900_;
	wire _0901_;
	wire _0902_;
	wire _0903_;
	wire _0904_;
	wire _0905_;
	wire _0906_;
	wire _0907_;
	wire _0908_;
	wire _0909_;
	wire _0910_;
	wire _0911_;
	wire _0912_;
	wire _0913_;
	wire _0914_;
	wire _0915_;
	wire _0916_;
	wire _0917_;
	wire _0918_;
	wire _0919_;
	wire _0920_;
	wire _0921_;
	wire _0922_;
	wire _0923_;
	wire _0924_;
	wire _0925_;
	wire _0926_;
	wire _0927_;
	wire _0928_;
	wire _0929_;
	wire _0930_;
	wire _0931_;
	wire _0932_;
	wire _0933_;
	wire _0934_;
	wire _0935_;
	wire _0936_;
	wire _0937_;
	wire _0938_;
	wire _0939_;
	wire _0940_;
	wire _0941_;
	wire _0942_;
	wire _0943_;
	wire _0944_;
	wire _0945_;
	wire _0946_;
	wire _0947_;
	wire _0948_;
	wire _0949_;
	wire _0950_;
	wire _0951_;
	wire _0952_;
	wire _0953_;
	wire _0954_;
	wire _0955_;
	wire _0956_;
	wire _0957_;
	wire _0958_;
	wire _0959_;
	wire _0960_;
	wire _0961_;
	wire _0962_;
	wire _0963_;
	wire _0964_;
	wire _0965_;
	wire _0966_;
	wire _0967_;
	wire _0968_;
	wire _0969_;
	wire _0970_;
	wire _0971_;
	wire _0972_;
	wire _0973_;
	wire _0974_;
	wire _0975_;
	wire _0976_;
	wire _0977_;
	wire _0978_;
	wire _0979_;
	wire _0980_;
	wire _0981_;
	wire _0982_;
	wire _0983_;
	wire _0984_;
	wire _0985_;
	wire _0986_;
	wire _0987_;
	wire _0988_;
	wire _0989_;
	wire _0990_;
	wire _0991_;
	wire _0992_;
	wire _0993_;
	wire _0994_;
	wire _0995_;
	wire _0996_;
	wire _0997_;
	wire _0998_;
	wire _0999_;
	wire _1000_;
	wire _1001_;
	wire _1002_;
	wire _1003_;
	wire _1004_;
	wire _1005_;
	wire _1006_;
	wire _1007_;
	wire _1008_;
	wire _1009_;
	wire _1010_;
	wire _1011_;
	wire _1012_;
	wire _1013_;
	wire _1014_;
	wire _1015_;
	wire _1016_;
	wire _1017_;
	wire _1018_;
	wire _1019_;
	wire _1020_;
	wire _1021_;
	wire _1022_;
	wire _1023_;
	wire _1024_;
	wire _1025_;
	wire _1026_;
	wire _1027_;
	wire _1028_;
	wire _1029_;
	wire _1030_;
	wire _1031_;
	wire _1032_;
	wire _1033_;
	wire _1034_;
	wire _1035_;
	wire _1036_;
	wire _1037_;
	wire _1038_;
	wire _1039_;
	wire _1040_;
	wire _1041_;
	wire _1042_;
	wire _1043_;
	wire _1044_;
	wire _1045_;
	wire _1046_;
	wire _1047_;
	wire _1048_;
	wire _1049_;
	wire _1050_;
	wire _1051_;
	wire _1052_;
	wire _1053_;
	wire _1054_;
	wire _1055_;
	wire _1056_;
	wire _1057_;
	wire _1058_;
	wire _1059_;
	wire _1060_;
	wire _1061_;
	wire _1062_;
	wire _1063_;
	wire _1064_;
	wire _1065_;
	wire _1066_;
	wire _1067_;
	wire _1068_;
	wire _1069_;
	wire _1070_;
	wire _1071_;
	wire _1072_;
	wire _1073_;
	wire _1074_;
	wire _1075_;
	wire _1076_;
	wire _1077_;
	wire _1078_;
	wire _1079_;
	wire _1080_;
	wire _1081_;
	wire _1082_;
	wire _1083_;
	wire _1084_;
	wire _1085_;
	wire _1086_;
	wire _1087_;
	wire _1088_;
	wire _1089_;
	wire _1090_;
	wire _1091_;
	wire _1092_;
	wire _1093_;
	wire _1094_;
	wire _1095_;
	wire _1096_;
	wire _1097_;
	wire _1098_;
	wire _1099_;
	wire _1100_;
	wire _1101_;
	wire _1102_;
	wire _1103_;
	wire _1104_;
	wire _1105_;
	wire _1106_;
	wire _1107_;
	wire _1108_;
	wire _1109_;
	wire _1110_;
	wire _1111_;
	wire _1112_;
	wire _1113_;
	wire _1114_;
	wire _1115_;
	wire _1116_;
	wire _1117_;
	wire _1118_;
	wire _1119_;
	wire _1120_;
	wire _1121_;
	wire _1122_;
	wire _1123_;
	wire _1124_;
	wire _1125_;
	wire _1126_;
	wire _1127_;
	wire _1128_;
	wire _1129_;
	wire _1130_;
	wire _1131_;
	wire _1132_;
	wire _1133_;
	wire _1134_;
	wire _1135_;
	wire _1136_;
	wire _1137_;
	wire _1138_;
	wire _1139_;
	wire _1140_;
	wire _1141_;
	wire _1142_;
	wire _1143_;
	wire _1144_;
	wire _1145_;
	wire _1146_;
	wire _1147_;
	wire _1148_;
	wire _1149_;
	wire _1150_;
	wire _1151_;
	wire _1152_;
	wire _1153_;
	wire _1154_;
	wire _1155_;
	wire _1156_;
	wire _1157_;
	wire _1158_;
	wire _1159_;
	wire _1160_;
	wire _1161_;
	wire _1162_;
	wire _1163_;
	wire _1164_;
	wire _1165_;
	wire _1166_;
	wire _1167_;
	wire _1168_;
	wire _1169_;
	wire _1170_;
	wire _1171_;
	wire _1172_;
	wire _1173_;
	wire _1174_;
	wire _1175_;
	wire _1176_;
	wire _1177_;
	wire _1178_;
	wire _1179_;
	wire _1180_;
	wire _1181_;
	wire _1182_;
	wire _1183_;
	wire _1184_;
	wire _1185_;
	wire _1186_;
	wire _1187_;
	wire _1188_;
	wire _1189_;
	wire _1190_;
	wire _1191_;
	wire _1192_;
	wire _1193_;
	wire _1194_;
	wire _1195_;
	wire _1196_;
	wire _1197_;
	wire _1198_;
	wire _1199_;
	wire _1200_;
	wire _1201_;
	wire _1202_;
	wire _1203_;
	wire _1204_;
	wire _1205_;
	wire _1206_;
	wire _1207_;
	wire _1208_;
	wire _1209_;
	wire _1210_;
	wire _1211_;
	wire _1212_;
	wire _1213_;
	wire _1214_;
	wire _1215_;
	wire _1216_;
	wire _1217_;
	wire _1218_;
	wire _1219_;
	wire _1220_;
	wire _1221_;
	wire _1222_;
	wire _1223_;
	wire _1224_;
	wire _1225_;
	wire _1226_;
	wire _1227_;
	wire _1228_;
	wire _1229_;
	wire _1230_;
	wire _1231_;
	wire _1232_;
	wire _1233_;
	wire _1234_;
	wire _1235_;
	wire _1236_;
	wire _1237_;
	wire _1238_;
	wire _1239_;
	wire _1240_;
	wire _1241_;
	wire _1242_;
	wire _1243_;
	wire _1244_;
	wire _1245_;
	wire _1246_;
	wire _1247_;
	wire _1248_;
	wire _1249_;
	wire _1250_;
	wire _1251_;
	wire _1252_;
	wire _1253_;
	wire _1254_;
	wire _1255_;
	wire _1256_;
	wire _1257_;
	wire _1258_;
	wire _1259_;
	wire _1260_;
	wire _1261_;
	wire _1262_;
	wire _1263_;
	wire _1264_;
	wire _1265_;
	wire _1266_;
	wire _1267_;
	wire _1268_;
	wire _1269_;
	wire _1270_;
	wire _1271_;
	wire _1272_;
	wire _1273_;
	wire _1274_;
	wire _1275_;
	wire _1276_;
	wire _1277_;
	wire _1278_;
	wire _1279_;
	wire _1280_;
	wire _1281_;
	wire _1282_;
	wire _1283_;
	wire _1284_;
	wire _1285_;
	wire _1286_;
	wire _1287_;
	wire _1288_;
	wire _1289_;
	wire _1290_;
	wire _1291_;
	wire _1292_;
	wire _1293_;
	wire _1294_;
	wire _1295_;
	wire _1296_;
	wire _1297_;
	wire _1298_;
	wire _1299_;
	wire _1300_;
	wire _1301_;
	wire _1302_;
	wire _1303_;
	wire _1304_;
	wire _1305_;
	wire _1306_;
	wire _1307_;
	wire _1308_;
	wire _1309_;
	wire _1310_;
	wire _1311_;
	wire _1312_;
	wire _1313_;
	wire _1314_;
	wire _1315_;
	wire _1316_;
	wire _1317_;
	wire _1318_;
	wire _1319_;
	wire _1320_;
	wire _1321_;
	wire _1322_;
	wire _1323_;
	wire _1324_;
	wire _1325_;
	wire _1326_;
	wire _1327_;
	wire _1328_;
	wire _1329_;
	wire _1330_;
	wire _1331_;
	wire _1332_;
	wire _1333_;
	wire _1334_;
	wire _1335_;
	wire _1336_;
	wire _1337_;
	wire _1338_;
	wire _1339_;
	wire _1340_;
	wire _1341_;
	wire _1342_;
	wire _1343_;
	wire _1344_;
	wire _1345_;
	wire _1346_;
	wire _1347_;
	wire _1348_;
	wire _1349_;
	wire _1350_;
	wire _1351_;
	wire _1352_;
	wire _1353_;
	wire _1354_;
	wire _1355_;
	wire _1356_;
	wire _1357_;
	wire _1358_;
	wire _1359_;
	wire _1360_;
	wire _1361_;
	wire _1362_;
	wire _1363_;
	wire _1364_;
	wire _1365_;
	wire _1366_;
	wire _1367_;
	wire _1368_;
	wire _1369_;
	wire _1370_;
	wire _1371_;
	wire _1372_;
	wire _1373_;
	wire _1374_;
	wire _1375_;
	wire _1376_;
	wire _1377_;
	wire _1378_;
	wire _1379_;
	wire _1380_;
	wire _1381_;
	wire _1382_;
	wire _1383_;
	wire _1384_;
	wire _1385_;
	wire _1386_;
	wire _1387_;
	wire _1388_;
	wire _1389_;
	wire _1390_;
	wire _1391_;
	wire _1392_;
	wire _1393_;
	wire _1394_;
	wire _1395_;
	wire _1396_;
	wire _1397_;
	wire _1398_;
	wire _1399_;
	wire _1400_;
	wire _1401_;
	wire _1402_;
	wire _1403_;
	wire _1404_;
	wire _1405_;
	wire _1406_;
	wire _1407_;
	wire _1408_;
	wire _1409_;
	wire _1410_;
	wire _1411_;
	wire _1412_;
	wire _1413_;
	wire _1414_;
	wire _1415_;
	wire _1416_;
	wire _1417_;
	wire _1418_;
	wire _1419_;
	wire _1420_;
	wire _1421_;
	wire _1422_;
	wire _1423_;
	wire _1424_;
	wire _1425_;
	wire _1426_;
	wire _1427_;
	wire _1428_;
	wire _1429_;
	wire _1430_;
	wire _1431_;
	wire _1432_;
	wire _1433_;
	wire _1434_;
	wire _1435_;
	wire _1436_;
	wire _1437_;
	wire _1438_;
	wire _1439_;
	wire _1440_;
	wire _1441_;
	wire _1442_;
	wire _1443_;
	wire _1444_;
	wire _1445_;
	wire _1446_;
	wire _1447_;
	wire _1448_;
	wire _1449_;
	wire _1450_;
	wire _1451_;
	wire _1452_;
	wire _1453_;
	wire _1454_;
	wire _1455_;
	wire _1456_;
	wire _1457_;
	wire _1458_;
	wire _1459_;
	wire _1460_;
	wire _1461_;
	wire _1462_;
	wire _1463_;
	wire _1464_;
	wire _1465_;
	wire _1466_;
	wire _1467_;
	wire _1468_;
	wire _1469_;
	wire _1470_;
	wire _1471_;
	wire _1472_;
	wire _1473_;
	wire _1474_;
	wire _1475_;
	wire _1476_;
	wire _1477_;
	wire _1478_;
	wire _1479_;
	wire _1480_;
	wire _1481_;
	wire _1482_;
	wire _1483_;
	wire _1484_;
	wire _1485_;
	wire _1486_;
	wire _1487_;
	wire _1488_;
	wire _1489_;
	wire _1490_;
	wire _1491_;
	wire _1492_;
	wire _1493_;
	wire _1494_;
	wire _1495_;
	wire _1496_;
	wire _1497_;
	wire _1498_;
	wire _1499_;
	wire _1500_;
	wire _1501_;
	wire _1502_;
	wire _1503_;
	wire _1504_;
	wire _1505_;
	wire _1506_;
	wire _1507_;
	wire _1508_;
	wire _1509_;
	wire _1510_;
	wire _1511_;
	wire _1512_;
	wire _1513_;
	wire _1514_;
	wire _1515_;
	wire _1516_;
	wire _1517_;
	wire _1518_;
	wire _1519_;
	wire _1520_;
	wire _1521_;
	wire _1522_;
	wire _1523_;
	wire _1524_;
	wire _1525_;
	wire _1526_;
	wire _1527_;
	wire _1528_;
	wire _1529_;
	wire _1530_;
	wire _1531_;
	wire _1532_;
	wire _1533_;
	wire _1534_;
	wire _1535_;
	wire _1536_;
	wire _1537_;
	wire _1538_;
	wire _1539_;
	wire _1540_;
	wire _1541_;
	wire _1542_;
	wire _1543_;
	wire _1544_;
	wire _1545_;
	wire _1546_;
	wire _1547_;
	wire _1548_;
	wire _1549_;
	wire _1550_;
	wire _1551_;
	wire _1552_;
	wire _1553_;
	wire _1554_;
	wire _1555_;
	wire _1556_;
	wire _1557_;
	wire _1558_;
	wire _1559_;
	wire _1560_;
	wire _1561_;
	wire _1562_;
	wire _1563_;
	wire _1564_;
	wire _1565_;
	wire _1566_;
	wire _1567_;
	wire _1568_;
	wire _1569_;
	wire _1570_;
	wire _1571_;
	wire _1572_;
	wire _1573_;
	wire _1574_;
	wire _1575_;
	wire _1576_;
	wire _1577_;
	wire _1578_;
	wire _1579_;
	wire _1580_;
	wire _1581_;
	wire _1582_;
	wire _1583_;
	wire _1584_;
	wire _1585_;
	wire _1586_;
	wire _1587_;
	wire _1588_;
	wire _1589_;
	wire _1590_;
	wire _1591_;
	wire _1592_;
	wire _1593_;
	wire _1594_;
	wire _1595_;
	wire _1596_;
	wire _1597_;
	wire _1598_;
	wire _1599_;
	wire _1600_;
	wire _1601_;
	wire _1602_;
	wire _1603_;
	wire _1604_;
	wire _1605_;
	wire _1606_;
	wire _1607_;
	wire _1608_;
	wire _1609_;
	wire _1610_;
	wire _1611_;
	wire _1612_;
	wire _1613_;
	wire _1614_;
	wire _1615_;
	wire _1616_;
	wire _1617_;
	wire _1618_;
	wire _1619_;
	wire _1620_;
	wire _1621_;
	wire _1622_;
	wire _1623_;
	wire _1624_;
	wire _1625_;
	wire _1626_;
	wire _1627_;
	wire _1628_;
	wire _1629_;
	wire _1630_;
	wire _1631_;
	wire _1632_;
	wire _1633_;
	wire _1634_;
	wire _1635_;
	wire _1636_;
	wire _1637_;
	wire _1638_;
	wire _1639_;
	wire _1640_;
	wire _1641_;
	wire _1642_;
	wire _1643_;
	wire _1644_;
	wire _1645_;
	wire _1646_;
	wire _1647_;
	wire _1648_;
	wire _1649_;
	wire _1650_;
	wire _1651_;
	wire _1652_;
	wire _1653_;
	wire _1654_;
	wire _1655_;
	wire _1656_;
	wire _1657_;
	wire _1658_;
	wire _1659_;
	wire _1660_;
	wire _1661_;
	wire _1662_;
	wire _1663_;
	wire _1664_;
	wire _1665_;
	wire _1666_;
	wire _1667_;
	wire _1668_;
	wire _1669_;
	wire _1670_;
	wire _1671_;
	wire _1672_;
	wire _1673_;
	wire _1674_;
	wire _1675_;
	wire _1676_;
	wire _1677_;
	wire _1678_;
	wire _1679_;
	wire _1680_;
	wire _1681_;
	wire _1682_;
	wire _1683_;
	wire _1684_;
	wire _1685_;
	wire _1686_;
	wire _1687_;
	wire _1688_;
	wire _1689_;
	wire _1690_;
	wire _1691_;
	wire _1692_;
	wire _1693_;
	wire _1694_;
	wire _1695_;
	wire _1696_;
	wire _1697_;
	wire _1698_;
	wire _1699_;
	wire _1700_;
	wire _1701_;
	wire _1702_;
	wire _1703_;
	wire _1704_;
	wire _1705_;
	wire _1706_;
	wire _1707_;
	wire _1708_;
	wire _1709_;
	wire _1710_;
	wire _1711_;
	wire _1712_;
	wire _1713_;
	wire _1714_;
	wire _1715_;
	wire _1716_;
	wire _1717_;
	wire _1718_;
	wire _1719_;
	wire _1720_;
	wire _1721_;
	wire _1722_;
	wire _1723_;
	wire _1724_;
	wire _1725_;
	wire _1726_;
	wire _1727_;
	wire _1728_;
	wire _1729_;
	wire _1730_;
	wire _1731_;
	wire _1732_;
	wire _1733_;
	wire _1734_;
	wire _1735_;
	wire _1736_;
	wire _1737_;
	wire _1738_;
	wire _1739_;
	wire _1740_;
	wire _1741_;
	wire _1742_;
	wire _1743_;
	wire _1744_;
	wire _1745_;
	wire _1746_;
	wire _1747_;
	wire _1748_;
	wire _1749_;
	wire _1750_;
	wire _1751_;
	wire _1752_;
	wire _1753_;
	wire _1754_;
	wire _1755_;
	wire _1756_;
	wire _1757_;
	wire _1758_;
	wire _1759_;
	wire _1760_;
	wire _1761_;
	wire _1762_;
	wire _1763_;
	wire _1764_;
	wire _1765_;
	wire _1766_;
	wire _1767_;
	wire _1768_;
	wire _1769_;
	wire _1770_;
	wire _1771_;
	wire _1772_;
	wire _1773_;
	wire _1774_;
	wire _1775_;
	wire _1776_;
	wire _1777_;
	wire _1778_;
	wire _1779_;
	wire _1780_;
	wire _1781_;
	wire _1782_;
	wire _1783_;
	wire _1784_;
	wire _1785_;
	wire _1786_;
	wire _1787_;
	wire _1788_;
	wire _1789_;
	wire _1790_;
	wire _1791_;
	wire _1792_;
	wire _1793_;
	wire _1794_;
	wire _1795_;
	wire _1796_;
	wire _1797_;
	wire _1798_;
	wire _1799_;
	wire _1800_;
	wire _1801_;
	wire _1802_;
	wire _1803_;
	wire _1804_;
	wire _1805_;
	wire _1806_;
	wire _1807_;
	wire _1808_;
	wire _1809_;
	wire _1810_;
	wire _1811_;
	wire _1812_;
	wire _1813_;
	wire _1814_;
	wire _1815_;
	wire _1816_;
	wire _1817_;
	wire _1818_;
	wire _1819_;
	wire _1820_;
	wire _1821_;
	wire _1822_;
	wire _1823_;
	wire _1824_;
	wire _1825_;
	wire _1826_;
	wire _1827_;
	wire _1828_;
	wire _1829_;
	wire _1830_;
	wire _1831_;
	wire _1832_;
	wire _1833_;
	wire _1834_;
	wire _1835_;
	wire _1836_;
	wire _1837_;
	wire _1838_;
	wire _1839_;
	wire _1840_;
	wire _1841_;
	wire _1842_;
	wire _1843_;
	wire _1844_;
	wire _1845_;
	wire _1846_;
	wire _1847_;
	wire _1848_;
	wire _1849_;
	wire _1850_;
	wire _1851_;
	wire _1852_;
	wire _1853_;
	wire _1854_;
	wire _1855_;
	wire _1856_;
	wire _1857_;
	wire _1858_;
	wire _1859_;
	wire _1860_;
	wire _1861_;
	wire _1862_;
	wire _1863_;
	wire _1864_;
	wire _1865_;
	wire _1866_;
	wire _1867_;
	wire _1868_;
	wire _1869_;
	wire _1870_;
	wire _1871_;
	wire _1872_;
	wire _1873_;
	wire _1874_;
	wire _1875_;
	wire _1876_;
	wire _1877_;
	wire _1878_;
	wire _1879_;
	wire _1880_;
	wire _1881_;
	wire _1882_;
	wire _1883_;
	wire _1884_;
	wire _1885_;
	wire _1886_;
	wire _1887_;
	wire _1888_;
	wire _1889_;
	wire _1890_;
	wire _1891_;
	wire _1892_;
	wire _1893_;
	wire _1894_;
	wire _1895_;
	wire _1896_;
	wire _1897_;
	wire _1898_;
	wire _1899_;
	wire _1900_;
	wire _1901_;
	wire _1902_;
	wire _1903_;
	wire _1904_;
	wire _1905_;
	wire _1906_;
	wire _1907_;
	wire _1908_;
	wire _1909_;
	wire _1910_;
	wire _1911_;
	wire _1912_;
	wire _1913_;
	wire _1914_;
	wire _1915_;
	wire _1916_;
	wire _1917_;
	wire _1918_;
	wire _1919_;
	wire _1920_;
	wire _1921_;
	wire _1922_;
	wire _1923_;
	wire _1924_;
	wire _1925_;
	wire _1926_;
	wire _1927_;
	wire _1928_;
	wire _1929_;
	wire _1930_;
	wire _1931_;
	wire _1932_;
	wire _1933_;
	wire _1934_;
	wire _1935_;
	wire _1936_;
	wire _1937_;
	wire _1938_;
	wire _1939_;
	wire _1940_;
	wire _1941_;
	wire _1942_;
	wire _1943_;
	wire _1944_;
	wire _1945_;
	wire _1946_;
	wire _1947_;
	wire _1948_;
	wire _1949_;
	wire _1950_;
	wire _1951_;
	wire _1952_;
	wire _1953_;
	wire _1954_;
	wire _1955_;
	wire _1956_;
	wire _1957_;
	wire _1958_;
	wire _1959_;
	wire _1960_;
	wire _1961_;
	wire _1962_;
	wire _1963_;
	wire _1964_;
	wire _1965_;
	wire _1966_;
	wire _1967_;
	wire _1968_;
	wire _1969_;
	wire _1970_;
	wire _1971_;
	wire _1972_;
	wire _1973_;
	wire _1974_;
	wire _1975_;
	wire _1976_;
	wire _1977_;
	wire _1978_;
	wire _1979_;
	wire _1980_;
	wire _1981_;
	wire _1982_;
	wire _1983_;
	wire _1984_;
	wire _1985_;
	wire _1986_;
	wire _1987_;
	wire _1988_;
	wire _1989_;
	wire _1990_;
	wire _1991_;
	wire _1992_;
	wire _1993_;
	wire _1994_;
	wire _1995_;
	wire _1996_;
	wire _1997_;
	wire _1998_;
	wire _1999_;
	wire _2000_;
	wire _2001_;
	wire _2002_;
	wire _2003_;
	wire _2004_;
	wire _2005_;
	wire _2006_;
	wire _2007_;
	wire _2008_;
	wire _2009_;
	wire _2010_;
	wire _2011_;
	wire _2012_;
	wire _2013_;
	wire _2014_;
	wire _2015_;
	wire _2016_;
	wire _2017_;
	wire _2018_;
	wire _2019_;
	wire _2020_;
	wire _2021_;
	wire _2022_;
	wire _2023_;
	wire _2024_;
	wire _2025_;
	wire _2026_;
	wire _2027_;
	wire _2028_;
	wire _2029_;
	wire _2030_;
	wire _2031_;
	wire _2032_;
	wire _2033_;
	wire _2034_;
	wire _2035_;
	wire _2036_;
	wire _2037_;
	wire _2038_;
	wire _2039_;
	wire _2040_;
	wire _2041_;
	wire _2042_;
	wire _2043_;
	wire _2044_;
	wire _2045_;
	wire _2046_;
	wire _2047_;
	wire _2048_;
	wire _2049_;
	wire _2050_;
	wire _2051_;
	wire _2052_;
	wire _2053_;
	wire _2054_;
	wire _2055_;
	wire _2056_;
	wire _2057_;
	wire _2058_;
	wire _2059_;
	wire _2060_;
	wire _2061_;
	wire _2062_;
	wire _2063_;
	wire _2064_;
	wire _2065_;
	wire _2066_;
	wire _2067_;
	wire _2068_;
	wire _2069_;
	wire _2070_;
	wire _2071_;
	wire _2072_;
	wire _2073_;
	wire _2074_;
	wire _2075_;
	wire _2076_;
	wire _2077_;
	wire _2078_;
	wire _2079_;
	wire _2080_;
	wire _2081_;
	wire _2082_;
	wire _2083_;
	wire _2084_;
	wire _2085_;
	wire _2086_;
	wire _2087_;
	wire _2088_;
	wire _2089_;
	wire _2090_;
	wire _2091_;
	wire _2092_;
	wire _2093_;
	wire _2094_;
	wire _2095_;
	wire _2096_;
	wire _2097_;
	wire _2098_;
	wire _2099_;
	wire _2100_;
	wire _2101_;
	wire _2102_;
	wire _2103_;
	wire _2104_;
	wire _2105_;
	wire _2106_;
	wire _2107_;
	wire _2108_;
	wire _2109_;
	wire _2110_;
	wire _2111_;
	wire _2112_;
	wire _2113_;
	wire _2114_;
	wire _2115_;
	wire _2116_;
	wire _2117_;
	wire _2118_;
	wire _2119_;
	wire _2120_;
	wire _2121_;
	wire _2122_;
	wire _2123_;
	wire _2124_;
	wire _2125_;
	wire _2126_;
	wire _2127_;
	wire _2128_;
	wire _2129_;
	wire _2130_;
	wire _2131_;
	wire _2132_;
	wire _2133_;
	wire _2134_;
	wire _2135_;
	wire _2136_;
	wire _2137_;
	wire _2138_;
	wire _2139_;
	wire _2140_;
	wire _2141_;
	wire _2142_;
	wire _2143_;
	wire _2144_;
	wire _2145_;
	wire _2146_;
	wire _2147_;
	wire _2148_;
	wire _2149_;
	wire _2150_;
	wire _2151_;
	wire _2152_;
	wire _2153_;
	wire _2154_;
	wire _2155_;
	wire _2156_;
	wire _2157_;
	wire _2158_;
	wire _2159_;
	wire _2160_;
	wire _2161_;
	wire _2162_;
	wire _2163_;
	wire _2164_;
	wire _2165_;
	wire _2166_;
	wire _2167_;
	wire _2168_;
	wire _2169_;
	wire _2170_;
	wire _2171_;
	wire _2172_;
	wire _2173_;
	wire _2174_;
	wire _2175_;
	wire _2176_;
	wire _2177_;
	wire _2178_;
	wire _2179_;
	wire _2180_;
	wire _2181_;
	wire _2182_;
	wire _2183_;
	wire _2184_;
	wire _2185_;
	wire _2186_;
	wire _2187_;
	wire _2188_;
	wire _2189_;
	wire _2190_;
	wire _2191_;
	wire _2192_;
	wire _2193_;
	wire _2194_;
	wire _2195_;
	wire _2196_;
	wire _2197_;
	wire _2198_;
	wire _2199_;
	wire _2200_;
	wire _2201_;
	wire _2202_;
	wire _2203_;
	wire _2204_;
	wire _2205_;
	wire _2206_;
	wire _2207_;
	wire _2208_;
	wire _2209_;
	wire _2210_;
	wire _2211_;
	wire _2212_;
	wire _2213_;
	wire _2214_;
	wire _2215_;
	wire _2216_;
	wire _2217_;
	wire _2218_;
	wire _2219_;
	wire _2220_;
	wire _2221_;
	wire _2222_;
	wire _2223_;
	wire _2224_;
	wire _2225_;
	wire _2226_;
	wire _2227_;
	wire _2228_;
	wire _2229_;
	wire _2230_;
	wire _2231_;
	wire _2232_;
	wire _2233_;
	wire _2234_;
	wire _2235_;
	wire _2236_;
	wire _2237_;
	wire _2238_;
	wire _2239_;
	wire _2240_;
	wire _2241_;
	wire _2242_;
	wire _2243_;
	wire _2244_;
	wire _2245_;
	wire _2246_;
	wire _2247_;
	wire _2248_;
	wire _2249_;
	wire _2250_;
	wire _2251_;
	wire _2252_;
	wire _2253_;
	wire _2254_;
	wire _2255_;
	wire _2256_;
	wire _2257_;
	wire _2258_;
	wire _2259_;
	wire _2260_;
	wire _2261_;
	wire _2262_;
	wire _2263_;
	wire _2264_;
	wire _2265_;
	wire _2266_;
	wire _2267_;
	wire _2268_;
	wire _2269_;
	wire _2270_;
	wire _2271_;
	wire _2272_;
	wire _2273_;
	wire _2274_;
	wire _2275_;
	wire _2276_;
	wire _2277_;
	wire _2278_;
	wire _2279_;
	wire _2280_;
	wire _2281_;
	wire _2282_;
	wire _2283_;
	wire _2284_;
	wire _2285_;
	wire _2286_;
	wire _2287_;
	wire _2288_;
	wire _2289_;
	wire _2290_;
	wire _2291_;
	wire _2292_;
	wire _2293_;
	wire _2294_;
	wire _2295_;
	wire _2296_;
	wire _2297_;
	wire _2298_;
	wire _2299_;
	wire _2300_;
	wire _2301_;
	wire _2302_;
	wire _2303_;
	wire _2304_;
	wire _2305_;
	wire _2306_;
	wire _2307_;
	wire _2308_;
	wire _2309_;
	wire _2310_;
	wire _2311_;
	wire _2312_;
	wire _2313_;
	wire _2314_;
	wire _2315_;
	wire _2316_;
	wire _2317_;
	wire _2318_;
	wire _2319_;
	wire _2320_;
	wire _2321_;
	wire _2322_;
	wire _2323_;
	wire _2324_;
	wire _2325_;
	wire _2326_;
	wire _2327_;
	wire _2328_;
	wire _2329_;
	wire _2330_;
	wire _2331_;
	wire _2332_;
	wire _2333_;
	wire _2334_;
	wire _2335_;
	wire _2336_;
	wire _2337_;
	wire _2338_;
	wire _2339_;
	wire _2340_;
	wire _2341_;
	wire _2342_;
	wire _2343_;
	wire _2344_;
	wire _2345_;
	wire _2346_;
	wire _2347_;
	wire _2348_;
	wire _2349_;
	wire _2350_;
	wire _2351_;
	wire _2352_;
	wire _2353_;
	wire _2354_;
	wire _2355_;
	wire _2356_;
	wire _2357_;
	wire _2358_;
	wire _2359_;
	wire _2360_;
	wire _2361_;
	wire _2362_;
	wire _2363_;
	wire _2364_;
	wire _2365_;
	wire _2366_;
	wire _2367_;
	wire _2368_;
	wire _2369_;
	wire _2370_;
	wire _2371_;
	wire _2372_;
	wire _2373_;
	wire _2374_;
	wire _2375_;
	wire _2376_;
	wire _2377_;
	wire _2378_;
	wire _2379_;
	wire _2380_;
	wire _2381_;
	wire _2382_;
	wire _2383_;
	wire _2384_;
	wire _2385_;
	wire _2386_;
	wire _2387_;
	wire _2388_;
	wire _2389_;
	wire _2390_;
	wire _2391_;
	wire _2392_;
	wire _2393_;
	wire _2394_;
	wire _2395_;
	wire _2396_;
	wire _2397_;
	wire _2398_;
	wire _2399_;
	wire _2400_;
	wire _2401_;
	wire _2402_;
	wire _2403_;
	wire _2404_;
	wire _2405_;
	wire _2406_;
	wire _2407_;
	wire _2408_;
	wire _2409_;
	wire _2410_;
	wire _2411_;
	wire _2412_;
	wire _2413_;
	wire _2414_;
	wire _2415_;
	wire _2416_;
	wire _2417_;
	wire _2418_;
	wire _2419_;
	wire _2420_;
	wire _2421_;
	wire _2422_;
	wire _2423_;
	wire _2424_;
	wire _2425_;
	wire _2426_;
	wire _2427_;
	wire _2428_;
	wire _2429_;
	wire _2430_;
	wire _2431_;
	wire _2432_;
	wire _2433_;
	wire _2434_;
	wire _2435_;
	wire _2436_;
	wire _2437_;
	wire _2438_;
	wire _2439_;
	wire _2440_;
	wire _2441_;
	wire _2442_;
	wire _2443_;
	wire _2444_;
	wire _2445_;
	wire _2446_;
	wire _2447_;
	wire _2448_;
	wire _2449_;
	wire _2450_;
	wire _2451_;
	wire _2452_;
	wire _2453_;
	wire _2454_;
	wire _2455_;
	wire _2456_;
	wire _2457_;
	wire _2458_;
	wire _2459_;
	wire _2460_;
	wire _2461_;
	wire _2462_;
	wire _2463_;
	wire _2464_;
	wire _2465_;
	wire _2466_;
	wire _2467_;
	wire _2468_;
	wire _2469_;
	wire _2470_;
	wire _2471_;
	wire _2472_;
	wire _2473_;
	wire _2474_;
	wire _2475_;
	wire _2476_;
	wire _2477_;
	wire _2478_;
	wire _2479_;
	wire _2480_;
	wire _2481_;
	wire _2482_;
	wire _2483_;
	wire _2484_;
	wire _2485_;
	wire _2486_;
	wire _2487_;
	wire _2488_;
	wire _2489_;
	wire _2490_;
	wire _2491_;
	wire _2492_;
	wire _2493_;
	wire _2494_;
	wire _2495_;
	wire _2496_;
	wire _2497_;
	wire _2498_;
	wire _2499_;
	wire _2500_;
	wire _2501_;
	wire _2502_;
	wire _2503_;
	wire _2504_;
	wire _2505_;
	wire _2506_;
	wire _2507_;
	wire _2508_;
	wire _2509_;
	wire _2510_;
	wire _2511_;
	wire _2512_;
	wire _2513_;
	wire _2514_;
	wire _2515_;
	wire _2516_;
	wire _2517_;
	wire _2518_;
	wire _2519_;
	wire _2520_;
	wire _2521_;
	wire _2522_;
	wire _2523_;
	wire _2524_;
	wire _2525_;
	wire _2526_;
	wire _2527_;
	wire _2528_;
	wire _2529_;
	wire _2530_;
	wire _2531_;
	wire _2532_;
	wire _2533_;
	wire _2534_;
	wire _2535_;
	wire _2536_;
	wire _2537_;
	wire _2538_;
	wire _2539_;
	wire _2540_;
	wire _2541_;
	wire _2542_;
	wire _2543_;
	wire _2544_;
	wire _2545_;
	wire _2546_;
	wire _2547_;
	wire _2548_;
	wire _2549_;
	wire _2550_;
	wire _2551_;
	wire _2552_;
	wire _2553_;
	wire _2554_;
	wire _2555_;
	wire _2556_;
	wire _2557_;
	wire _2558_;
	wire _2559_;
	wire _2560_;
	wire _2561_;
	wire _2562_;
	wire _2563_;
	wire _2564_;
	wire _2565_;
	wire _2566_;
	wire _2567_;
	wire _2568_;
	wire _2569_;
	wire _2570_;
	wire _2571_;
	wire _2572_;
	wire _2573_;
	wire _2574_;
	wire _2575_;
	wire _2576_;
	wire _2577_;
	wire _2578_;
	wire _2579_;
	wire _2580_;
	wire _2581_;
	wire _2582_;
	wire _2583_;
	wire _2584_;
	wire _2585_;
	wire _2586_;
	wire _2587_;
	wire _2588_;
	wire _2589_;
	wire _2590_;
	wire _2591_;
	wire _2592_;
	wire _2593_;
	wire _2594_;
	wire _2595_;
	wire _2596_;
	wire _2597_;
	wire _2598_;
	wire _2599_;
	wire _2600_;
	wire _2601_;
	wire _2602_;
	wire _2603_;
	wire _2604_;
	wire _2605_;
	wire _2606_;
	wire _2607_;
	wire _2608_;
	wire _2609_;
	wire _2610_;
	wire _2611_;
	wire _2612_;
	wire _2613_;
	wire _2614_;
	wire _2615_;
	wire _2616_;
	wire _2617_;
	wire _2618_;
	wire _2619_;
	wire _2620_;
	wire _2621_;
	wire _2622_;
	wire _2623_;
	wire _2624_;
	wire _2625_;
	wire _2626_;
	wire _2627_;
	wire _2628_;
	wire _2629_;
	wire _2630_;
	wire _2631_;
	wire _2632_;
	wire _2633_;
	wire _2634_;
	wire _2635_;
	wire _2636_;
	wire _2637_;
	wire _2638_;
	wire _2639_;
	wire _2640_;
	wire _2641_;
	wire _2642_;
	wire _2643_;
	wire _2644_;
	wire _2645_;
	wire _2646_;
	wire _2647_;
	wire _2648_;
	wire _2649_;
	wire _2650_;
	wire _2651_;
	wire _2652_;
	wire _2653_;
	wire _2654_;
	wire _2655_;
	wire _2656_;
	wire _2657_;
	wire _2658_;
	wire _2659_;
	wire _2660_;
	wire _2661_;
	wire _2662_;
	wire _2663_;
	wire _2664_;
	wire _2665_;
	wire _2666_;
	wire _2667_;
	wire _2668_;
	wire _2669_;
	wire _2670_;
	wire _2671_;
	wire _2672_;
	wire _2673_;
	wire _2674_;
	wire _2675_;
	wire _2676_;
	wire _2677_;
	wire _2678_;
	wire _2679_;
	wire _2680_;
	wire _2681_;
	wire _2682_;
	wire _2683_;
	wire _2684_;
	wire _2685_;
	wire _2686_;
	wire _2687_;
	wire _2688_;
	wire _2689_;
	wire _2690_;
	wire _2691_;
	wire _2692_;
	wire _2693_;
	wire _2694_;
	wire _2695_;
	wire _2696_;
	wire _2697_;
	wire _2698_;
	wire _2699_;
	wire _2700_;
	wire _2701_;
	wire _2702_;
	wire _2703_;
	wire _2704_;
	wire _2705_;
	wire _2706_;
	wire _2707_;
	wire _2708_;
	wire _2709_;
	wire _2710_;
	wire _2711_;
	wire _2712_;
	wire _2713_;
	wire _2714_;
	wire _2715_;
	wire _2716_;
	wire _2717_;
	wire _2718_;
	wire _2719_;
	wire _2720_;
	wire _2721_;
	wire _2722_;
	wire _2723_;
	wire _2724_;
	wire _2725_;
	wire _2726_;
	wire _2727_;
	wire _2728_;
	wire _2729_;
	wire _2730_;
	wire _2731_;
	wire _2732_;
	wire _2733_;
	wire _2734_;
	wire _2735_;
	wire _2736_;
	wire _2737_;
	wire _2738_;
	wire _2739_;
	wire _2740_;
	wire _2741_;
	wire _2742_;
	wire _2743_;
	wire _2744_;
	wire _2745_;
	wire _2746_;
	wire _2747_;
	wire _2748_;
	wire _2749_;
	wire _2750_;
	wire _2751_;
	wire _2752_;
	wire _2753_;
	wire _2754_;
	wire _2755_;
	wire _2756_;
	wire _2757_;
	wire _2758_;
	wire _2759_;
	wire _2760_;
	wire _2761_;
	wire _2762_;
	wire _2763_;
	wire _2764_;
	wire _2765_;
	wire _2766_;
	wire _2767_;
	wire _2768_;
	wire _2769_;
	wire _2770_;
	wire _2771_;
	wire _2772_;
	wire _2773_;
	wire _2774_;
	wire _2775_;
	wire _2776_;
	wire _2777_;
	wire _2778_;
	wire _2779_;
	wire _2780_;
	wire _2781_;
	wire _2782_;
	wire _2783_;
	wire _2784_;
	wire _2785_;
	wire _2786_;
	wire _2787_;
	wire _2788_;
	wire _2789_;
	wire _2790_;
	wire _2791_;
	wire _2792_;
	wire _2793_;
	wire _2794_;
	wire _2795_;
	wire _2796_;
	wire _2797_;
	wire _2798_;
	wire _2799_;
	wire _2800_;
	wire _2801_;
	wire _2802_;
	wire _2803_;
	wire _2804_;
	wire _2805_;
	wire _2806_;
	wire _2807_;
	wire _2808_;
	wire _2809_;
	wire _2810_;
	wire _2811_;
	wire _2812_;
	wire _2813_;
	wire _2814_;
	wire _2815_;
	wire _2816_;
	wire _2817_;
	wire _2818_;
	wire _2819_;
	wire _2820_;
	wire _2821_;
	wire _2822_;
	wire _2823_;
	wire _2824_;
	wire _2825_;
	wire _2826_;
	wire _2827_;
	wire _2828_;
	wire _2829_;
	wire _2830_;
	wire _2831_;
	wire _2832_;
	wire _2833_;
	wire _2834_;
	wire _2835_;
	wire _2836_;
	wire _2837_;
	wire _2838_;
	wire _2839_;
	wire _2840_;
	wire _2841_;
	wire _2842_;
	wire _2843_;
	wire _2844_;
	wire _2845_;
	wire _2846_;
	wire _2847_;
	wire _2848_;
	wire _2849_;
	wire _2850_;
	wire _2851_;
	wire _2852_;
	wire _2853_;
	wire _2854_;
	wire _2855_;
	wire _2856_;
	wire _2857_;
	wire _2858_;
	wire _2859_;
	wire _2860_;
	wire _2861_;
	wire _2862_;
	wire _2863_;
	wire _2864_;
	wire _2865_;
	wire _2866_;
	wire _2867_;
	wire _2868_;
	wire _2869_;
	wire _2870_;
	wire _2871_;
	wire _2872_;
	wire _2873_;
	wire _2874_;
	wire _2875_;
	wire _2876_;
	wire _2877_;
	wire _2878_;
	wire _2879_;
	wire _2880_;
	wire _2881_;
	wire _2882_;
	wire _2883_;
	wire _2884_;
	wire _2885_;
	wire _2886_;
	wire _2887_;
	wire _2888_;
	wire _2889_;
	wire _2890_;
	wire _2891_;
	wire _2892_;
	wire _2893_;
	wire _2894_;
	wire _2895_;
	wire _2896_;
	wire _2897_;
	wire _2898_;
	wire _2899_;
	wire _2900_;
	wire _2901_;
	wire _2902_;
	wire _2903_;
	wire _2904_;
	wire _2905_;
	wire _2906_;
	wire _2907_;
	wire _2908_;
	wire _2909_;
	wire _2910_;
	wire _2911_;
	wire _2912_;
	wire _2913_;
	wire _2914_;
	wire _2915_;
	wire _2916_;
	wire _2917_;
	wire _2918_;
	wire _2919_;
	wire _2920_;
	wire _2921_;
	wire _2922_;
	wire _2923_;
	wire _2924_;
	wire _2925_;
	wire _2926_;
	wire _2927_;
	wire _2928_;
	wire _2929_;
	wire _2930_;
	wire _2931_;
	wire _2932_;
	wire _2933_;
	wire _2934_;
	wire _2935_;
	wire _2936_;
	wire _2937_;
	wire _2938_;
	wire _2939_;
	wire _2940_;
	wire _2941_;
	wire _2942_;
	wire _2943_;
	wire _2944_;
	wire _2945_;
	wire _2946_;
	wire _2947_;
	wire _2948_;
	wire _2949_;
	wire _2950_;
	wire _2951_;
	wire _2952_;
	wire _2953_;
	wire _2954_;
	wire _2955_;
	wire _2956_;
	wire _2957_;
	wire _2958_;
	wire _2959_;
	wire _2960_;
	wire _2961_;
	wire _2962_;
	wire _2963_;
	wire _2964_;
	wire _2965_;
	wire _2966_;
	wire _2967_;
	wire _2968_;
	wire _2969_;
	wire _2970_;
	wire _2971_;
	wire _2972_;
	wire _2973_;
	wire _2974_;
	wire _2975_;
	wire _2976_;
	wire _2977_;
	wire _2978_;
	wire _2979_;
	wire _2980_;
	wire _2981_;
	wire _2982_;
	wire _2983_;
	wire _2984_;
	wire _2985_;
	wire _2986_;
	wire _2987_;
	wire _2988_;
	wire _2989_;
	wire _2990_;
	wire _2991_;
	wire _2992_;
	wire _2993_;
	wire _2994_;
	wire _2995_;
	wire _2996_;
	wire _2997_;
	wire _2998_;
	wire _2999_;
	wire _3000_;
	wire _3001_;
	wire _3002_;
	wire _3003_;
	wire _3004_;
	wire _3005_;
	wire _3006_;
	wire _3007_;
	wire _3008_;
	wire _3009_;
	wire _3010_;
	wire _3011_;
	wire _3012_;
	wire _3013_;
	wire _3014_;
	wire _3015_;
	wire _3016_;
	wire _3017_;
	wire _3018_;
	wire _3019_;
	wire _3020_;
	wire _3021_;
	wire _3022_;
	wire _3023_;
	wire _3024_;
	wire _3025_;
	wire _3026_;
	wire _3027_;
	wire _3028_;
	wire _3029_;
	wire _3030_;
	wire _3031_;
	wire _3032_;
	wire _3033_;
	wire _3034_;
	wire _3035_;
	wire _3036_;
	wire _3037_;
	wire _3038_;
	wire _3039_;
	wire _3040_;
	wire _3041_;
	wire _3042_;
	wire _3043_;
	wire _3044_;
	wire _3045_;
	wire _3046_;
	wire _3047_;
	wire _3048_;
	wire _3049_;
	wire _3050_;
	wire _3051_;
	wire _3052_;
	wire _3053_;
	wire _3054_;
	wire _3055_;
	wire _3056_;
	wire _3057_;
	wire _3058_;
	wire _3059_;
	wire _3060_;
	wire _3061_;
	wire _3062_;
	wire _3063_;
	wire _3064_;
	wire _3065_;
	wire _3066_;
	wire _3067_;
	wire _3068_;
	wire _3069_;
	wire _3070_;
	wire _3071_;
	wire _3072_;
	wire _3073_;
	wire _3074_;
	wire _3075_;
	wire _3076_;
	wire _3077_;
	wire _3078_;
	wire _3079_;
	wire _3080_;
	wire _3081_;
	wire _3082_;
	wire _3083_;
	wire _3084_;
	wire _3085_;
	wire _3086_;
	wire _3087_;
	wire _3088_;
	wire _3089_;
	wire _3090_;
	wire _3091_;
	wire _3092_;
	wire _3093_;
	wire _3094_;
	wire _3095_;
	wire _3096_;
	wire _3097_;
	wire _3098_;
	wire _3099_;
	wire _3100_;
	wire _3101_;
	wire _3102_;
	wire _3103_;
	wire _3104_;
	wire _3105_;
	wire _3106_;
	wire _3107_;
	wire _3108_;
	wire _3109_;
	wire _3110_;
	wire _3111_;
	wire _3112_;
	wire _3113_;
	wire _3114_;
	wire _3115_;
	wire _3116_;
	wire _3117_;
	wire _3118_;
	wire _3119_;
	wire _3120_;
	wire _3121_;
	wire _3122_;
	wire _3123_;
	wire _3124_;
	wire _3125_;
	wire _3126_;
	wire _3127_;
	wire _3128_;
	wire _3129_;
	wire _3130_;
	wire _3131_;
	wire _3132_;
	wire _3133_;
	wire _3134_;
	wire _3135_;
	wire _3136_;
	wire _3137_;
	wire _3138_;
	wire _3139_;
	wire _3140_;
	wire _3141_;
	wire _3142_;
	wire _3143_;
	wire _3144_;
	wire _3145_;
	wire _3146_;
	wire _3147_;
	wire _3148_;
	wire _3149_;
	wire _3150_;
	wire _3151_;
	wire _3152_;
	wire _3153_;
	wire _3154_;
	wire _3155_;
	wire _3156_;
	wire _3157_;
	wire _3158_;
	wire _3159_;
	wire _3160_;
	wire _3161_;
	wire _3162_;
	wire _3163_;
	wire _3164_;
	wire _3165_;
	wire _3166_;
	wire _3167_;
	wire _3168_;
	wire _3169_;
	wire _3170_;
	wire _3171_;
	wire _3172_;
	wire _3173_;
	wire _3174_;
	wire _3175_;
	wire _3176_;
	wire _3177_;
	wire _3178_;
	wire _3179_;
	wire _3180_;
	wire _3181_;
	wire _3182_;
	wire _3183_;
	wire _3184_;
	wire _3185_;
	wire _3186_;
	wire _3187_;
	wire _3188_;
	wire _3189_;
	wire _3190_;
	wire _3191_;
	wire _3192_;
	wire _3193_;
	wire _3194_;
	wire _3195_;
	wire _3196_;
	wire _3197_;
	wire _3198_;
	wire _3199_;
	wire _3200_;
	wire _3201_;
	wire _3202_;
	wire _3203_;
	wire _3204_;
	wire _3205_;
	wire _3206_;
	wire _3207_;
	wire _3208_;
	wire _3209_;
	wire _3210_;
	wire _3211_;
	wire _3212_;
	wire _3213_;
	wire _3214_;
	wire _3215_;
	wire _3216_;
	wire _3217_;
	wire _3218_;
	wire _3219_;
	wire _3220_;
	wire _3221_;
	wire _3222_;
	wire _3223_;
	wire _3224_;
	wire _3225_;
	wire _3226_;
	wire _3227_;
	wire _3228_;
	wire _3229_;
	wire _3230_;
	wire _3231_;
	wire _3232_;
	wire _3233_;
	wire _3234_;
	wire _3235_;
	wire _3236_;
	wire _3237_;
	wire _3238_;
	wire _3239_;
	wire _3240_;
	wire _3241_;
	wire _3242_;
	wire _3243_;
	wire _3244_;
	wire _3245_;
	wire _3246_;
	wire _3247_;
	wire _3248_;
	wire _3249_;
	wire _3250_;
	wire _3251_;
	wire _3252_;
	wire _3253_;
	wire _3254_;
	wire _3255_;
	wire _3256_;
	wire _3257_;
	wire _3258_;
	wire _3259_;
	wire _3260_;
	wire _3261_;
	wire _3262_;
	wire _3263_;
	wire _3264_;
	wire _3265_;
	wire _3266_;
	wire _3267_;
	wire _3268_;
	wire _3269_;
	wire _3270_;
	wire _3271_;
	wire _3272_;
	wire _3273_;
	wire _3274_;
	wire _3275_;
	wire _3276_;
	wire _3277_;
	wire _3278_;
	wire _3279_;
	wire _3280_;
	wire _3281_;
	wire _3282_;
	wire _3283_;
	wire _3284_;
	wire _3285_;
	wire _3286_;
	wire _3287_;
	wire _3288_;
	wire _3289_;
	wire _3290_;
	wire _3291_;
	wire _3292_;
	wire _3293_;
	wire _3294_;
	wire _3295_;
	wire _3296_;
	wire _3297_;
	wire _3298_;
	wire _3299_;
	wire _3300_;
	wire _3301_;
	wire _3302_;
	wire _3303_;
	wire _3304_;
	wire _3305_;
	wire _3306_;
	wire _3307_;
	wire _3308_;
	wire _3309_;
	wire _3310_;
	wire _3311_;
	wire _3312_;
	wire _3313_;
	wire _3314_;
	wire _3315_;
	wire _3316_;
	wire _3317_;
	wire _3318_;
	wire _3319_;
	wire _3320_;
	wire _3321_;
	wire _3322_;
	wire _3323_;
	wire _3324_;
	wire _3325_;
	wire _3326_;
	wire _3327_;
	wire _3328_;
	wire _3329_;
	wire _3330_;
	wire _3331_;
	wire _3332_;
	wire _3333_;
	wire _3334_;
	wire _3335_;
	wire _3336_;
	wire _3337_;
	wire _3338_;
	wire _3339_;
	wire _3340_;
	wire _3341_;
	wire _3342_;
	wire _3343_;
	wire _3344_;
	wire _3345_;
	wire _3346_;
	wire _3347_;
	wire _3348_;
	wire _3349_;
	wire _3350_;
	wire _3351_;
	wire _3352_;
	wire _3353_;
	wire _3354_;
	wire _3355_;
	wire _3356_;
	wire _3357_;
	wire _3358_;
	wire _3359_;
	wire _3360_;
	wire _3361_;
	wire _3362_;
	wire _3363_;
	wire _3364_;
	wire _3365_;
	wire _3366_;
	wire _3367_;
	wire _3368_;
	wire _3369_;
	wire _3370_;
	wire _3371_;
	wire _3372_;
	wire _3373_;
	wire _3374_;
	wire _3375_;
	wire _3376_;
	wire _3377_;
	wire _3378_;
	wire _3379_;
	wire _3380_;
	wire _3381_;
	wire _3382_;
	wire _3383_;
	wire _3384_;
	wire _3385_;
	wire _3386_;
	wire _3387_;
	wire _3388_;
	wire _3389_;
	wire _3390_;
	wire _3391_;
	wire _3392_;
	wire _3393_;
	wire _3394_;
	wire _3395_;
	wire _3396_;
	wire _3397_;
	wire _3398_;
	wire _3399_;
	wire _3400_;
	wire _3401_;
	wire _3402_;
	wire _3403_;
	wire _3404_;
	wire _3405_;
	wire _3406_;
	wire _3407_;
	wire _3408_;
	wire _3409_;
	wire _3410_;
	wire _3411_;
	wire _3412_;
	wire _3413_;
	wire _3414_;
	wire _3415_;
	wire _3416_;
	wire _3417_;
	wire _3418_;
	wire _3419_;
	wire _3420_;
	wire _3421_;
	wire _3422_;
	wire _3423_;
	wire _3424_;
	wire _3425_;
	wire _3426_;
	wire _3427_;
	wire _3428_;
	wire _3429_;
	wire _3430_;
	wire _3431_;
	wire _3432_;
	wire _3433_;
	wire _3434_;
	wire _3435_;
	wire _3436_;
	wire _3437_;
	wire _3438_;
	wire _3439_;
	wire _3440_;
	wire _3441_;
	wire _3442_;
	wire _3443_;
	wire _3444_;
	wire _3445_;
	wire _3446_;
	wire _3447_;
	wire _3448_;
	wire _3449_;
	wire _3450_;
	wire _3451_;
	wire _3452_;
	wire _3453_;
	wire _3454_;
	wire _3455_;
	wire _3456_;
	wire _3457_;
	wire _3458_;
	wire _3459_;
	wire _3460_;
	wire _3461_;
	wire _3462_;
	wire _3463_;
	wire _3464_;
	wire _3465_;
	wire _3466_;
	wire _3467_;
	wire _3468_;
	wire _3469_;
	wire _3470_;
	wire _3471_;
	wire _3472_;
	wire _3473_;
	wire _3474_;
	wire _3475_;
	wire _3476_;
	wire _3477_;
	wire _3478_;
	wire _3479_;
	wire _3480_;
	wire _3481_;
	wire _3482_;
	wire _3483_;
	wire _3484_;
	wire _3485_;
	wire _3486_;
	wire _3487_;
	wire _3488_;
	wire _3489_;
	wire _3490_;
	wire _3491_;
	wire _3492_;
	wire _3493_;
	wire _3494_;
	wire _3495_;
	wire _3496_;
	wire _3497_;
	wire _3498_;
	wire _3499_;
	wire _3500_;
	wire _3501_;
	wire _3502_;
	wire _3503_;
	wire _3504_;
	wire _3505_;
	wire _3506_;
	wire _3507_;
	wire _3508_;
	wire _3509_;
	wire _3510_;
	wire _3511_;
	wire _3512_;
	wire _3513_;
	wire _3514_;
	wire _3515_;
	wire _3516_;
	wire _3517_;
	wire _3518_;
	wire _3519_;
	wire _3520_;
	wire _3521_;
	wire _3522_;
	wire _3523_;
	wire _3524_;
	wire _3525_;
	wire _3526_;
	wire _3527_;
	wire _3528_;
	wire _3529_;
	wire _3530_;
	wire _3531_;
	wire _3532_;
	wire _3533_;
	wire _3534_;
	wire _3535_;
	wire _3536_;
	wire _3537_;
	wire _3538_;
	wire _3539_;
	wire _3540_;
	wire _3541_;
	wire _3542_;
	wire _3543_;
	wire _3544_;
	wire _3545_;
	wire _3546_;
	wire _3547_;
	wire _3548_;
	wire _3549_;
	wire _3550_;
	wire _3551_;
	wire _3552_;
	wire _3553_;
	wire _3554_;
	wire _3555_;
	wire _3556_;
	wire _3557_;
	wire _3558_;
	wire _3559_;
	wire _3560_;
	wire _3561_;
	wire _3562_;
	wire _3563_;
	wire _3564_;
	wire _3565_;
	wire _3566_;
	wire _3567_;
	wire _3568_;
	wire _3569_;
	wire _3570_;
	wire _3571_;
	wire _3572_;
	wire _3573_;
	wire _3574_;
	wire _3575_;
	wire _3576_;
	wire _3577_;
	wire _3578_;
	wire _3579_;
	wire _3580_;
	wire _3581_;
	wire _3582_;
	wire _3583_;
	wire _3584_;
	wire _3585_;
	wire _3586_;
	wire _3587_;
	wire _3588_;
	wire _3589_;
	wire _3590_;
	wire _3591_;
	wire _3592_;
	wire _3593_;
	wire _3594_;
	wire _3595_;
	wire _3596_;
	wire _3597_;
	wire _3598_;
	wire _3599_;
	wire _3600_;
	wire _3601_;
	wire _3602_;
	wire _3603_;
	wire _3604_;
	wire _3605_;
	wire _3606_;
	wire _3607_;
	wire _3608_;
	wire _3609_;
	wire _3610_;
	wire _3611_;
	wire _3612_;
	wire _3613_;
	wire _3614_;
	wire _3615_;
	wire _3616_;
	wire _3617_;
	wire _3618_;
	wire _3619_;
	wire _3620_;
	wire _3621_;
	wire _3622_;
	wire _3623_;
	wire _3624_;
	wire _3625_;
	wire _3626_;
	wire _3627_;
	wire _3628_;
	wire _3629_;
	wire _3630_;
	wire _3631_;
	wire _3632_;
	wire _3633_;
	wire _3634_;
	wire _3635_;
	wire _3636_;
	wire _3637_;
	wire _3638_;
	wire _3639_;
	wire _3640_;
	wire _3641_;
	wire _3642_;
	wire _3643_;
	wire _3644_;
	wire _3645_;
	wire _3646_;
	wire _3647_;
	wire _3648_;
	wire _3649_;
	wire _3650_;
	wire _3651_;
	wire _3652_;
	wire _3653_;
	wire _3654_;
	wire _3655_;
	wire _3656_;
	wire _3657_;
	wire _3658_;
	wire _3659_;
	wire _3660_;
	wire _3661_;
	wire _3662_;
	wire _3663_;
	wire _3664_;
	wire _3665_;
	wire _3666_;
	wire _3667_;
	wire _3668_;
	wire _3669_;
	wire _3670_;
	wire _3671_;
	wire _3672_;
	wire _3673_;
	wire _3674_;
	wire _3675_;
	wire _3676_;
	wire _3677_;
	wire _3678_;
	wire _3679_;
	wire _3680_;
	wire _3681_;
	wire _3682_;
	wire _3683_;
	wire _3684_;
	wire _3685_;
	wire _3686_;
	wire _3687_;
	wire _3688_;
	wire _3689_;
	wire _3690_;
	wire _3691_;
	wire _3692_;
	wire _3693_;
	wire _3694_;
	wire _3695_;
	wire _3696_;
	wire _3697_;
	wire _3698_;
	wire _3699_;
	wire _3700_;
	wire _3701_;
	wire _3702_;
	wire _3703_;
	wire _3704_;
	wire _3705_;
	wire _3706_;
	wire _3707_;
	wire _3708_;
	wire _3709_;
	wire _3710_;
	wire _3711_;
	wire _3712_;
	wire _3713_;
	wire _3714_;
	wire _3715_;
	wire _3716_;
	wire _3717_;
	wire _3718_;
	wire _3719_;
	wire _3720_;
	wire _3721_;
	wire _3722_;
	wire _3723_;
	wire _3724_;
	wire _3725_;
	wire _3726_;
	wire _3727_;
	wire _3728_;
	wire _3729_;
	wire _3730_;
	wire _3731_;
	wire _3732_;
	wire _3733_;
	wire _3734_;
	wire _3735_;
	wire _3736_;
	wire _3737_;
	wire _3738_;
	wire _3739_;
	wire _3740_;
	wire _3741_;
	wire _3742_;
	wire _3743_;
	wire _3744_;
	wire _3745_;
	wire _3746_;
	wire _3747_;
	wire _3748_;
	wire _3749_;
	wire _3750_;
	wire _3751_;
	wire _3752_;
	wire _3753_;
	wire _3754_;
	wire _3755_;
	wire _3756_;
	wire [3:0] _3757_;
	wire [4:0] _3758_;
	input wire [13:0] io_in;
	output wire [13:0] io_out;
	wire \mchip.clock ;
	reg [3:0] \mchip.count ;
	reg [3:0] \mchip.i ;
	wire \mchip.inst_add.add_valid ;
	wire [15:0] \mchip.inst_add.input_a ;
	wire [15:0] \mchip.inst_add.input_b ;
	wire [4:0] \mchip.inst_add.temp_3 ;
	wire [4:0] \mchip.inst_mul.expo_1_temp ;
	wire [4:0] \mchip.inst_mul.expo_2_temp ;
	wire [9:0] \mchip.inst_mul.frac_1 ;
	wire [9:0] \mchip.inst_mul.frac_2 ;
	wire [15:0] \mchip.inst_mul.input_a ;
	wire [15:0] \mchip.inst_mul.input_b ;
	wire \mchip.inst_mul.mul_valid ;
	wire \mchip.inst_mul.sign_1 ;
	wire \mchip.inst_mul.sign_2 ;
	wire [20:0] \mchip.inst_mul.temp_f_1 ;
	wire [10:0] \mchip.inst_mul.temp_f_2 ;
	wire [20:0] \mchip.inst_mul.temp_value[0] ;
	wire [20:0] \mchip.inst_mul.temp_value[10] ;
	wire [20:0] \mchip.inst_mul.temp_value[1] ;
	wire [20:0] \mchip.inst_mul.temp_value[2] ;
	wire [20:0] \mchip.inst_mul.temp_value[3] ;
	wire [20:0] \mchip.inst_mul.temp_value[4] ;
	wire [20:0] \mchip.inst_mul.temp_value[5] ;
	wire [20:0] \mchip.inst_mul.temp_value[6] ;
	wire [20:0] \mchip.inst_mul.temp_value[7] ;
	wire [20:0] \mchip.inst_mul.temp_value[8] ;
	wire [20:0] \mchip.inst_mul.temp_value[9] ;
	wire [11:0] \mchip.io_in ;
	wire [11:0] \mchip.io_out ;
	wire [31:0] \mchip.j ;
	wire \mchip.reset ;
	reg [15:0] \mchip.result ;
	wire \mchip.select ;
	wire \mchip.temp_valid_add ;
	wire \mchip.temp_valid_mul ;
	reg [15:0] \mchip.tmp_input_A ;
	reg [15:0] \mchip.tmp_input_B ;
	reg \mchip.valid ;
	reg [15:0] \mchip.value_A ;
	reg [15:0] \mchip.value_B ;
	assign _3757_[0] = ~\mchip.count [0];
	assign _0931_ = \mchip.count [2] | \mchip.count [3];
	assign _0942_ = ~(\mchip.count [1] | \mchip.count [0]);
	assign _3758_[4] = _0942_ & ~_0931_;
	assign _0963_ = \mchip.count [2] & ~\mchip.count [3];
	assign _0974_ = \mchip.count [0] | ~\mchip.count [1];
	assign _0985_ = _0963_ & ~_0974_;
	assign _0996_ = io_in[13] | ~io_in[9];
	assign _0007_ = _0985_ & ~_0996_;
	assign _1017_ = ~io_in[9];
	assign _1028_ = ~(\mchip.i [1] | \mchip.i [2]);
	assign _0008_ = _1017_ & ~_1028_;
	assign _1049_ = ~(\mchip.i [3] | \mchip.i [2]);
	assign _0009_ = _1017_ & ~_1049_;
	assign _1070_ = io_in[13] | io_in[9];
	assign _1081_ = \mchip.i [1] & ~_1070_;
	assign _1092_ = \mchip.i [3] & ~_0996_;
	assign _0003_ = _1092_ | _1081_;
	assign _1113_ = ~_0985_;
	assign _0005_ = (io_in[9] ? _1113_ : \mchip.i [2]);
	assign _0006_ = \mchip.i [0] & ~io_in[9];
	assign _1144_ = \mchip.i [0] & ~_1070_;
	assign _1155_ = \mchip.i [2] & ~_0996_;
	assign _0002_ = _1155_ | _1144_;
	assign _0004_ = io_in[9] & ~_0985_;
	assign _1186_ = \mchip.i [2] & ~_1070_;
	assign _1197_ = \mchip.i [1] & ~_0996_;
	assign _0001_ = _1197_ | _1186_;
	assign _1218_ = \mchip.i [0] & ~_0996_;
	assign _1229_ = \mchip.i [3] & ~_1070_;
	assign _1240_ = _1229_ | io_in[13];
	assign _0000_ = _1240_ | _1218_;
	assign _0051_ = ~(io_in[9] & \mchip.count [0]);
	assign _1271_ = \mchip.count [1] & \mchip.count [0];
	assign _3758_[1] = _1271_ | _0942_;
	assign _0052_ = io_in[9] & ~_3758_[1];
	assign _1302_ = ~(_1271_ ^ \mchip.count [2]);
	assign _0053_ = io_in[9] & ~_1302_;
	assign _1323_ = ~(_1271_ & \mchip.count [2]);
	assign _1334_ = _1323_ ^ \mchip.count [3];
	assign _0054_ = io_in[9] & ~_1334_;
	assign _0043_ = (\mchip.i [1] ? \mchip.result [8] : \mchip.result [0]);
	assign _0044_ = (\mchip.i [1] ? \mchip.result [9] : \mchip.result [1]);
	assign _0045_ = (\mchip.i [1] ? \mchip.result [10] : \mchip.result [2]);
	assign _0046_ = (\mchip.i [1] ? \mchip.result [11] : \mchip.result [3]);
	assign _0047_ = (\mchip.i [1] ? \mchip.result [12] : \mchip.result [4]);
	assign _0048_ = (\mchip.i [1] ? \mchip.result [13] : \mchip.result [5]);
	assign _0049_ = (\mchip.i [1] ? \mchip.result [14] : \mchip.result [6]);
	assign _0050_ = (\mchip.i [1] ? \mchip.result [15] : \mchip.result [7]);
	assign _0042_ = \mchip.valid  & ~\mchip.i [3];
	assign _1455_ = ~\mchip.value_B [11];
	assign _1466_ = ~\mchip.value_B [10];
	assign _1477_ = ~\mchip.value_B [14];
	assign _1488_ = \mchip.value_B [12] | \mchip.value_B [13];
	assign _1499_ = \mchip.value_B [10] | \mchip.value_B [11];
	assign _1510_ = _1499_ | _1488_;
	assign _1521_ = _1477_ & ~_1510_;
	assign _1532_ = _1521_ & ~_1466_;
	assign _1543_ = _1532_ & ~_1455_;
	assign _1554_ = _1543_ & \mchip.value_B [12];
	assign _1565_ = _1554_ ^ \mchip.value_B [13];
	assign _1576_ = ~\mchip.value_A [11];
	assign _1587_ = ~\mchip.value_A [10];
	assign _1598_ = ~\mchip.value_A [14];
	assign _1609_ = \mchip.value_A [12] | \mchip.value_A [13];
	assign _1620_ = \mchip.value_A [10] | \mchip.value_A [11];
	assign _1631_ = _1620_ | _1609_;
	assign _1642_ = _1598_ & ~_1631_;
	assign _1653_ = _1642_ & ~_1587_;
	assign _1664_ = _1653_ & ~_1576_;
	assign _1675_ = _1664_ & \mchip.value_A [12];
	assign _1686_ = _1675_ ^ \mchip.value_A [13];
	assign _1697_ = _1686_ & _1565_;
	assign _1708_ = ~(\mchip.value_B [12] & \mchip.value_B [13]);
	assign _1719_ = _1543_ & ~_1708_;
	assign _1730_ = _1719_ ^ \mchip.value_B [14];
	assign _1741_ = ~(\mchip.value_A [12] & \mchip.value_A [13]);
	assign _1752_ = _1664_ & ~_1741_;
	assign _1763_ = _1752_ ^ \mchip.value_A [14];
	assign _1774_ = ~(_1763_ ^ _1730_);
	assign _1785_ = _1774_ & _1697_;
	assign _1796_ = _1686_ ^ _1565_;
	assign _1807_ = _1543_ ^ \mchip.value_B [12];
	assign _1818_ = _1664_ ^ \mchip.value_A [12];
	assign _1829_ = _1818_ & _1807_;
	assign _1840_ = _1829_ & _1796_;
	assign _1851_ = _1818_ ^ _1807_;
	assign _1862_ = _1532_ ^ \mchip.value_B [11];
	assign _1873_ = _1653_ ^ \mchip.value_A [11];
	assign _1884_ = _1873_ & _1862_;
	assign _1895_ = _1884_ & _1851_;
	assign _1906_ = _1829_ ^ _1796_;
	assign _1917_ = _1906_ & _1895_;
	assign _1928_ = _1917_ | _1840_;
	assign _1939_ = _1521_ ^ \mchip.value_B [10];
	assign _1950_ = _1642_ ^ \mchip.value_A [10];
	assign _1961_ = ~(_1950_ | _1939_);
	assign _1972_ = _1873_ ^ _1862_;
	assign _1983_ = _1972_ & ~_1961_;
	assign _1994_ = _1884_ ^ _1851_;
	assign _2005_ = ~(_1994_ & _1906_);
	assign _2016_ = _1983_ & ~_2005_;
	assign _2027_ = _2016_ | _1928_;
	assign _2038_ = _1774_ ^ _1697_;
	assign _2049_ = _2038_ & _2027_;
	assign _2060_ = ~(_2049_ | _1785_);
	assign _2071_ = ~(_1763_ | _1730_);
	assign _2082_ = ~_2071_;
	assign _2093_ = _2082_ ^ _2060_;
	assign _2104_ = ~(_2071_ & _2038_);
	assign _2115_ = _2027_ & ~_2104_;
	assign _2126_ = _2082_ | _1785_;
	assign _2137_ = _2126_ | _2115_;
	assign _2148_ = ~(_2137_ & _2093_);
	assign _2159_ = ~(\mchip.value_B [0] | \mchip.value_B [1]);
	assign _2170_ = \mchip.value_B [2] | \mchip.value_B [3];
	assign _2181_ = _2159_ & ~_2170_;
	assign _2192_ = \mchip.value_B [7] | \mchip.value_B [6];
	assign _2203_ = \mchip.value_B [5] | \mchip.value_B [4];
	assign _2214_ = _2203_ | _2192_;
	assign _2225_ = _2181_ & ~_2214_;
	assign _2236_ = \mchip.value_B [9] | \mchip.value_B [8];
	assign _2246_ = _2236_ | ~_2225_;
	assign _2257_ = ~(\mchip.value_B [10] & \mchip.value_B [11]);
	assign _2268_ = _2257_ | _1708_;
	assign _2279_ = _2268_ | _1477_;
	assign _2290_ = ~(_2279_ | _2246_);
	assign _2300_ = ~(\mchip.value_A [9] | \mchip.value_A [8]);
	assign _2311_ = ~(\mchip.value_A [0] | \mchip.value_A [1]);
	assign _2322_ = \mchip.value_A [2] | \mchip.value_A [3];
	assign _2333_ = _2311_ & ~_2322_;
	assign _2344_ = \mchip.value_A [7] | \mchip.value_A [6];
	assign _2355_ = \mchip.value_A [4] | \mchip.value_A [5];
	assign _2365_ = _2355_ | _2344_;
	assign _2376_ = _2333_ & ~_2365_;
	assign _2387_ = _2376_ & _2300_;
	assign _2398_ = ~(\mchip.value_A [10] & \mchip.value_A [11]);
	assign _2409_ = _2398_ | _1741_;
	assign _2419_ = _2409_ | _1598_;
	assign _2430_ = _2387_ & ~_2419_;
	assign _2441_ = _2430_ | _2290_;
	assign _2452_ = _2148_ & ~_2441_;
	assign _2463_ = \mchip.value_B [6] & ~_1642_;
	assign _2473_ = \mchip.value_A [9] & \mchip.value_B [7];
	assign _2484_ = _2473_ & _2463_;
	assign _2495_ = \mchip.value_A [8] & \mchip.value_B [8];
	assign _2506_ = _2473_ ^ _2463_;
	assign _2516_ = _2506_ & _2495_;
	assign _2527_ = ~(_2516_ | _2484_);
	assign _2538_ = \mchip.value_A [9] & \mchip.value_B [8];
	assign _2549_ = \mchip.value_B [7] & ~_1642_;
	assign _2560_ = _2549_ ^ _2538_;
	assign _2570_ = \mchip.value_A [8] & \mchip.value_B [9];
	assign _2581_ = _2570_ ^ _2560_;
	assign _2592_ = _2581_ & ~_2527_;
	assign _2603_ = \mchip.value_A [7] & ~_1521_;
	assign _2613_ = ~(_2581_ ^ _2527_);
	assign _2624_ = _2613_ & _2603_;
	assign _2635_ = ~(_2624_ | _2592_);
	assign _2646_ = _2549_ & _2538_;
	assign _2656_ = _2570_ & _2560_;
	assign _2667_ = ~(_2656_ | _2646_);
	assign _2678_ = \mchip.value_A [9] & \mchip.value_B [9];
	assign _2688_ = \mchip.value_B [8] & ~_1642_;
	assign _2699_ = _2688_ ^ _2678_;
	assign _2710_ = \mchip.value_A [8] & ~_1521_;
	assign _2721_ = _2710_ ^ _2699_;
	assign _2731_ = ~(_2721_ ^ _2667_);
	assign _2742_ = ~(_2731_ ^ _2635_);
	assign _2752_ = \mchip.value_B [5] & ~_1642_;
	assign _2763_ = \mchip.value_A [9] & \mchip.value_B [6];
	assign _2773_ = _2763_ & _2752_;
	assign _2784_ = \mchip.value_A [8] & \mchip.value_B [7];
	assign _2794_ = _2763_ ^ _2752_;
	assign _2805_ = _2794_ & _2784_;
	assign _2816_ = ~(_2805_ | _2773_);
	assign _2826_ = _2506_ ^ _2495_;
	assign _2835_ = _2816_ | ~_2826_;
	assign _2846_ = \mchip.value_A [6] & ~_1521_;
	assign _2857_ = \mchip.value_A [7] & \mchip.value_B [9];
	assign _2860_ = _2857_ ^ _2846_;
	assign _2871_ = ~(_2826_ ^ _2816_);
	assign _2882_ = _2871_ & _2860_;
	assign _2893_ = _2835_ & ~_2882_;
	assign _2904_ = _2613_ ^ _2603_;
	assign _2915_ = _2893_ | ~_2904_;
	assign _2926_ = _2857_ & _2846_;
	assign _2936_ = ~(_2904_ ^ _2893_);
	assign _2946_ = _2936_ & _2926_;
	assign _2957_ = _2915_ & ~_2946_;
	assign _2967_ = _2742_ & ~_2957_;
	assign _2977_ = _2731_ & ~_2635_;
	assign _2987_ = _2721_ & ~_2667_;
	assign _2997_ = ~_2678_;
	assign _3006_ = _2688_ & ~_2997_;
	assign _3016_ = _2710_ & _2699_;
	assign _3025_ = ~(_3016_ | _3006_);
	assign _3034_ = \mchip.value_A [9] & ~_1521_;
	assign _3043_ = \mchip.value_B [9] & ~_1642_;
	assign _3053_ = _3043_ ^ _3034_;
	assign _3063_ = ~(_3053_ ^ _3025_);
	assign _3073_ = _3063_ ^ _2987_;
	assign _3083_ = _3073_ ^ _2977_;
	assign _3094_ = _3083_ ^ _2967_;
	assign _3103_ = _2936_ ^ _2926_;
	assign _3113_ = \mchip.value_B [4] & ~_1642_;
	assign _3122_ = \mchip.value_A [9] & \mchip.value_B [5];
	assign _3131_ = _3122_ & _3113_;
	assign _3140_ = \mchip.value_A [8] & \mchip.value_B [6];
	assign _3148_ = _3122_ ^ _3113_;
	assign _3152_ = _3148_ & _3140_;
	assign _3153_ = ~(_3152_ | _3131_);
	assign _3154_ = _2794_ ^ _2784_;
	assign _3155_ = _3153_ | ~_3154_;
	assign _3156_ = \mchip.value_A [5] & ~_1521_;
	assign _3157_ = \mchip.value_A [6] & \mchip.value_B [9];
	assign _3158_ = \mchip.value_A [7] & \mchip.value_B [8];
	assign _3159_ = _3158_ ^ _3157_;
	assign _3160_ = _3159_ ^ _3156_;
	assign _3161_ = ~(_3154_ ^ _3153_);
	assign _3162_ = _3161_ & _3160_;
	assign _3163_ = _3155_ & ~_3162_;
	assign _3164_ = _2871_ ^ _2860_;
	assign _3165_ = _3163_ | ~_3164_;
	assign _3166_ = _3158_ & _3157_;
	assign _3167_ = _3159_ & _3156_;
	assign _3168_ = _3167_ | _3166_;
	assign _3169_ = ~(_3164_ ^ _3163_);
	assign _3170_ = _3169_ & _3168_;
	assign _3171_ = _3165_ & ~_3170_;
	assign _3172_ = _3103_ & ~_3171_;
	assign _3173_ = ~(_2957_ ^ _2742_);
	assign _3174_ = _3173_ & _3172_;
	assign _3175_ = _3174_ & _3094_;
	assign _3176_ = _3173_ ^ _3172_;
	assign _3177_ = _3169_ ^ _3168_;
	assign _3178_ = \mchip.value_B [3] & ~_1642_;
	assign _3179_ = \mchip.value_A [9] & \mchip.value_B [4];
	assign _3180_ = _3179_ & _3178_;
	assign _3181_ = \mchip.value_A [8] & \mchip.value_B [5];
	assign _3182_ = _3179_ ^ _3178_;
	assign _3183_ = _3182_ & _3181_;
	assign _3184_ = ~(_3183_ | _3180_);
	assign _3185_ = _3148_ ^ _3140_;
	assign _3186_ = _3184_ | ~_3185_;
	assign _3187_ = \mchip.value_B [9] & \mchip.value_A [5];
	assign _3188_ = \mchip.value_A [6] & \mchip.value_B [8];
	assign _3189_ = \mchip.value_A [7] & \mchip.value_B [7];
	assign _3190_ = _3189_ ^ _3188_;
	assign _3191_ = _3190_ ^ _3187_;
	assign _3192_ = ~(_3185_ ^ _3184_);
	assign _3193_ = _3192_ & _3191_;
	assign _3194_ = _3186_ & ~_3193_;
	assign _3195_ = _3161_ ^ _3160_;
	assign _3196_ = _3194_ | ~_3195_;
	assign _3197_ = _3189_ & _3188_;
	assign _3198_ = _3190_ & _3187_;
	assign _3199_ = _3198_ | _3197_;
	assign _3200_ = ~(_3195_ ^ _3194_);
	assign _3201_ = _3200_ & _3199_;
	assign _3202_ = _3196_ & ~_3201_;
	assign _3203_ = _3177_ & ~_3202_;
	assign _3204_ = ~(_3171_ ^ _3103_);
	assign _3205_ = _3204_ & _3203_;
	assign _3206_ = _3205_ & _3176_;
	assign _3207_ = _3174_ ^ _3094_;
	assign _3208_ = _3207_ & _3206_;
	assign _3209_ = _3208_ | _3175_;
	assign _3210_ = _3205_ ^ _3176_;
	assign _3211_ = _3210_ & _3207_;
	assign _3212_ = \mchip.value_B [2] & ~_1642_;
	assign _3213_ = \mchip.value_A [9] & \mchip.value_B [3];
	assign _3214_ = _3213_ & _3212_;
	assign _3215_ = \mchip.value_A [8] & \mchip.value_B [4];
	assign _3216_ = _3213_ ^ _3212_;
	assign _3217_ = _3216_ & _3215_;
	assign _3218_ = ~(_3217_ | _3214_);
	assign _3219_ = _3182_ ^ _3181_;
	assign _3220_ = _3219_ & ~_3218_;
	assign _3221_ = \mchip.value_B [8] & \mchip.value_A [5];
	assign _3222_ = \mchip.value_A [6] & \mchip.value_B [7];
	assign _3223_ = \mchip.value_A [7] & \mchip.value_B [6];
	assign _3224_ = _3223_ ^ _3222_;
	assign _3225_ = _3224_ ^ _3221_;
	assign _3226_ = ~(_3219_ ^ _3218_);
	assign _3227_ = _3226_ & _3225_;
	assign _3228_ = ~(_3227_ | _3220_);
	assign _3229_ = _3192_ ^ _3191_;
	assign _3230_ = _3229_ & ~_3228_;
	assign _3231_ = \mchip.value_A [3] & ~_1521_;
	assign _3232_ = \mchip.value_B [9] & \mchip.value_A [4];
	assign _3233_ = _3232_ & _3231_;
	assign _3234_ = \mchip.value_A [4] & ~_1521_;
	assign _3235_ = ~(_3223_ & _3222_);
	assign _3236_ = _3224_ & _3221_;
	assign _3237_ = _3235_ & ~_3236_;
	assign _3238_ = ~(_3237_ ^ _3234_);
	assign _3239_ = _3238_ ^ _3233_;
	assign _3240_ = ~(_3229_ ^ _3228_);
	assign _3241_ = _3240_ & _3239_;
	assign _3242_ = ~(_3241_ | _3230_);
	assign _3243_ = _3200_ ^ _3199_;
	assign _3244_ = _3243_ & ~_3242_;
	assign _3245_ = _3234_ & ~_3237_;
	assign _3246_ = _3238_ & _3233_;
	assign _3247_ = _3246_ | _3245_;
	assign _3248_ = ~(_3243_ ^ _3242_);
	assign _3249_ = _3248_ & _3247_;
	assign _3250_ = ~(_3249_ | _3244_);
	assign _3251_ = ~(_3202_ ^ _3177_);
	assign _3252_ = _3250_ | ~_3251_;
	assign _3253_ = _3204_ ^ _3203_;
	assign _3254_ = _3252_ | ~_3253_;
	assign _3255_ = ~(_3251_ ^ _3250_);
	assign _3256_ = _3248_ ^ _3247_;
	assign _3257_ = \mchip.value_B [1] & ~_1642_;
	assign _3258_ = \mchip.value_A [9] & \mchip.value_B [2];
	assign _3259_ = _3258_ & _3257_;
	assign _3260_ = \mchip.value_A [8] & \mchip.value_B [3];
	assign _3261_ = _3258_ ^ _3257_;
	assign _3262_ = _3261_ & _3260_;
	assign _3263_ = ~(_3262_ | _3259_);
	assign _3264_ = _3216_ ^ _3215_;
	assign _3265_ = _3264_ & ~_3263_;
	assign _3266_ = \mchip.value_B [7] & \mchip.value_A [5];
	assign _3267_ = \mchip.value_A [6] & \mchip.value_B [6];
	assign _3268_ = \mchip.value_A [7] & \mchip.value_B [5];
	assign _3269_ = _3268_ ^ _3267_;
	assign _3270_ = _3269_ ^ _3266_;
	assign _3271_ = ~(_3264_ ^ _3263_);
	assign _3272_ = _3271_ & _3270_;
	assign _3273_ = ~(_3272_ | _3265_);
	assign _3274_ = _3226_ ^ _3225_;
	assign _3275_ = _3273_ | ~_3274_;
	assign _3276_ = \mchip.value_B [8] & \mchip.value_A [4];
	assign _3277_ = \mchip.value_B [9] & \mchip.value_A [3];
	assign _3278_ = _3277_ & _3276_;
	assign _3279_ = \mchip.value_A [2] & ~_1521_;
	assign _3280_ = _3277_ ^ _3276_;
	assign _3281_ = _3280_ & _3279_;
	assign _3282_ = _3281_ | _3278_;
	assign _3283_ = _3232_ ^ _3231_;
	assign _3284_ = ~(_3268_ & _3267_);
	assign _3285_ = _3269_ & _3266_;
	assign _3286_ = _3284_ & ~_3285_;
	assign _3287_ = ~(_3286_ ^ _3283_);
	assign _3288_ = _3287_ ^ _3282_;
	assign _3289_ = ~(_3274_ ^ _3273_);
	assign _3290_ = _3289_ & _3288_;
	assign _3291_ = _3275_ & ~_3290_;
	assign _3292_ = _3240_ ^ _3239_;
	assign _3293_ = _3291_ | ~_3292_;
	assign _3294_ = _3283_ & ~_3286_;
	assign _3295_ = _3287_ & _3282_;
	assign _3296_ = _3295_ | _3294_;
	assign _3297_ = ~(_3292_ ^ _3291_);
	assign _3298_ = _3297_ & _3296_;
	assign _3299_ = _3293_ & ~_3298_;
	assign _3300_ = _3256_ & ~_3299_;
	assign _3301_ = _3300_ & _3255_;
	assign _3302_ = ~(_3253_ ^ _3252_);
	assign _3303_ = _3302_ & _3301_;
	assign _3304_ = _3254_ & ~_3303_;
	assign _3305_ = _3211_ & ~_3304_;
	assign _3306_ = _3305_ | _3209_;
	assign _3307_ = ~(_3300_ ^ _3255_);
	assign _3308_ = _3302_ & ~_3307_;
	assign _3309_ = _3308_ & _3211_;
	assign _3310_ = _3299_ ^ _3256_;
	assign _3311_ = _3297_ ^ _3296_;
	assign _3312_ = \mchip.value_B [0] & ~_1642_;
	assign _3313_ = \mchip.value_A [9] & \mchip.value_B [1];
	assign _3314_ = _3313_ & _3312_;
	assign _3315_ = \mchip.value_B [2] & \mchip.value_A [8];
	assign _3316_ = _3313_ ^ _3312_;
	assign _3317_ = _3316_ & _3315_;
	assign _3318_ = ~(_3317_ | _3314_);
	assign _3319_ = _3261_ ^ _3260_;
	assign _3320_ = _3319_ & ~_3318_;
	assign _3321_ = \mchip.value_B [6] & \mchip.value_A [5];
	assign _3322_ = \mchip.value_A [6] & \mchip.value_B [5];
	assign _3323_ = \mchip.value_A [7] & \mchip.value_B [4];
	assign _3324_ = _3323_ ^ _3322_;
	assign _3325_ = _3324_ ^ _3321_;
	assign _3326_ = ~(_3319_ ^ _3318_);
	assign _3327_ = _3326_ & _3325_;
	assign _3328_ = ~(_3327_ | _3320_);
	assign _3329_ = _3271_ ^ _3270_;
	assign _3330_ = _3328_ | ~_3329_;
	assign _3331_ = \mchip.value_B [7] & \mchip.value_A [4];
	assign _3332_ = \mchip.value_B [8] & \mchip.value_A [3];
	assign _3333_ = _3332_ & _3331_;
	assign _3334_ = \mchip.value_B [9] & \mchip.value_A [2];
	assign _3335_ = _3332_ ^ _3331_;
	assign _3336_ = _3335_ & _3334_;
	assign _3337_ = _3336_ | _3333_;
	assign _3338_ = _3280_ ^ _3279_;
	assign _3339_ = ~(_3323_ & _3322_);
	assign _3340_ = _3324_ & _3321_;
	assign _3341_ = _3339_ & ~_3340_;
	assign _3342_ = ~(_3341_ ^ _3338_);
	assign _3343_ = _3342_ ^ _3337_;
	assign _3344_ = ~(_3329_ ^ _3328_);
	assign _3345_ = _3344_ & _3343_;
	assign _3346_ = _3330_ & ~_3345_;
	assign _3347_ = _3289_ ^ _3288_;
	assign _3348_ = _3346_ | ~_3347_;
	assign _3349_ = _3338_ & ~_3341_;
	assign _3350_ = _3342_ & _3337_;
	assign _3351_ = _3350_ | _3349_;
	assign _3352_ = ~(_3347_ ^ _3346_);
	assign _3353_ = _3352_ & _3351_;
	assign _3354_ = _3348_ & ~_3353_;
	assign _3355_ = _3311_ & ~_3354_;
	assign _3356_ = _3310_ | ~_3355_;
	assign _3357_ = ~(_3354_ ^ _3311_);
	assign _3358_ = \mchip.value_B [0] & \mchip.value_A [9];
	assign _3359_ = \mchip.value_B [1] & \mchip.value_A [8];
	assign _3360_ = _3359_ & _3358_;
	assign _3361_ = \mchip.value_B [2] & \mchip.value_A [7];
	assign _3362_ = _3359_ ^ _3358_;
	assign _3363_ = _3362_ & _3361_;
	assign _3364_ = ~(_3363_ | _3360_);
	assign _3365_ = _3316_ ^ _3315_;
	assign _3366_ = _3365_ & ~_3364_;
	assign _3367_ = \mchip.value_B [5] & \mchip.value_A [5];
	assign _3368_ = \mchip.value_A [6] & \mchip.value_B [4];
	assign _3369_ = \mchip.value_A [7] & \mchip.value_B [3];
	assign _3370_ = _3369_ ^ _3368_;
	assign _3371_ = _3370_ ^ _3367_;
	assign _3372_ = ~(_3365_ ^ _3364_);
	assign _3373_ = _3372_ & _3371_;
	assign _3374_ = ~(_3373_ | _3366_);
	assign _3375_ = _3326_ ^ _3325_;
	assign _3376_ = _3375_ & ~_3374_;
	assign _3377_ = \mchip.value_B [6] & \mchip.value_A [4];
	assign _3378_ = \mchip.value_B [7] & \mchip.value_A [3];
	assign _3379_ = _3378_ & _3377_;
	assign _3380_ = \mchip.value_A [2] & \mchip.value_B [8];
	assign _3381_ = ~_3380_;
	assign _3382_ = _3378_ ^ _3377_;
	assign _3383_ = _3382_ & ~_3381_;
	assign _3384_ = _3383_ | _3379_;
	assign _3385_ = _3335_ ^ _3334_;
	assign _3386_ = ~(_3369_ & _3368_);
	assign _3387_ = _3370_ & _3367_;
	assign _3388_ = _3386_ & ~_3387_;
	assign _3389_ = ~(_3388_ ^ _3385_);
	assign _3390_ = _3389_ ^ _3384_;
	assign _3391_ = ~(_3375_ ^ _3374_);
	assign _3392_ = _3391_ & _3390_;
	assign _3393_ = ~(_3392_ | _3376_);
	assign _3394_ = _3344_ ^ _3343_;
	assign _3395_ = _3394_ & ~_3393_;
	assign _3396_ = _3385_ & ~_3388_;
	assign _3397_ = _3389_ & _3384_;
	assign _3398_ = _3397_ | _3396_;
	assign _3399_ = ~(_3394_ ^ _3393_);
	assign _3400_ = _3399_ & _3398_;
	assign _3401_ = ~(_3400_ | _3395_);
	assign _3402_ = _3352_ ^ _3351_;
	assign _3403_ = _3402_ & ~_3401_;
	assign _3404_ = _3403_ & _3357_;
	assign _3405_ = ~(_3355_ ^ _3310_);
	assign _3406_ = _3405_ & _3404_;
	assign _3407_ = _3356_ & ~_3406_;
	assign _3408_ = _3403_ ^ _3357_;
	assign _3409_ = _3408_ & _3405_;
	assign _3410_ = \mchip.value_B [0] & \mchip.value_A [8];
	assign _3411_ = \mchip.value_B [1] & \mchip.value_A [7];
	assign _3412_ = _3411_ & _3410_;
	assign _3413_ = \mchip.value_B [2] & \mchip.value_A [6];
	assign _3414_ = _3411_ ^ _3410_;
	assign _3415_ = _3414_ & _3413_;
	assign _3416_ = ~(_3415_ | _3412_);
	assign _3417_ = _3362_ ^ _3361_;
	assign _3418_ = _3417_ & ~_3416_;
	assign _3419_ = \mchip.value_B [5] & \mchip.value_A [4];
	assign _3420_ = \mchip.value_B [4] & \mchip.value_A [5];
	assign _3421_ = \mchip.value_A [6] & \mchip.value_B [3];
	assign _3422_ = _3421_ ^ _3420_;
	assign _3423_ = _3422_ ^ _3419_;
	assign _3424_ = ~(_3417_ ^ _3416_);
	assign _3425_ = _3424_ & _3423_;
	assign _3426_ = ~(_3425_ | _3418_);
	assign _3427_ = _3372_ ^ _3371_;
	assign _3428_ = _3427_ & ~_3426_;
	assign _3429_ = \mchip.value_B [6] & \mchip.value_A [3];
	assign _3430_ = \mchip.value_A [2] & \mchip.value_B [7];
	assign _3431_ = _3430_ & _3429_;
	assign _3432_ = \mchip.value_A [1] & \mchip.value_B [8];
	assign _3433_ = ~_3432_;
	assign _3434_ = _3430_ ^ _3429_;
	assign _3435_ = _3434_ & ~_3433_;
	assign _3436_ = _3435_ | _3431_;
	assign _3437_ = _3382_ ^ _3381_;
	assign _3438_ = _3421_ & _3420_;
	assign _3439_ = ~(_3422_ & _3419_);
	assign _3440_ = _3439_ & ~_3438_;
	assign _3441_ = _3440_ ^ _3437_;
	assign _3442_ = _3441_ ^ _3436_;
	assign _3443_ = ~(_3427_ ^ _3426_);
	assign _3444_ = _3443_ & _3442_;
	assign _3445_ = ~(_3444_ | _3428_);
	assign _3446_ = _3391_ ^ _3390_;
	assign _3447_ = _3446_ & ~_3445_;
	assign _3448_ = \mchip.value_A [1] & ~_1521_;
	assign _3449_ = _3440_ | _3437_;
	assign _3450_ = _3441_ & _3436_;
	assign _3451_ = _3449_ & ~_3450_;
	assign _3452_ = ~(_3451_ ^ _3448_);
	assign _3453_ = ~(_3446_ ^ _3445_);
	assign _3454_ = _3453_ & _3452_;
	assign _3455_ = ~(_3454_ | _3447_);
	assign _3456_ = _3399_ ^ _3398_;
	assign _3457_ = _3455_ | ~_3456_;
	assign _3458_ = _3448_ & ~_3451_;
	assign _3459_ = ~(_3456_ ^ _3455_);
	assign _3460_ = _3459_ & _3458_;
	assign _3461_ = _3457_ & ~_3460_;
	assign _3462_ = ~(_3402_ ^ _3401_);
	assign _3463_ = _3461_ | ~_3462_;
	assign _3464_ = \mchip.value_B [0] & \mchip.value_A [7];
	assign _3465_ = \mchip.value_B [1] & \mchip.value_A [6];
	assign _3466_ = _3465_ & _3464_;
	assign _3467_ = \mchip.value_B [2] & \mchip.value_A [5];
	assign _3468_ = _3465_ ^ _3464_;
	assign _3469_ = _3468_ & _3467_;
	assign _3470_ = ~(_3469_ | _3466_);
	assign _3471_ = _3414_ ^ _3413_;
	assign _3472_ = _3471_ & ~_3470_;
	assign _3473_ = \mchip.value_A [3] & \mchip.value_B [5];
	assign _3474_ = \mchip.value_A [4] & \mchip.value_B [4];
	assign _3475_ = \mchip.value_A [5] & \mchip.value_B [3];
	assign _3476_ = _3475_ ^ _3474_;
	assign _3477_ = _3476_ ^ _3473_;
	assign _3478_ = ~(_3471_ ^ _3470_);
	assign _3479_ = _3478_ & _3477_;
	assign _3480_ = ~(_3479_ | _3472_);
	assign _3481_ = _3424_ ^ _3423_;
	assign _3482_ = _3481_ & ~_3480_;
	assign _3483_ = \mchip.value_A [2] & \mchip.value_B [6];
	assign _3484_ = \mchip.value_B [7] & \mchip.value_A [1];
	assign _3485_ = _3484_ & _3483_;
	assign _3486_ = \mchip.value_A [0] & \mchip.value_B [8];
	assign _3487_ = ~_3486_;
	assign _3488_ = _3484_ ^ _3483_;
	assign _3489_ = _3488_ & ~_3487_;
	assign _3490_ = _3489_ | _3485_;
	assign _3491_ = _3434_ ^ _3433_;
	assign _3492_ = _3475_ & _3474_;
	assign _3493_ = ~(_3476_ & _3473_);
	assign _3494_ = _3493_ & ~_3492_;
	assign _3495_ = _3494_ ^ _3491_;
	assign _3496_ = _3495_ ^ _3490_;
	assign _3497_ = ~(_3481_ ^ _3480_);
	assign _3498_ = _3497_ & _3496_;
	assign _3499_ = ~(_3498_ | _3482_);
	assign _3500_ = _3443_ ^ _3442_;
	assign _3501_ = _3500_ & ~_3499_;
	assign _3502_ = \mchip.value_A [0] & ~_1521_;
	assign _3503_ = \mchip.value_B [9] & \mchip.value_A [1];
	assign _3504_ = _3494_ | _3491_;
	assign _3505_ = _3495_ & _3490_;
	assign _3506_ = _3504_ & ~_3505_;
	assign _3507_ = ~(_3506_ ^ _3503_);
	assign _3508_ = _3507_ ^ _3502_;
	assign _3509_ = ~(_3500_ ^ _3499_);
	assign _3510_ = _3509_ & _3508_;
	assign _3511_ = ~(_3510_ | _3501_);
	assign _3512_ = _3453_ ^ _3452_;
	assign _3513_ = _3512_ & ~_3511_;
	assign _3514_ = _3503_ & ~_3506_;
	assign _3515_ = _3507_ & _3502_;
	assign _3516_ = _3515_ | _3514_;
	assign _3517_ = ~(_3512_ ^ _3511_);
	assign _3518_ = _3517_ & _3516_;
	assign _3519_ = ~(_3518_ | _3513_);
	assign _3520_ = _3459_ ^ _3458_;
	assign _3521_ = _3520_ & ~_3519_;
	assign _3522_ = ~_3521_;
	assign _3523_ = ~(_3462_ ^ _3461_);
	assign _3524_ = _3523_ & ~_3522_;
	assign _3525_ = _3463_ & ~_3524_;
	assign _3526_ = _3409_ & ~_3525_;
	assign _3527_ = _3407_ & ~_3526_;
	assign _3528_ = _3520_ ^ _3519_;
	assign _3529_ = _3523_ & ~_3528_;
	assign _3530_ = _3529_ & _3409_;
	assign _3531_ = \mchip.value_B [0] & \mchip.value_A [6];
	assign _3532_ = \mchip.value_B [1] & \mchip.value_A [5];
	assign _3533_ = _3532_ & _3531_;
	assign _3534_ = \mchip.value_B [2] & \mchip.value_A [4];
	assign _3535_ = _3532_ ^ _3531_;
	assign _3536_ = _3535_ & _3534_;
	assign _3537_ = ~(_3536_ | _3533_);
	assign _3538_ = _3468_ ^ _3467_;
	assign _3539_ = _3538_ & ~_3537_;
	assign _3540_ = \mchip.value_A [2] & \mchip.value_B [5];
	assign _3541_ = \mchip.value_A [3] & \mchip.value_B [4];
	assign _3542_ = \mchip.value_A [4] & \mchip.value_B [3];
	assign _3543_ = _3542_ ^ _3541_;
	assign _3544_ = _3543_ ^ _3540_;
	assign _3545_ = ~(_3538_ ^ _3537_);
	assign _3546_ = _3545_ & _3544_;
	assign _3547_ = ~(_3546_ | _3539_);
	assign _3548_ = _3478_ ^ _3477_;
	assign _3549_ = _3548_ & ~_3547_;
	assign _3550_ = \mchip.value_A [0] & \mchip.value_B [7];
	assign _3551_ = \mchip.value_B [6] & \mchip.value_A [1];
	assign _3552_ = _3551_ & _3550_;
	assign _3553_ = _3488_ ^ _3487_;
	assign _3554_ = _3542_ & _3541_;
	assign _3555_ = ~(_3543_ & _3540_);
	assign _3556_ = _3555_ & ~_3554_;
	assign _3557_ = _3556_ ^ _3553_;
	assign _3558_ = _3557_ ^ _3552_;
	assign _3559_ = ~(_3548_ ^ _3547_);
	assign _3560_ = _3559_ & _3558_;
	assign _3561_ = ~(_3560_ | _3549_);
	assign _3562_ = _3497_ ^ _3496_;
	assign _3563_ = _3562_ & ~_3561_;
	assign _3564_ = \mchip.value_B [9] & \mchip.value_A [0];
	assign _3565_ = _3556_ | _3553_;
	assign _3566_ = _3557_ & _3552_;
	assign _3567_ = _3565_ & ~_3566_;
	assign _3568_ = ~(_3567_ ^ _3564_);
	assign _3569_ = ~(_3562_ ^ _3561_);
	assign _3570_ = _3569_ & _3568_;
	assign _3571_ = ~(_3570_ | _3563_);
	assign _3572_ = _3509_ ^ _3508_;
	assign _3573_ = _3571_ | ~_3572_;
	assign _3574_ = _3564_ & ~_3567_;
	assign _3575_ = ~(_3572_ ^ _3571_);
	assign _3576_ = _3575_ & _3574_;
	assign _3577_ = _3573_ & ~_3576_;
	assign _3578_ = _3517_ ^ _3516_;
	assign _3579_ = _3577_ | ~_3578_;
	assign _3580_ = _3575_ ^ _3574_;
	assign _3581_ = _3569_ ^ _3568_;
	assign _3582_ = \mchip.value_B [0] & \mchip.value_A [5];
	assign _3583_ = \mchip.value_B [1] & \mchip.value_A [4];
	assign _3584_ = _3583_ & _3582_;
	assign _3585_ = \mchip.value_B [2] & \mchip.value_A [3];
	assign _3586_ = _3583_ ^ _3582_;
	assign _3587_ = _3586_ & _3585_;
	assign _3588_ = ~(_3587_ | _3584_);
	assign _3589_ = _3535_ ^ _3534_;
	assign _3590_ = _3589_ & ~_3588_;
	assign _3591_ = \mchip.value_A [1] & \mchip.value_B [5];
	assign _3592_ = \mchip.value_A [2] & \mchip.value_B [4];
	assign _3593_ = \mchip.value_A [3] & \mchip.value_B [3];
	assign _3594_ = _3593_ ^ _3592_;
	assign _3595_ = _3594_ ^ _3591_;
	assign _3596_ = ~(_3589_ ^ _3588_);
	assign _3597_ = _3596_ & _3595_;
	assign _3598_ = ~(_3597_ | _3590_);
	assign _3599_ = _3545_ ^ _3544_;
	assign _3600_ = _3598_ | ~_3599_;
	assign _3601_ = _3551_ ^ _3550_;
	assign _3602_ = _3593_ & _3592_;
	assign _3603_ = ~(_3594_ & _3591_);
	assign _3604_ = _3603_ & ~_3602_;
	assign _3605_ = ~(_3604_ ^ _3601_);
	assign _3606_ = ~(_3599_ ^ _3598_);
	assign _3607_ = _3606_ & _3605_;
	assign _3608_ = _3600_ & ~_3607_;
	assign _3609_ = _3559_ ^ _3558_;
	assign _3610_ = _3608_ | ~_3609_;
	assign _3611_ = _3601_ & ~_3604_;
	assign _3612_ = ~(_3609_ ^ _3608_);
	assign _3613_ = _3612_ & _3611_;
	assign _3614_ = _3610_ & ~_3613_;
	assign _3615_ = _3581_ & ~_3614_;
	assign _3616_ = _3615_ & _3580_;
	assign _3617_ = ~_3616_;
	assign _3618_ = ~(_3578_ ^ _3577_);
	assign _3619_ = _3618_ & ~_3617_;
	assign _3620_ = _3579_ & ~_3619_;
	assign _3621_ = ~(_3615_ ^ _3580_);
	assign _3622_ = _3618_ & ~_3621_;
	assign _3623_ = _3614_ ^ _3581_;
	assign _3624_ = _3612_ ^ _3611_;
	assign _3625_ = \mchip.value_B [0] & \mchip.value_A [4];
	assign _3626_ = \mchip.value_B [1] & \mchip.value_A [3];
	assign _3627_ = _3626_ & _3625_;
	assign _3628_ = \mchip.value_B [2] & \mchip.value_A [2];
	assign _3629_ = _3626_ ^ _3625_;
	assign _3630_ = _3629_ & _3628_;
	assign _3631_ = ~(_3630_ | _3627_);
	assign _3632_ = _3586_ ^ _3585_;
	assign _3633_ = _3632_ & ~_3631_;
	assign _3634_ = \mchip.value_A [0] & \mchip.value_B [5];
	assign _3635_ = \mchip.value_A [1] & \mchip.value_B [4];
	assign _3636_ = \mchip.value_A [2] & \mchip.value_B [3];
	assign _3637_ = _3636_ ^ _3635_;
	assign _3638_ = _3637_ ^ _3634_;
	assign _3639_ = ~(_3632_ ^ _3631_);
	assign _3640_ = _3639_ & _3638_;
	assign _3641_ = ~(_3640_ | _3633_);
	assign _3642_ = _3596_ ^ _3595_;
	assign _3643_ = _3641_ | ~_3642_;
	assign _3644_ = \mchip.value_A [0] & \mchip.value_B [6];
	assign _3645_ = _3636_ & _3635_;
	assign _3646_ = ~(_3637_ & _3634_);
	assign _3647_ = _3646_ & ~_3645_;
	assign _3648_ = ~(_3647_ ^ _3644_);
	assign _3649_ = ~(_3642_ ^ _3641_);
	assign _3650_ = _3649_ & _3648_;
	assign _3651_ = _3643_ & ~_3650_;
	assign _3652_ = _3606_ ^ _3605_;
	assign _3653_ = _3651_ | ~_3652_;
	assign _3654_ = _3644_ & ~_3647_;
	assign _3655_ = ~(_3652_ ^ _3651_);
	assign _3656_ = _3655_ & _3654_;
	assign _3657_ = _3653_ & ~_3656_;
	assign _3658_ = _3624_ & ~_3657_;
	assign _3659_ = _3623_ | ~_3658_;
	assign _3660_ = ~(_3657_ ^ _3624_);
	assign _3661_ = _3649_ ^ _3648_;
	assign _3662_ = \mchip.value_B [0] & \mchip.value_A [3];
	assign _3663_ = \mchip.value_B [1] & \mchip.value_A [2];
	assign _3664_ = _3663_ & _3662_;
	assign _3665_ = \mchip.value_B [2] & \mchip.value_A [1];
	assign _3666_ = _3663_ ^ _3662_;
	assign _3667_ = _3666_ & _3665_;
	assign _3668_ = ~(_3667_ | _3664_);
	assign _3669_ = _3629_ ^ _3628_;
	assign _3670_ = _3669_ & ~_3668_;
	assign _3671_ = \mchip.value_A [0] & \mchip.value_B [4];
	assign _3672_ = \mchip.value_A [1] & \mchip.value_B [3];
	assign _3673_ = _3672_ ^ _3671_;
	assign _3674_ = ~(_3669_ ^ _3668_);
	assign _3675_ = _3674_ & _3673_;
	assign _3676_ = ~(_3675_ | _3670_);
	assign _3677_ = _3639_ ^ _3638_;
	assign _3678_ = _3676_ | ~_3677_;
	assign _3679_ = _3672_ & _3671_;
	assign _3680_ = ~(_3677_ ^ _3676_);
	assign _3681_ = _3680_ & _3679_;
	assign _3682_ = _3678_ & ~_3681_;
	assign _3683_ = _3661_ & ~_3682_;
	assign _3684_ = _3655_ ^ _3654_;
	assign _3685_ = _3684_ & _3683_;
	assign _3686_ = _3685_ & _3660_;
	assign _3687_ = ~(_3658_ ^ _3623_);
	assign _3688_ = _3687_ & _3686_;
	assign _3689_ = _3659_ & ~_3688_;
	assign _3690_ = _3622_ & ~_3689_;
	assign _3691_ = _3620_ & ~_3690_;
	assign _3692_ = _3530_ & ~_3691_;
	assign _3693_ = _3527_ & ~_3692_;
	assign _3694_ = ~(_3685_ ^ _3660_);
	assign _3695_ = _3694_ | ~_3687_;
	assign _3696_ = _3622_ & ~_3695_;
	assign _3697_ = _3696_ & _3530_;
	assign _3698_ = _3684_ ^ _3683_;
	assign _3699_ = _3674_ ^ _3673_;
	assign _3700_ = \mchip.value_B [0] & \mchip.value_A [2];
	assign _3701_ = \mchip.value_B [1] & \mchip.value_A [1];
	assign _3702_ = _3701_ & _3700_;
	assign _3703_ = \mchip.value_B [2] & \mchip.value_A [0];
	assign _3704_ = _3701_ ^ _3700_;
	assign _3705_ = _3704_ & _3703_;
	assign _3706_ = ~(_3705_ | _3702_);
	assign _3707_ = _3666_ ^ _3665_;
	assign _3708_ = _3706_ | ~_3707_;
	assign _3709_ = \mchip.value_A [0] & \mchip.value_B [3];
	assign _3710_ = ~(_3707_ ^ _3706_);
	assign _3711_ = _3710_ & _3709_;
	assign _3712_ = _3708_ & ~_3711_;
	assign _3713_ = _3699_ & ~_3712_;
	assign _3714_ = ~_3713_;
	assign _3715_ = _3680_ ^ _3679_;
	assign _3716_ = _3715_ & ~_3714_;
	assign _3717_ = ~(_3682_ ^ _3661_);
	assign _3718_ = _3717_ & _3716_;
	assign _3719_ = ~(_3718_ & _3698_);
	assign _3720_ = \mchip.value_B [1] & \mchip.value_A [0];
	assign _3721_ = \mchip.value_B [0] & \mchip.value_A [1];
	assign _3722_ = _3721_ & _3720_;
	assign _3723_ = ~_3722_;
	assign _3724_ = _3704_ ^ _3703_;
	assign _3725_ = _3724_ & ~_3723_;
	assign _3726_ = ~_3725_;
	assign _3727_ = _3710_ ^ _3709_;
	assign _3728_ = _3727_ & ~_3726_;
	assign _3729_ = ~_3728_;
	assign _3730_ = ~(_3712_ ^ _3699_);
	assign _3731_ = _3730_ & ~_3729_;
	assign _3732_ = ~_3731_;
	assign _3733_ = _3715_ ^ _3713_;
	assign _3734_ = _3733_ & ~_3732_;
	assign _3735_ = ~_3734_;
	assign _3736_ = _3717_ ^ _3716_;
	assign _3737_ = _3736_ & ~_3735_;
	assign _3738_ = _3718_ ^ _3698_;
	assign _3739_ = _3738_ & _3737_;
	assign _3740_ = _3719_ & ~_3739_;
	assign _3741_ = _3697_ & ~_3740_;
	assign _3742_ = _3693_ & ~_3741_;
	assign _3743_ = _3309_ & ~_3742_;
	assign _3744_ = _3743_ | _3306_;
	assign _3745_ = _3083_ & _2967_;
	assign _3746_ = _3073_ & _2977_;
	assign _3747_ = _3063_ & _2987_;
	assign _3748_ = _3053_ & ~_3025_;
	assign _3749_ = _3043_ & _3034_;
	assign _3750_ = ~(_1642_ | _1521_);
	assign _3751_ = _3750_ ^ _3749_;
	assign _3752_ = _3751_ ^ _3748_;
	assign _3753_ = _3752_ ^ _3747_;
	assign _3754_ = _3753_ ^ _3746_;
	assign _3755_ = _3754_ ^ _3745_;
	assign _3756_ = _3755_ ^ _3744_;
	assign _0071_ = _3754_ & _3745_;
	assign _0072_ = _3755_ & _3744_;
	assign _0073_ = ~(_0072_ | _0071_);
	assign _0074_ = _3753_ & _3746_;
	assign _0075_ = _3752_ & _3747_;
	assign _0076_ = _3750_ & _3749_;
	assign _0077_ = _3751_ & _3748_;
	assign _0078_ = _0077_ ^ _0076_;
	assign _0079_ = _0078_ ^ _0075_;
	assign _0080_ = _0079_ ^ _0074_;
	assign _0081_ = ~(_0080_ ^ _0073_);
	assign _0082_ = ~(_1994_ & _1983_);
	assign _0083_ = _0082_ & ~_1895_;
	assign _0084_ = ~(_0083_ ^ _1906_);
	assign _0085_ = _1994_ ^ _1983_;
	assign _0086_ = ~(_1972_ ^ _1961_);
	assign _0087_ = ~(_1950_ ^ _1939_);
	assign _0088_ = ~_0087_;
	assign _0089_ = _0088_ & ~_0086_;
	assign _0090_ = _0089_ & ~_0085_;
	assign _0091_ = ~(_0084_ ^ _0090_);
	assign _0092_ = (_2137_ ? _0084_ : _0091_);
	assign _0093_ = ~(_0089_ ^ _0085_);
	assign _0094_ = (_2137_ ? _0085_ : _0093_);
	assign _0095_ = _0094_ | _0092_;
	assign _0096_ = _0087_ ^ _0086_;
	assign _0097_ = (_2137_ ? _0086_ : _0096_);
	assign _0098_ = _0097_ | _0088_;
	assign _0099_ = ~(_0098_ | _0095_);
	assign _0100_ = _0084_ | _0085_;
	assign _0101_ = _0089_ & ~_0100_;
	assign _0102_ = _2038_ ^ _2027_;
	assign _0103_ = _0102_ | ~_0101_;
	assign _0104_ = _0103_ ^ _2093_;
	assign _0105_ = (_2137_ ? _2093_ : _0104_);
	assign _0106_ = ~(_0102_ ^ _0101_);
	assign _0107_ = (_2137_ ? _0102_ : _0106_);
	assign _0108_ = _0107_ | _0105_;
	assign _0109_ = _0099_ & ~_0108_;
	assign _0110_ = _0109_ & _0081_;
	assign _0111_ = _0097_ | _0087_;
	assign _0112_ = _0111_ | _0095_;
	assign _0113_ = ~(_0112_ | _0108_);
	assign _0114_ = _3756_ & _0113_;
	assign _0115_ = ~(_0114_ | _0110_);
	assign _0116_ = ~(_0094_ & _0092_);
	assign _0117_ = ~(_0097_ & _0088_);
	assign _0118_ = _0117_ | _0116_;
	assign _0119_ = ~(_0118_ | _0108_);
	assign _0120_ = ~(_0097_ & _0087_);
	assign _0121_ = _0120_ | _0116_;
	assign _0122_ = ~(_0121_ | _0108_);
	assign _0123_ = ~(_0122_ | _0119_);
	assign _0124_ = _0116_ | _0111_;
	assign _0125_ = ~(_0124_ | _0108_);
	assign _0126_ = _0116_ | _0098_;
	assign _0127_ = ~(_0126_ | _0108_);
	assign _0128_ = _0127_ | _0125_;
	assign _0129_ = _0123_ & ~_0128_;
	assign _0130_ = _0094_ | ~_0092_;
	assign _0131_ = _0130_ | _0111_;
	assign _0132_ = ~(_0131_ | _0108_);
	assign _0133_ = _0130_ | _0098_;
	assign _0134_ = ~(_0133_ | _0108_);
	assign _0135_ = _0134_ | _0132_;
	assign _0136_ = _0130_ | _0117_;
	assign _0137_ = ~(_0136_ | _0108_);
	assign _0138_ = _0130_ | _0120_;
	assign _0139_ = ~(_0138_ | _0108_);
	assign _0140_ = _0139_ | _0137_;
	assign _0141_ = _0140_ | _0135_;
	assign _0142_ = _0129_ & ~_0141_;
	assign _0143_ = _0113_ | _0109_;
	assign _0144_ = _0117_ | _0095_;
	assign _0145_ = ~(_0144_ | _0108_);
	assign _0146_ = _0120_ | _0095_;
	assign _0147_ = ~(_0146_ | _0108_);
	assign _0148_ = _0147_ | _0145_;
	assign _0149_ = _0148_ | _0143_;
	assign _0150_ = _0092_ | ~_0094_;
	assign _0151_ = _0150_ | _0111_;
	assign _0152_ = ~(_0151_ | _0108_);
	assign _0153_ = _0150_ | _0098_;
	assign _0154_ = ~(_0153_ | _0108_);
	assign _0155_ = _0154_ | _0152_;
	assign _0156_ = _0150_ | _0117_;
	assign _0157_ = ~(_0156_ | _0108_);
	assign _0158_ = _0150_ | _0120_;
	assign _0159_ = ~(_0158_ | _0108_);
	assign _0160_ = _0159_ | _0157_;
	assign _0161_ = _0160_ | _0155_;
	assign _0162_ = _0161_ | _0149_;
	assign _0163_ = _0142_ & ~_0162_;
	assign _0164_ = ~(_0163_ | _0115_);
	assign _0165_ = (_2137_ ? _3756_ : _0164_);
	assign _0166_ = ~_3210_;
	assign _0167_ = _3308_ & ~_3742_;
	assign _0168_ = _3304_ & ~_0167_;
	assign _0169_ = _0168_ | _0166_;
	assign _0170_ = _0169_ & ~_3206_;
	assign _0171_ = ~(_0170_ ^ _3207_);
	assign _0172_ = ~(_0145_ & _0081_);
	assign _0173_ = ~_0113_;
	assign _0174_ = _0171_ & ~_0173_;
	assign _0175_ = _3756_ & _0109_;
	assign _0176_ = _0175_ | _0174_;
	assign _0177_ = _0172_ & ~_0176_;
	assign _0178_ = ~(_0177_ | _0163_);
	assign _0179_ = (_2137_ ? _0171_ : _0178_);
	assign _0180_ = _0179_ | _0165_;
	assign _0181_ = _0168_ ^ _0166_;
	assign _0182_ = ~(_0147_ & _0081_);
	assign _0183_ = _0145_ & _3756_;
	assign _0184_ = _0182_ & ~_0183_;
	assign _0185_ = _0181_ & ~_0173_;
	assign _0186_ = _0171_ & _0109_;
	assign _0187_ = _0186_ | _0185_;
	assign _0188_ = _0184_ & ~_0187_;
	assign _0189_ = ~(_0188_ | _0163_);
	assign _0190_ = (_2137_ ? _0181_ : _0189_);
	assign _0191_ = _3742_ | _3307_;
	assign _0192_ = _0191_ & ~_3301_;
	assign _0193_ = ~(_0192_ ^ _3302_);
	assign _0194_ = ~(_0152_ & _0081_);
	assign _0195_ = _0193_ & ~_0173_;
	assign _0196_ = _0181_ & _0109_;
	assign _0197_ = _0196_ | _0195_;
	assign _0198_ = _0171_ & _0145_;
	assign _0199_ = _0147_ & _3756_;
	assign _0200_ = _0199_ | _0198_;
	assign _0201_ = _0200_ | _0197_;
	assign _0202_ = _0194_ & ~_0201_;
	assign _0203_ = ~(_0202_ | _0163_);
	assign _0204_ = (_2137_ ? _0193_ : _0203_);
	assign _0205_ = _0204_ | _0190_;
	assign _0206_ = _3742_ ^ _3307_;
	assign _0207_ = ~(_0154_ & _0081_);
	assign _0208_ = _0152_ & _3756_;
	assign _0209_ = _0207_ & ~_0208_;
	assign _0210_ = _0206_ & ~_0173_;
	assign _0211_ = _0193_ & _0109_;
	assign _0212_ = _0211_ | _0210_;
	assign _0213_ = _0181_ & _0145_;
	assign _0214_ = _0171_ & _0147_;
	assign _0215_ = _0214_ | _0213_;
	assign _0216_ = _0215_ | _0212_;
	assign _0217_ = _0209_ & ~_0216_;
	assign _0218_ = ~(_0217_ | _0163_);
	assign _0219_ = (_2137_ ? _0206_ : _0218_);
	assign _0220_ = ~_3408_;
	assign _0221_ = _3696_ & ~_3740_;
	assign _0222_ = _3691_ & ~_0221_;
	assign _0223_ = _3529_ & ~_0222_;
	assign _0224_ = _3525_ & ~_0223_;
	assign _0225_ = _0224_ | _0220_;
	assign _0226_ = _0225_ & ~_3404_;
	assign _0227_ = ~(_0226_ ^ _3405_);
	assign _0228_ = ~(_0157_ & _0081_);
	assign _0229_ = _0171_ & _0152_;
	assign _0230_ = _0154_ & _3756_;
	assign _0231_ = _0230_ | _0229_;
	assign _0232_ = _0228_ & ~_0231_;
	assign _0233_ = _0227_ & ~_0173_;
	assign _0234_ = _0206_ & _0109_;
	assign _0235_ = _0234_ | _0233_;
	assign _0236_ = _0193_ & _0145_;
	assign _0237_ = _0181_ & _0147_;
	assign _0238_ = _0237_ | _0236_;
	assign _0239_ = _0238_ | _0235_;
	assign _0240_ = _0232_ & ~_0239_;
	assign _0241_ = ~(_0240_ | _0163_);
	assign _0242_ = (_2137_ ? _0227_ : _0241_);
	assign _0243_ = _0242_ | _0219_;
	assign _0244_ = _0243_ | _0205_;
	assign _0245_ = _0224_ ^ _0220_;
	assign _0246_ = ~(_0159_ & _0081_);
	assign _0247_ = _0157_ & _3756_;
	assign _0248_ = _0246_ & ~_0247_;
	assign _0249_ = _0181_ & _0152_;
	assign _0250_ = _0171_ & _0154_;
	assign _0251_ = _0250_ | _0249_;
	assign _0252_ = _0248_ & ~_0251_;
	assign _0253_ = _0245_ & ~_0173_;
	assign _0254_ = _0227_ & _0109_;
	assign _0255_ = _0254_ | _0253_;
	assign _0256_ = _0206_ & _0145_;
	assign _0257_ = _0193_ & _0147_;
	assign _0258_ = _0257_ | _0256_;
	assign _0259_ = _0258_ | _0255_;
	assign _0260_ = _0252_ & ~_0259_;
	assign _0261_ = ~(_0260_ | _0163_);
	assign _0262_ = (_2137_ ? _0245_ : _0261_);
	assign _0263_ = ~(_0222_ | _3528_);
	assign _0264_ = _3522_ & ~_0263_;
	assign _0265_ = ~(_0264_ ^ _3523_);
	assign _0266_ = ~(_0132_ & _0081_);
	assign _0267_ = _0265_ & ~_0173_;
	assign _0268_ = _0245_ & _0109_;
	assign _0269_ = _0268_ | _0267_;
	assign _0270_ = _0227_ & _0145_;
	assign _0271_ = _0206_ & _0147_;
	assign _0272_ = _0271_ | _0270_;
	assign _0273_ = _0272_ | _0269_;
	assign _0274_ = _0193_ & _0152_;
	assign _0275_ = _0181_ & _0154_;
	assign _0276_ = _0275_ | _0274_;
	assign _0277_ = _0171_ & _0157_;
	assign _0278_ = _0159_ & _3756_;
	assign _0279_ = _0278_ | _0277_;
	assign _0280_ = _0279_ | _0276_;
	assign _0281_ = _0280_ | _0273_;
	assign _0282_ = _0266_ & ~_0281_;
	assign _0283_ = ~(_0282_ | _0163_);
	assign _0284_ = (_2137_ ? _0265_ : _0283_);
	assign _0285_ = _0284_ | _0262_;
	assign _0286_ = _0222_ ^ _3528_;
	assign _0287_ = ~(_0134_ & _0081_);
	assign _0288_ = _0132_ & _3756_;
	assign _0289_ = _0287_ & ~_0288_;
	assign _0290_ = _0286_ & ~_0173_;
	assign _0291_ = _0265_ & _0109_;
	assign _0292_ = _0291_ | _0290_;
	assign _0293_ = _0245_ & _0145_;
	assign _0294_ = _0227_ & _0147_;
	assign _0295_ = _0294_ | _0293_;
	assign _0296_ = _0295_ | _0292_;
	assign _0297_ = _0206_ & _0152_;
	assign _0298_ = _0193_ & _0154_;
	assign _0299_ = _0298_ | _0297_;
	assign _0300_ = _0181_ & _0157_;
	assign _0301_ = _0171_ & _0159_;
	assign _0302_ = _0301_ | _0300_;
	assign _0303_ = _0302_ | _0299_;
	assign _0304_ = _0303_ | _0296_;
	assign _0305_ = _0289_ & ~_0304_;
	assign _0306_ = ~(_0305_ | _0163_);
	assign _0307_ = (_2137_ ? _0286_ : _0306_);
	assign _0308_ = ~(_3740_ | _3695_);
	assign _0309_ = _3689_ & ~_0308_;
	assign _0310_ = ~(_0309_ | _3621_);
	assign _0311_ = _3617_ & ~_0310_;
	assign _0312_ = ~(_0311_ ^ _3618_);
	assign _0313_ = ~(_0312_ & _0113_);
	assign _0314_ = _0286_ & _0109_;
	assign _0315_ = _0313_ & ~_0314_;
	assign _0316_ = _0265_ & _0145_;
	assign _0317_ = _0245_ & _0147_;
	assign _0318_ = _0317_ | _0316_;
	assign _0319_ = _0315_ & ~_0318_;
	assign _0320_ = _0227_ & _0152_;
	assign _0321_ = _0206_ & _0154_;
	assign _0322_ = _0321_ | _0320_;
	assign _0323_ = _0193_ & _0157_;
	assign _0324_ = _0181_ & _0159_;
	assign _0325_ = _0324_ | _0323_;
	assign _0326_ = _0325_ | _0322_;
	assign _0327_ = _0319_ & ~_0326_;
	assign _0328_ = _0171_ & _0132_;
	assign _0329_ = _0134_ & _3756_;
	assign _0330_ = _0329_ | _0328_;
	assign _0331_ = _0137_ & _0081_;
	assign _0332_ = _0331_ | _0330_;
	assign _0333_ = _0327_ & ~_0332_;
	assign _0334_ = ~(_0333_ | _0163_);
	assign _0335_ = (_2137_ ? _0312_ : _0334_);
	assign _0336_ = _0335_ | _0307_;
	assign _0337_ = _0336_ | _0285_;
	assign _0338_ = _0337_ | _0244_;
	assign _0339_ = _0338_ | _0180_;
	assign _0340_ = ~(_0339_ | _2137_);
	assign _0341_ = ~_0206_;
	assign _0342_ = _0193_ & ~_0341_;
	assign _0343_ = ~(_0245_ & _0227_);
	assign _0344_ = _0342_ & ~_0343_;
	assign _0345_ = _0286_ & _0265_;
	assign _0346_ = _3740_ | _3694_;
	assign _0347_ = _0346_ & ~_3686_;
	assign _0348_ = ~(_0347_ ^ _3687_);
	assign _0349_ = _0309_ ^ _3621_;
	assign _0350_ = ~(_0349_ & _0348_);
	assign _0351_ = _0312_ & ~_0350_;
	assign _0352_ = ~(_0351_ & _0345_);
	assign _0353_ = _0344_ & ~_0352_;
	assign _0354_ = ~(_0181_ & _0171_);
	assign _0355_ = _0353_ & ~_0354_;
	assign _0356_ = ~(_0355_ ^ _3756_);
	assign _0357_ = _0355_ & _3756_;
	assign _0358_ = _0357_ ^ _0081_;
	assign _0359_ = _0358_ | ~_0356_;
	assign _0360_ = _3727_ ^ _3725_;
	assign _0361_ = ~_0360_;
	assign _0362_ = _0113_ & ~_0361_;
	assign _0363_ = _3730_ ^ _3728_;
	assign _0364_ = ~_0363_;
	assign _0365_ = _0109_ & ~_0364_;
	assign _0366_ = _0365_ | _0362_;
	assign _0367_ = _3733_ ^ _3731_;
	assign _0368_ = ~_0367_;
	assign _0369_ = _0145_ & ~_0368_;
	assign _0370_ = _3736_ ^ _3734_;
	assign _0371_ = ~_0370_;
	assign _0372_ = _0147_ & ~_0371_;
	assign _0373_ = _0372_ | _0369_;
	assign _0374_ = _0373_ | _0366_;
	assign _0375_ = _3738_ ^ _3737_;
	assign _0376_ = ~_0375_;
	assign _0377_ = _0152_ & ~_0376_;
	assign _0378_ = _3740_ ^ _3694_;
	assign _0379_ = ~_0378_;
	assign _0380_ = _0154_ & ~_0379_;
	assign _0381_ = _0380_ | _0377_;
	assign _0382_ = _0348_ & _0157_;
	assign _0383_ = _0349_ & _0159_;
	assign _0384_ = _0383_ | _0382_;
	assign _0385_ = _0384_ | _0381_;
	assign _0386_ = _0385_ | _0374_;
	assign _0387_ = _0312_ & _0132_;
	assign _0388_ = _0286_ & _0134_;
	assign _0389_ = _0388_ | _0387_;
	assign _0390_ = _0265_ & _0137_;
	assign _0391_ = _0245_ & _0139_;
	assign _0392_ = _0391_ | _0390_;
	assign _0393_ = _0392_ | _0389_;
	assign _0394_ = _0227_ & _0125_;
	assign _0395_ = _0206_ & _0127_;
	assign _0396_ = _0395_ | _0394_;
	assign _0397_ = _0193_ & _0119_;
	assign _0398_ = _0181_ & _0122_;
	assign _0399_ = _0398_ | _0397_;
	assign _0400_ = _0399_ | _0396_;
	assign _0401_ = _0400_ | _0393_;
	assign _0402_ = _0401_ | _0386_;
	assign _0403_ = (_0163_ ? _0171_ : _0402_);
	assign _0404_ = (_2137_ ? _0360_ : _0403_);
	assign _0405_ = _3724_ ^ _3722_;
	assign _0406_ = ~_0405_;
	assign _0407_ = _0113_ & ~_0406_;
	assign _0408_ = _0109_ & ~_0361_;
	assign _0409_ = _0408_ | _0407_;
	assign _0410_ = _0145_ & ~_0364_;
	assign _0411_ = _0147_ & ~_0368_;
	assign _0412_ = _0411_ | _0410_;
	assign _0413_ = _0412_ | _0409_;
	assign _0414_ = _0152_ & ~_0371_;
	assign _0415_ = _0154_ & ~_0376_;
	assign _0416_ = _0415_ | _0414_;
	assign _0417_ = _0157_ & ~_0379_;
	assign _0418_ = _0348_ & _0159_;
	assign _0419_ = _0418_ | _0417_;
	assign _0420_ = _0419_ | _0416_;
	assign _0421_ = _0420_ | _0413_;
	assign _0422_ = _0349_ & _0132_;
	assign _0423_ = _0312_ & _0134_;
	assign _0424_ = _0423_ | _0422_;
	assign _0425_ = _0286_ & _0137_;
	assign _0426_ = _0265_ & _0139_;
	assign _0427_ = _0426_ | _0425_;
	assign _0428_ = _0427_ | _0424_;
	assign _0429_ = _0245_ & _0125_;
	assign _0430_ = _0227_ & _0127_;
	assign _0431_ = _0430_ | _0429_;
	assign _0432_ = _0206_ & _0119_;
	assign _0433_ = _0193_ & _0122_;
	assign _0434_ = _0433_ | _0432_;
	assign _0435_ = _0434_ | _0431_;
	assign _0436_ = _0435_ | _0428_;
	assign _0437_ = _0436_ | _0421_;
	assign _0438_ = (_0163_ ? _0181_ : _0437_);
	assign _0439_ = (_2137_ ? _0405_ : _0438_);
	assign _0440_ = _0439_ & ~_0404_;
	assign _0441_ = ~(_0119_ & _0081_);
	assign _0442_ = _0171_ & _0125_;
	assign _0443_ = _0127_ & _3756_;
	assign _0444_ = _0443_ | _0442_;
	assign _0445_ = _0441_ & ~_0444_;
	assign _0446_ = _0227_ & _0132_;
	assign _0447_ = _0206_ & _0134_;
	assign _0448_ = _0447_ | _0446_;
	assign _0449_ = _0193_ & _0137_;
	assign _0450_ = _0181_ & _0139_;
	assign _0451_ = _0450_ | _0449_;
	assign _0452_ = _0451_ | _0448_;
	assign _0453_ = _0445_ & ~_0452_;
	assign _0454_ = _0113_ & ~_0376_;
	assign _0455_ = _0109_ & ~_0379_;
	assign _0456_ = _0455_ | _0454_;
	assign _0457_ = _0348_ & _0145_;
	assign _0458_ = _0349_ & _0147_;
	assign _0459_ = _0458_ | _0457_;
	assign _0460_ = _0459_ | _0456_;
	assign _0461_ = _0312_ & _0152_;
	assign _0462_ = _0286_ & _0154_;
	assign _0463_ = _0462_ | _0461_;
	assign _0464_ = _0265_ & _0157_;
	assign _0465_ = _0245_ & _0159_;
	assign _0466_ = _0465_ | _0464_;
	assign _0467_ = _0466_ | _0463_;
	assign _0468_ = _0467_ | _0460_;
	assign _0469_ = _0453_ & ~_0468_;
	assign _0470_ = ~(_0469_ | _0163_);
	assign _0471_ = (_2137_ ? _0375_ : _0470_);
	assign _0472_ = ~(_0122_ & _0081_);
	assign _0473_ = _0119_ & _3756_;
	assign _0474_ = _0472_ & ~_0473_;
	assign _0475_ = _0181_ & _0125_;
	assign _0476_ = _0171_ & _0127_;
	assign _0477_ = _0476_ | _0475_;
	assign _0478_ = _0474_ & ~_0477_;
	assign _0479_ = _0245_ & _0132_;
	assign _0480_ = _0227_ & _0134_;
	assign _0481_ = _0480_ | _0479_;
	assign _0482_ = _0206_ & _0137_;
	assign _0483_ = _0193_ & _0139_;
	assign _0484_ = _0483_ | _0482_;
	assign _0485_ = _0484_ | _0481_;
	assign _0486_ = _0478_ & ~_0485_;
	assign _0487_ = _0113_ & ~_0371_;
	assign _0488_ = _0109_ & ~_0376_;
	assign _0489_ = _0488_ | _0487_;
	assign _0490_ = _0145_ & ~_0379_;
	assign _0491_ = _0348_ & _0147_;
	assign _0492_ = _0491_ | _0490_;
	assign _0493_ = _0492_ | _0489_;
	assign _0494_ = _0349_ & _0152_;
	assign _0495_ = _0312_ & _0154_;
	assign _0496_ = _0495_ | _0494_;
	assign _0497_ = _0286_ & _0157_;
	assign _0498_ = _0265_ & _0159_;
	assign _0499_ = _0498_ | _0497_;
	assign _0500_ = _0499_ | _0496_;
	assign _0501_ = _0500_ | _0493_;
	assign _0502_ = _0486_ & ~_0501_;
	assign _0503_ = ~(_0502_ | _0163_);
	assign _0504_ = (_2137_ ? _0370_ : _0503_);
	assign _0505_ = _0504_ | _0471_;
	assign _0506_ = _0113_ & ~_0368_;
	assign _0507_ = _0109_ & ~_0371_;
	assign _0508_ = _0507_ | _0506_;
	assign _0509_ = _0145_ & ~_0376_;
	assign _0510_ = _0147_ & ~_0379_;
	assign _0511_ = _0510_ | _0509_;
	assign _0512_ = _0511_ | _0508_;
	assign _0513_ = _0348_ & _0152_;
	assign _0514_ = _0349_ & _0154_;
	assign _0515_ = _0514_ | _0513_;
	assign _0516_ = _0312_ & _0157_;
	assign _0517_ = _0286_ & _0159_;
	assign _0518_ = _0517_ | _0516_;
	assign _0519_ = _0518_ | _0515_;
	assign _0520_ = _0519_ | _0512_;
	assign _0521_ = _0265_ & _0132_;
	assign _0522_ = _0245_ & _0134_;
	assign _0523_ = _0522_ | _0521_;
	assign _0524_ = _0227_ & _0137_;
	assign _0525_ = _0206_ & _0139_;
	assign _0526_ = _0525_ | _0524_;
	assign _0527_ = _0526_ | _0523_;
	assign _0528_ = _0193_ & _0125_;
	assign _0529_ = _0181_ & _0127_;
	assign _0530_ = _0529_ | _0528_;
	assign _0531_ = _0171_ & _0119_;
	assign _0532_ = _0122_ & _3756_;
	assign _0533_ = _0532_ | _0531_;
	assign _0534_ = _0533_ | _0530_;
	assign _0535_ = _0534_ | _0527_;
	assign _0536_ = _0535_ | _0520_;
	assign _0537_ = (_0163_ ? _0081_ : _0536_);
	assign _0538_ = (_2137_ ? _0367_ : _0537_);
	assign _0539_ = _0113_ & ~_0364_;
	assign _0540_ = _0109_ & ~_0368_;
	assign _0541_ = _0540_ | _0539_;
	assign _0542_ = _0145_ & ~_0371_;
	assign _0543_ = _0147_ & ~_0376_;
	assign _0544_ = _0543_ | _0542_;
	assign _0545_ = _0544_ | _0541_;
	assign _0546_ = _0152_ & ~_0379_;
	assign _0547_ = _0348_ & _0154_;
	assign _0548_ = _0547_ | _0546_;
	assign _0549_ = _0349_ & _0157_;
	assign _0550_ = _0312_ & _0159_;
	assign _0551_ = _0550_ | _0549_;
	assign _0552_ = _0551_ | _0548_;
	assign _0553_ = _0552_ | _0545_;
	assign _0554_ = _0286_ & _0132_;
	assign _0555_ = _0265_ & _0134_;
	assign _0556_ = _0555_ | _0554_;
	assign _0557_ = _0245_ & _0137_;
	assign _0558_ = _0227_ & _0139_;
	assign _0559_ = _0558_ | _0557_;
	assign _0560_ = _0559_ | _0556_;
	assign _0561_ = _0206_ & _0125_;
	assign _0562_ = _0193_ & _0127_;
	assign _0563_ = _0562_ | _0561_;
	assign _0564_ = _0181_ & _0119_;
	assign _0565_ = _0171_ & _0122_;
	assign _0566_ = _0565_ | _0564_;
	assign _0567_ = _0566_ | _0563_;
	assign _0568_ = _0567_ | _0560_;
	assign _0569_ = _0568_ | _0553_;
	assign _0570_ = (_0163_ ? _3756_ : _0569_);
	assign _0571_ = (_2137_ ? _0363_ : _0570_);
	assign _0572_ = _0571_ | _0538_;
	assign _0573_ = _0572_ | _0505_;
	assign _0574_ = _0440_ & ~_0573_;
	assign _0575_ = _0262_ | _0242_;
	assign _0576_ = _0307_ | _0284_;
	assign _0577_ = _0576_ | _0575_;
	assign _0578_ = ~(_0139_ & _0081_);
	assign _0579_ = _0137_ & _3756_;
	assign _0580_ = _0578_ & ~_0579_;
	assign _0581_ = _0181_ & _0132_;
	assign _0582_ = _0171_ & _0134_;
	assign _0583_ = _0582_ | _0581_;
	assign _0584_ = _0580_ & ~_0583_;
	assign _0585_ = _0349_ & _0113_;
	assign _0586_ = _0312_ & _0109_;
	assign _0587_ = _0586_ | _0585_;
	assign _0588_ = _0286_ & _0145_;
	assign _0589_ = _0265_ & _0147_;
	assign _0590_ = _0589_ | _0588_;
	assign _0591_ = _0590_ | _0587_;
	assign _0592_ = _0245_ & _0152_;
	assign _0593_ = _0227_ & _0154_;
	assign _0594_ = _0593_ | _0592_;
	assign _0595_ = _0206_ & _0157_;
	assign _0596_ = _0193_ & _0159_;
	assign _0597_ = _0596_ | _0595_;
	assign _0598_ = _0597_ | _0594_;
	assign _0599_ = _0598_ | _0591_;
	assign _0600_ = _0584_ & ~_0599_;
	assign _0601_ = ~(_0600_ | _0163_);
	assign _0602_ = (_2137_ ? _0349_ : _0601_);
	assign _0603_ = _0602_ | _0335_;
	assign _0604_ = ~(_0125_ & _0081_);
	assign _0605_ = _0193_ & _0132_;
	assign _0606_ = _0181_ & _0134_;
	assign _0607_ = _0606_ | _0605_;
	assign _0608_ = _0171_ & _0137_;
	assign _0609_ = _0139_ & _3756_;
	assign _0610_ = _0609_ | _0608_;
	assign _0611_ = _0610_ | _0607_;
	assign _0612_ = _0604_ & ~_0611_;
	assign _0613_ = _0348_ & _0113_;
	assign _0614_ = _0349_ & _0109_;
	assign _0615_ = _0614_ | _0613_;
	assign _0616_ = _0312_ & _0145_;
	assign _0617_ = _0286_ & _0147_;
	assign _0618_ = _0617_ | _0616_;
	assign _0619_ = _0618_ | _0615_;
	assign _0620_ = _0265_ & _0152_;
	assign _0621_ = _0245_ & _0154_;
	assign _0622_ = _0621_ | _0620_;
	assign _0623_ = _0227_ & _0157_;
	assign _0624_ = _0206_ & _0159_;
	assign _0625_ = _0624_ | _0623_;
	assign _0626_ = _0625_ | _0622_;
	assign _0627_ = _0626_ | _0619_;
	assign _0628_ = _0612_ & ~_0627_;
	assign _0629_ = ~(_0628_ | _0163_);
	assign _0630_ = (_2137_ ? _0348_ : _0629_);
	assign _0631_ = ~(_0127_ & _0081_);
	assign _0632_ = _0125_ & _3756_;
	assign _0633_ = _0631_ & ~_0632_;
	assign _0634_ = _0206_ & _0132_;
	assign _0635_ = _0193_ & _0134_;
	assign _0636_ = _0635_ | _0634_;
	assign _0637_ = _0181_ & _0137_;
	assign _0638_ = _0171_ & _0139_;
	assign _0639_ = _0638_ | _0637_;
	assign _0640_ = _0639_ | _0636_;
	assign _0641_ = _0633_ & ~_0640_;
	assign _0642_ = _0113_ & ~_0379_;
	assign _0643_ = _0348_ & _0109_;
	assign _0644_ = _0643_ | _0642_;
	assign _0645_ = _0349_ & _0145_;
	assign _0646_ = _0312_ & _0147_;
	assign _0647_ = _0646_ | _0645_;
	assign _0648_ = _0647_ | _0644_;
	assign _0649_ = _0286_ & _0152_;
	assign _0650_ = _0265_ & _0154_;
	assign _0651_ = _0650_ | _0649_;
	assign _0652_ = _0245_ & _0157_;
	assign _0653_ = _0227_ & _0159_;
	assign _0654_ = _0653_ | _0652_;
	assign _0655_ = _0654_ | _0651_;
	assign _0656_ = _0655_ | _0648_;
	assign _0657_ = _0641_ & ~_0656_;
	assign _0658_ = ~(_0657_ | _0163_);
	assign _0659_ = (_2137_ ? _0378_ : _0658_);
	assign _0660_ = _0659_ | _0630_;
	assign _0661_ = _0660_ | _0603_;
	assign _0662_ = _0661_ | _0577_;
	assign _0663_ = _0574_ & ~_0662_;
	assign _0664_ = ~(_0113_ & _0081_);
	assign _0665_ = ~(_0664_ | _0163_);
	assign _0666_ = (_2137_ ? _0081_ : _0665_);
	assign _0667_ = _0666_ | _0165_;
	assign _0668_ = _0190_ | _0179_;
	assign _0669_ = _0219_ | _0204_;
	assign _0670_ = _0669_ | _0668_;
	assign _0671_ = _0670_ | _0667_;
	assign _0672_ = _0663_ & ~_0671_;
	assign _0673_ = ~(\mchip.value_B [0] & \mchip.value_A [0]);
	assign _0674_ = ~(_0227_ & _0122_);
	assign _0675_ = _0245_ & _0119_;
	assign _0676_ = _0674_ & ~_0675_;
	assign _0677_ = _0286_ & _0125_;
	assign _0678_ = _0265_ & _0127_;
	assign _0679_ = _0678_ | _0677_;
	assign _0680_ = _0676_ & ~_0679_;
	assign _0681_ = _0132_ & ~_0379_;
	assign _0682_ = _0348_ & _0134_;
	assign _0683_ = _0682_ | _0681_;
	assign _0684_ = _0349_ & _0137_;
	assign _0685_ = _0312_ & _0139_;
	assign _0686_ = _0685_ | _0684_;
	assign _0687_ = _0686_ | _0683_;
	assign _0688_ = _0680_ & ~_0687_;
	assign _0689_ = _0113_ & ~_0673_;
	assign _0690_ = _3721_ ^ _3720_;
	assign _0691_ = ~_0690_;
	assign _0692_ = _0109_ & ~_0691_;
	assign _0693_ = _0692_ | _0689_;
	assign _0694_ = _0145_ & ~_0406_;
	assign _0695_ = _0147_ & ~_0361_;
	assign _0696_ = _0695_ | _0694_;
	assign _0697_ = _0696_ | _0693_;
	assign _0698_ = _0152_ & ~_0364_;
	assign _0699_ = _0154_ & ~_0368_;
	assign _0700_ = _0699_ | _0698_;
	assign _0701_ = _0157_ & ~_0371_;
	assign _0702_ = _0159_ & ~_0376_;
	assign _0703_ = _0702_ | _0701_;
	assign _0704_ = _0703_ | _0700_;
	assign _0705_ = _0704_ | _0697_;
	assign _0706_ = _0688_ & ~_0705_;
	assign _0707_ = (_0163_ ? _0341_ : _0706_);
	assign _0708_ = (_2137_ ? _0673_ : _0707_);
	assign _0709_ = _0672_ & ~_0708_;
	assign _0710_ = _0538_ | ~_0571_;
	assign _0711_ = _0710_ | _0505_;
	assign _0712_ = _0711_ | _0662_;
	assign _0713_ = _0712_ | _0671_;
	assign _0714_ = _0439_ & ~_0713_;
	assign _0715_ = _0113_ & ~_0691_;
	assign _0716_ = _0109_ & ~_0406_;
	assign _0717_ = _0716_ | _0715_;
	assign _0718_ = _0145_ & ~_0361_;
	assign _0719_ = _0147_ & ~_0364_;
	assign _0720_ = _0719_ | _0718_;
	assign _0721_ = _0720_ | _0717_;
	assign _0722_ = _0152_ & ~_0368_;
	assign _0723_ = _0154_ & ~_0371_;
	assign _0724_ = _0723_ | _0722_;
	assign _0725_ = _0157_ & ~_0376_;
	assign _0726_ = _0159_ & ~_0379_;
	assign _0727_ = _0726_ | _0725_;
	assign _0728_ = _0727_ | _0724_;
	assign _0729_ = _0728_ | _0721_;
	assign _0730_ = _0348_ & _0132_;
	assign _0731_ = _0349_ & _0134_;
	assign _0732_ = _0731_ | _0730_;
	assign _0733_ = _0312_ & _0137_;
	assign _0734_ = _0286_ & _0139_;
	assign _0735_ = _0734_ | _0733_;
	assign _0736_ = _0735_ | _0732_;
	assign _0737_ = _0265_ & _0125_;
	assign _0738_ = _0245_ & _0127_;
	assign _0739_ = _0738_ | _0737_;
	assign _0740_ = _0227_ & _0119_;
	assign _0741_ = _0206_ & _0122_;
	assign _0742_ = _0741_ | _0740_;
	assign _0743_ = _0742_ | _0739_;
	assign _0744_ = _0743_ | _0736_;
	assign _0745_ = _0744_ | _0729_;
	assign _0746_ = (_0163_ ? _0193_ : _0745_);
	assign _0747_ = (_2137_ ? _0690_ : _0746_);
	assign _0748_ = _0573_ | ~_0404_;
	assign _0749_ = _0748_ | _0662_;
	assign _0750_ = _0749_ | _0671_;
	assign _0751_ = _0747_ & ~_0750_;
	assign _0752_ = _0751_ | _0714_;
	assign _0753_ = ~(_0752_ | _0709_);
	assign _0754_ = _0630_ | ~_0659_;
	assign _0755_ = _0754_ | _0603_;
	assign _0756_ = _0755_ | _0577_;
	assign _0757_ = _0756_ | _0671_;
	assign _0758_ = _0504_ & ~_0757_;
	assign _0759_ = _0662_ | ~_0471_;
	assign _0760_ = _0759_ | _0671_;
	assign _0761_ = _0538_ & ~_0760_;
	assign _0762_ = _0761_ | _0758_;
	assign _0763_ = _0471_ | ~_0504_;
	assign _0764_ = _0763_ | _0662_;
	assign _0765_ = _0764_ | _0671_;
	assign _0766_ = _0571_ & ~_0765_;
	assign _0767_ = _0505_ | ~_0538_;
	assign _0768_ = _0767_ | _0662_;
	assign _0769_ = _0768_ | _0671_;
	assign _0770_ = _0404_ & ~_0769_;
	assign _0771_ = _0770_ | _0766_;
	assign _0772_ = _0771_ | _0762_;
	assign _0773_ = _0753_ & ~_0772_;
	assign _0774_ = _0204_ | ~_0219_;
	assign _0775_ = _0774_ | _0668_;
	assign _0776_ = _0775_ | _0667_;
	assign _0777_ = _0262_ & ~_0776_;
	assign _0778_ = _0671_ | ~_0242_;
	assign _0779_ = _0284_ & ~_0778_;
	assign _0780_ = _0779_ | _0777_;
	assign _0781_ = _0242_ | ~_0262_;
	assign _0782_ = _0781_ | _0671_;
	assign _0783_ = _0307_ & ~_0782_;
	assign _0784_ = _0575_ | ~_0284_;
	assign _0785_ = _0784_ | _0671_;
	assign _0786_ = _0335_ & ~_0785_;
	assign _0787_ = _0786_ | _0783_;
	assign _0788_ = _0787_ | _0780_;
	assign _0789_ = _0284_ | ~_0307_;
	assign _0790_ = _0789_ | _0575_;
	assign _0791_ = _0790_ | _0671_;
	assign _0792_ = _0602_ & ~_0791_;
	assign _0793_ = _0577_ | ~_0335_;
	assign _0794_ = _0793_ | _0671_;
	assign _0795_ = _0630_ & ~_0794_;
	assign _0796_ = _0795_ | _0792_;
	assign _0797_ = _0335_ | ~_0602_;
	assign _0798_ = _0797_ | _0577_;
	assign _0799_ = _0798_ | _0671_;
	assign _0800_ = _0659_ & ~_0799_;
	assign _0801_ = _0603_ | ~_0630_;
	assign _0802_ = _0801_ | _0577_;
	assign _0803_ = _0802_ | _0671_;
	assign _0804_ = _0471_ & ~_0803_;
	assign _0805_ = _0804_ | _0800_;
	assign _0806_ = _0805_ | _0796_;
	assign _0807_ = _0806_ | _0788_;
	assign _0808_ = _0773_ & ~_0807_;
	assign _0809_ = _0667_ | ~_0179_;
	assign _0810_ = _0204_ & ~_0809_;
	assign _0811_ = _0179_ | ~_0190_;
	assign _0812_ = _0811_ | _0667_;
	assign _0813_ = _0219_ & ~_0812_;
	assign _0814_ = _0668_ | ~_0204_;
	assign _0815_ = _0814_ | _0667_;
	assign _0816_ = _0242_ & ~_0815_;
	assign _0817_ = _0816_ | _0813_;
	assign _0818_ = _0817_ | _0810_;
	assign _0819_ = _0808_ & ~_0818_;
	assign _0820_ = _0760_ & _0757_;
	assign _0821_ = ~(_0769_ & _0765_);
	assign _0822_ = _0820_ & ~_0821_;
	assign _0823_ = ~(_0750_ & _0713_);
	assign _0824_ = _0439_ | _0404_;
	assign _0825_ = _0824_ | ~_0747_;
	assign _0826_ = _0825_ | _0573_;
	assign _0827_ = _0826_ | _0662_;
	assign _0828_ = ~(_0827_ | _0671_);
	assign _0829_ = _0828_ | _0672_;
	assign _0830_ = _0829_ | _0823_;
	assign _0831_ = _0822_ & ~_0830_;
	assign _0832_ = ~(_0778_ & _0776_);
	assign _0833_ = ~(_0785_ & _0782_);
	assign _0834_ = _0833_ | _0832_;
	assign _0835_ = ~(_0794_ & _0791_);
	assign _0836_ = ~(_0803_ & _0799_);
	assign _0837_ = _0836_ | _0835_;
	assign _0838_ = _0837_ | _0834_;
	assign _0839_ = _0831_ & ~_0838_;
	assign _0840_ = _0815_ & _0812_;
	assign _0841_ = ~(_0840_ & _0809_);
	assign _0842_ = _0839_ & ~_0841_;
	assign _0843_ = ~(_0842_ | _0819_);
	assign _0844_ = _0708_ | ~_0828_;
	assign _0845_ = _0747_ & _0672_;
	assign _0846_ = _0844_ & ~_0845_;
	assign _0847_ = _0404_ & ~_0713_;
	assign _0848_ = _0439_ & ~_0750_;
	assign _0849_ = _0848_ | _0847_;
	assign _0850_ = _0846_ & ~_0849_;
	assign _0851_ = _0471_ & ~_0757_;
	assign _0852_ = _0504_ & ~_0760_;
	assign _0853_ = _0852_ | _0851_;
	assign _0854_ = _0538_ & ~_0765_;
	assign _0855_ = _0571_ & ~_0769_;
	assign _0856_ = _0855_ | _0854_;
	assign _0857_ = _0856_ | _0853_;
	assign _0858_ = _0850_ & ~_0857_;
	assign _0859_ = _0242_ & ~_0776_;
	assign _0860_ = _0262_ & ~_0778_;
	assign _0861_ = _0860_ | _0859_;
	assign _0862_ = _0284_ & ~_0782_;
	assign _0863_ = _0307_ & ~_0785_;
	assign _0864_ = _0863_ | _0862_;
	assign _0865_ = _0864_ | _0861_;
	assign _0866_ = _0335_ & ~_0791_;
	assign _0867_ = _0602_ & ~_0794_;
	assign _0868_ = _0867_ | _0866_;
	assign _0869_ = _0630_ & ~_0799_;
	assign _0870_ = _0659_ & ~_0803_;
	assign _0871_ = _0870_ | _0869_;
	assign _0872_ = _0871_ | _0868_;
	assign _0873_ = _0872_ | _0865_;
	assign _0874_ = _0858_ & ~_0873_;
	assign _0875_ = _0190_ & ~_0809_;
	assign _0876_ = _0204_ & ~_0812_;
	assign _0877_ = _0219_ & ~_0815_;
	assign _0878_ = _0877_ | _0876_;
	assign _0879_ = _0878_ | _0875_;
	assign _0880_ = _0874_ & ~_0879_;
	assign _0881_ = _0880_ | _0842_;
	assign _0882_ = _0843_ | ~_0881_;
	assign _0883_ = _0713_ | _0708_;
	assign _0884_ = _0571_ & ~_0757_;
	assign _0885_ = _0404_ & ~_0760_;
	assign _0886_ = _0885_ | _0884_;
	assign _0887_ = _0439_ & ~_0765_;
	assign _0888_ = _0747_ & ~_0769_;
	assign _0889_ = _0888_ | _0887_;
	assign _0890_ = _0889_ | _0886_;
	assign _0891_ = _0883_ & ~_0890_;
	assign _0892_ = _0307_ & ~_0776_;
	assign _0893_ = _0335_ & ~_0778_;
	assign _0894_ = _0893_ | _0892_;
	assign _0895_ = _0602_ & ~_0782_;
	assign _0896_ = _0630_ & ~_0785_;
	assign _0897_ = _0896_ | _0895_;
	assign _0898_ = _0897_ | _0894_;
	assign _0899_ = _0659_ & ~_0791_;
	assign _0900_ = _0471_ & ~_0794_;
	assign _0901_ = _0900_ | _0899_;
	assign _0902_ = _0504_ & ~_0799_;
	assign _0903_ = _0538_ & ~_0803_;
	assign _0904_ = _0903_ | _0902_;
	assign _0905_ = _0904_ | _0901_;
	assign _0906_ = _0905_ | _0898_;
	assign _0907_ = _0891_ & ~_0906_;
	assign _0908_ = _0242_ & ~_0809_;
	assign _0909_ = _0262_ & ~_0812_;
	assign _0910_ = _0284_ & ~_0815_;
	assign _0911_ = _0910_ | _0909_;
	assign _0912_ = _0911_ | _0908_;
	assign _0913_ = _0907_ & ~_0912_;
	assign _0914_ = ~(_0913_ | _0842_);
	assign _0915_ = _0750_ | _0708_;
	assign _0916_ = _0747_ & ~_0713_;
	assign _0917_ = _0915_ & ~_0916_;
	assign _0918_ = _0538_ & ~_0757_;
	assign _0919_ = _0571_ & ~_0760_;
	assign _0920_ = _0919_ | _0918_;
	assign _0921_ = _0404_ & ~_0765_;
	assign _0922_ = _0439_ & ~_0769_;
	assign _0923_ = _0922_ | _0921_;
	assign _0924_ = _0923_ | _0920_;
	assign _0925_ = _0917_ & ~_0924_;
	assign _0926_ = _0284_ & ~_0776_;
	assign _0927_ = _0307_ & ~_0778_;
	assign _0928_ = _0927_ | _0926_;
	assign _0929_ = _0335_ & ~_0782_;
	assign _0930_ = _0602_ & ~_0785_;
	assign _0932_ = _0930_ | _0929_;
	assign _0933_ = _0932_ | _0928_;
	assign _0934_ = _0630_ & ~_0791_;
	assign _0935_ = _0659_ & ~_0794_;
	assign _0936_ = _0935_ | _0934_;
	assign _0937_ = _0471_ & ~_0799_;
	assign _0938_ = _0504_ & ~_0803_;
	assign _0939_ = _0938_ | _0937_;
	assign _0940_ = _0939_ | _0936_;
	assign _0941_ = _0940_ | _0933_;
	assign _0943_ = _0925_ & ~_0941_;
	assign _0944_ = _0219_ & ~_0809_;
	assign _0945_ = _0242_ & ~_0812_;
	assign _0946_ = _0262_ & ~_0815_;
	assign _0947_ = _0946_ | _0945_;
	assign _0948_ = _0947_ | _0944_;
	assign _0949_ = _0943_ & ~_0948_;
	assign _0950_ = ~(_0949_ | _0842_);
	assign _0951_ = _0950_ | _0914_;
	assign _0952_ = _0765_ | _0708_;
	assign _0953_ = _0439_ & ~_0757_;
	assign _0954_ = _0747_ & ~_0760_;
	assign _0955_ = _0954_ | _0953_;
	assign _0956_ = _0952_ & ~_0955_;
	assign _0957_ = _0602_ & ~_0776_;
	assign _0958_ = _0630_ & ~_0778_;
	assign _0959_ = _0958_ | _0957_;
	assign _0960_ = _0659_ & ~_0782_;
	assign _0961_ = _0471_ & ~_0785_;
	assign _0962_ = _0961_ | _0960_;
	assign _0964_ = _0962_ | _0959_;
	assign _0965_ = _0504_ & ~_0791_;
	assign _0966_ = _0538_ & ~_0794_;
	assign _0967_ = _0966_ | _0965_;
	assign _0968_ = _0571_ & ~_0799_;
	assign _0969_ = _0404_ & ~_0803_;
	assign _0970_ = _0969_ | _0968_;
	assign _0971_ = _0970_ | _0967_;
	assign _0972_ = _0971_ | _0964_;
	assign _0973_ = _0956_ & ~_0972_;
	assign _0975_ = _0284_ & ~_0809_;
	assign _0976_ = _0307_ & ~_0812_;
	assign _0977_ = _0335_ & ~_0815_;
	assign _0978_ = _0977_ | _0976_;
	assign _0979_ = _0978_ | _0975_;
	assign _0980_ = _0973_ & ~_0979_;
	assign _0981_ = ~(_0980_ | _0842_);
	assign _0982_ = _0769_ | _0708_;
	assign _0983_ = _0747_ & ~_0765_;
	assign _0984_ = _0982_ & ~_0983_;
	assign _0986_ = _0404_ & ~_0757_;
	assign _0987_ = _0439_ & ~_0760_;
	assign _0988_ = _0987_ | _0986_;
	assign _0989_ = _0984_ & ~_0988_;
	assign _0990_ = _0335_ & ~_0776_;
	assign _0991_ = _0602_ & ~_0778_;
	assign _0992_ = _0991_ | _0990_;
	assign _0993_ = _0630_ & ~_0782_;
	assign _0994_ = _0659_ & ~_0785_;
	assign _0995_ = _0994_ | _0993_;
	assign _0997_ = _0995_ | _0992_;
	assign _0998_ = _0471_ & ~_0791_;
	assign _0999_ = _0504_ & ~_0794_;
	assign _1000_ = _0999_ | _0998_;
	assign _1001_ = _0538_ & ~_0799_;
	assign _1002_ = _0571_ & ~_0803_;
	assign _1003_ = _1002_ | _1001_;
	assign _1004_ = _1003_ | _1000_;
	assign _1005_ = _1004_ | _0997_;
	assign _1006_ = _0989_ & ~_1005_;
	assign _1007_ = _0262_ & ~_0809_;
	assign _1008_ = _0284_ & ~_0812_;
	assign _1009_ = _0307_ & ~_0815_;
	assign _1010_ = _1009_ | _1008_;
	assign _1011_ = _1010_ | _1007_;
	assign _1012_ = _1006_ & ~_1011_;
	assign _1013_ = ~(_1012_ | _0842_);
	assign _1014_ = _1013_ | _0981_;
	assign _1015_ = _1014_ | _0951_;
	assign _1016_ = _0757_ | _0708_;
	assign _1018_ = _0659_ & ~_0776_;
	assign _1019_ = _0471_ & ~_0778_;
	assign _1020_ = _1019_ | _1018_;
	assign _1021_ = _0504_ & ~_0782_;
	assign _1022_ = _0538_ & ~_0785_;
	assign _1023_ = _1022_ | _1021_;
	assign _1024_ = _1023_ | _1020_;
	assign _1025_ = _0571_ & ~_0791_;
	assign _1026_ = _0404_ & ~_0794_;
	assign _1027_ = _1026_ | _1025_;
	assign _1029_ = _0439_ & ~_0799_;
	assign _1030_ = _0747_ & ~_0803_;
	assign _1031_ = _1030_ | _1029_;
	assign _1032_ = _1031_ | _1027_;
	assign _1033_ = _1032_ | _1024_;
	assign _1034_ = _1016_ & ~_1033_;
	assign _1035_ = _0335_ & ~_0809_;
	assign _1036_ = _0602_ & ~_0812_;
	assign _1037_ = _0630_ & ~_0815_;
	assign _1038_ = _1037_ | _1036_;
	assign _1039_ = _1038_ | _1035_;
	assign _1040_ = _1034_ & ~_1039_;
	assign _1041_ = ~(_1040_ | _0842_);
	assign _1042_ = _0760_ | _0708_;
	assign _1043_ = _0747_ & ~_0757_;
	assign _1044_ = _1042_ & ~_1043_;
	assign _1045_ = _0630_ & ~_0776_;
	assign _1046_ = _0659_ & ~_0778_;
	assign _1047_ = _1046_ | _1045_;
	assign _1048_ = _0471_ & ~_0782_;
	assign _1050_ = _0504_ & ~_0785_;
	assign _1051_ = _1050_ | _1048_;
	assign _1052_ = _1051_ | _1047_;
	assign _1053_ = _0538_ & ~_0791_;
	assign _1054_ = _0571_ & ~_0794_;
	assign _1055_ = _1054_ | _1053_;
	assign _1056_ = _0404_ & ~_0799_;
	assign _1057_ = _0439_ & ~_0803_;
	assign _1058_ = _1057_ | _1056_;
	assign _1059_ = _1058_ | _1055_;
	assign _1060_ = _1059_ | _1052_;
	assign _1061_ = _1044_ & ~_1060_;
	assign _1062_ = _0307_ & ~_0809_;
	assign _1063_ = _0335_ & ~_0812_;
	assign _1064_ = _0602_ & ~_0815_;
	assign _1065_ = _1064_ | _1063_;
	assign _1066_ = _1065_ | _1062_;
	assign _1067_ = _1061_ & ~_1066_;
	assign _1068_ = ~(_1067_ | _0842_);
	assign _1069_ = _1068_ | _1041_;
	assign _1071_ = _0799_ | _0708_;
	assign _1072_ = _0439_ & ~_0791_;
	assign _1073_ = _0747_ & ~_0794_;
	assign _1074_ = _1073_ | _1072_;
	assign _1075_ = _1071_ & ~_1074_;
	assign _1076_ = _0504_ & ~_0776_;
	assign _1077_ = _0538_ & ~_0778_;
	assign _1078_ = _1077_ | _1076_;
	assign _1079_ = _0571_ & ~_0782_;
	assign _1080_ = _0404_ & ~_0785_;
	assign _1082_ = _1080_ | _1079_;
	assign _1083_ = _1082_ | _1078_;
	assign _1084_ = _1075_ & ~_1083_;
	assign _1085_ = _0630_ & ~_0809_;
	assign _1086_ = _0659_ & ~_0812_;
	assign _1087_ = _0471_ & ~_0815_;
	assign _1088_ = _1087_ | _1086_;
	assign _1089_ = _1088_ | _1085_;
	assign _1090_ = _1084_ & ~_1089_;
	assign _1091_ = _1090_ | _0842_;
	assign _1093_ = _0803_ | _0708_;
	assign _1094_ = _0747_ & ~_0799_;
	assign _1095_ = _1093_ & ~_1094_;
	assign _1096_ = _0404_ & ~_0791_;
	assign _1097_ = _0439_ & ~_0794_;
	assign _1098_ = _1097_ | _1096_;
	assign _1099_ = _1095_ & ~_1098_;
	assign _1100_ = _0471_ & ~_0776_;
	assign _1101_ = _0504_ & ~_0778_;
	assign _1102_ = _1101_ | _1100_;
	assign _1103_ = _0538_ & ~_0782_;
	assign _1104_ = _0571_ & ~_0785_;
	assign _1105_ = _1104_ | _1103_;
	assign _1106_ = _1105_ | _1102_;
	assign _1107_ = _1099_ & ~_1106_;
	assign _1108_ = _0602_ & ~_0809_;
	assign _1109_ = _0630_ & ~_0812_;
	assign _1110_ = _0659_ & ~_0815_;
	assign _1111_ = _1110_ | _1109_;
	assign _1112_ = _1111_ | _1108_;
	assign _1114_ = _1107_ & ~_1112_;
	assign _1115_ = ~(_1114_ | _0842_);
	assign _1116_ = _1115_ | ~_1091_;
	assign _1117_ = _1116_ | _1069_;
	assign _1118_ = _1117_ | _1015_;
	assign _1119_ = _1118_ | _0882_;
	assign _1120_ = ~(_1119_ | _0359_);
	assign _1121_ = _1120_ | _0340_;
	assign _1122_ = _1488_ | \mchip.value_B [14];
	assign _1123_ = _2236_ | _1499_;
	assign _1124_ = _1123_ | _1122_;
	assign _1125_ = _2225_ & ~_1124_;
	assign _1126_ = _1609_ | \mchip.value_A [14];
	assign _1127_ = _1620_ | ~_2300_;
	assign _1128_ = _1127_ | _1126_;
	assign _1129_ = _2376_ & ~_1128_;
	assign _1130_ = _1129_ | _1125_;
	assign _1131_ = _1130_ | _1121_;
	assign _1132_ = _2452_ & ~_1131_;
	assign _1133_ = ~_0335_;
	assign _1134_ = _0350_ ^ _0312_;
	assign _1135_ = ~(_0349_ ^ _0348_);
	assign _1136_ = (_0358_ ? _1134_ : _1135_);
	assign _1137_ = _0822_ & ~_0834_;
	assign _1138_ = ~(_1137_ | _0842_);
	assign _1139_ = _1138_ & ~_0094_;
	assign _1140_ = _0836_ | _0833_;
	assign _1141_ = _0829_ | _0821_;
	assign _1142_ = _1141_ | _1140_;
	assign _1143_ = _0840_ & ~_1142_;
	assign _1145_ = ~(_1143_ | _0842_);
	assign _1146_ = _1145_ & ~_0097_;
	assign _1147_ = _0750_ & ~_0828_;
	assign _1148_ = ~(_0769_ & _0760_);
	assign _1149_ = _1147_ & ~_1148_;
	assign _1150_ = ~(_0785_ & _0778_);
	assign _1151_ = ~(_0803_ & _0794_);
	assign _1152_ = _1151_ | _1150_;
	assign _1153_ = _1149_ & ~_1152_;
	assign _1154_ = ~(_0815_ & _0809_);
	assign _1156_ = _1153_ & ~_1154_;
	assign _1157_ = ~(_1156_ | _0842_);
	assign _1158_ = _1157_ | ~_0087_;
	assign _1159_ = ~(_1145_ ^ _0097_);
	assign _1160_ = _1159_ & _1158_;
	assign _1161_ = _1160_ | _1146_;
	assign _1162_ = ~(_1138_ ^ _0094_);
	assign _1163_ = _1162_ & _1161_;
	assign _1164_ = ~(_1163_ | _1139_);
	assign _1165_ = ~_0092_;
	assign _1166_ = _0822_ & ~_0837_;
	assign _1167_ = ~(_1166_ | _0842_);
	assign _1168_ = _1167_ ^ _1165_;
	assign _1169_ = _1168_ ^ _1164_;
	assign _1170_ = _1162_ ^ _1161_;
	assign _1171_ = _1170_ | ~_1169_;
	assign _1172_ = _1157_ ^ _0087_;
	assign _1173_ = _1159_ ^ _1158_;
	assign _1174_ = _1173_ | _1172_;
	assign _1175_ = _1174_ | _1171_;
	assign _1176_ = _1167_ & _1165_;
	assign _1177_ = _1168_ & _1139_;
	assign _1178_ = _1177_ | _1176_;
	assign _1179_ = ~(_1168_ & _1162_);
	assign _1180_ = _1161_ & ~_1179_;
	assign _1181_ = _1180_ | _1178_;
	assign _1182_ = _0830_ & ~_0842_;
	assign _1183_ = ~(_1182_ ^ _0107_);
	assign _1184_ = _1183_ ^ _1181_;
	assign _1185_ = _1184_ | _1175_;
	assign _1187_ = _1185_ | _1091_;
	assign _1188_ = ~_1115_;
	assign _1189_ = _1173_ | ~_1172_;
	assign _1190_ = _1189_ | _1171_;
	assign _1191_ = ~(_1190_ | _1184_);
	assign _1192_ = _1191_ & ~_1188_;
	assign _1193_ = _1187_ & ~_1192_;
	assign _1194_ = _1172_ | ~_1173_;
	assign _1195_ = _1194_ | _1171_;
	assign _1196_ = _1195_ | _1184_;
	assign _1198_ = _1041_ & ~_1196_;
	assign _1199_ = ~(_1173_ & _1172_);
	assign _1200_ = _1199_ | _1171_;
	assign _1201_ = _1200_ | _1184_;
	assign _1202_ = _1068_ & ~_1201_;
	assign _1203_ = _1202_ | _1198_;
	assign _1204_ = ~(_1170_ & _1169_);
	assign _1205_ = _1204_ | _1174_;
	assign _1206_ = _1205_ | _1184_;
	assign _1207_ = _0981_ & ~_1206_;
	assign _1208_ = _1204_ | _1189_;
	assign _1209_ = _1208_ | _1184_;
	assign _1210_ = _1013_ & ~_1209_;
	assign _1211_ = _1210_ | _1207_;
	assign _1212_ = _1211_ | _1203_;
	assign _1213_ = _1204_ | _1194_;
	assign _1214_ = _1213_ | _1184_;
	assign _1215_ = _0914_ & ~_1214_;
	assign _1216_ = _1204_ | _1199_;
	assign _1217_ = _1216_ | _1184_;
	assign _1219_ = _0950_ & ~_1217_;
	assign _1220_ = _1219_ | _1215_;
	assign _1221_ = _1170_ | _1169_;
	assign _1222_ = _1221_ | _1174_;
	assign _1223_ = _1222_ | _1184_;
	assign _1224_ = _0843_ & ~_1223_;
	assign _1225_ = _1221_ | _1189_;
	assign _1226_ = ~(_1225_ | _1184_);
	assign _1227_ = _1226_ & ~_0881_;
	assign _1228_ = _1227_ | _1224_;
	assign _1230_ = _1228_ | _1220_;
	assign _1231_ = _1230_ | _1212_;
	assign _1232_ = _1193_ & ~_1231_;
	assign _1233_ = _1223_ & ~_1226_;
	assign _1234_ = ~(_1217_ & _1214_);
	assign _1235_ = _1233_ & ~_1234_;
	assign _1236_ = ~(_1201_ & _1196_);
	assign _1237_ = ~(_1209_ & _1206_);
	assign _1238_ = _1237_ | _1236_;
	assign _1239_ = _1235_ & ~_1238_;
	assign _1241_ = _1191_ | ~_1185_;
	assign _1242_ = _1239_ & ~_1241_;
	assign _1243_ = _1242_ | _1232_;
	assign _1244_ = _1183_ & ~_0105_;
	assign _1245_ = _1172_ | ~_1159_;
	assign _1246_ = _1245_ | _1179_;
	assign _1247_ = _1244_ & ~_1246_;
	assign _1248_ = _0107_ | ~_1182_;
	assign _1249_ = _1248_ | _0105_;
	assign _1250_ = _1244_ & _1181_;
	assign _1251_ = _1249_ & ~_1250_;
	assign _1252_ = _1251_ | _1247_;
	assign _1253_ = (_1252_ ? _1091_ : _1243_);
	assign _1254_ = (_0359_ ? _1136_ : _1253_);
	assign _1255_ = (_2137_ ? _1254_ : _1133_);
	assign _1256_ = _1132_ & ~_1255_;
	assign _1257_ = ~(\mchip.value_A [15] ^ \mchip.value_B [15]);
	assign _1258_ = ~(\mchip.value_B [14] | \mchip.value_A [14]);
	assign _1259_ = ~(\mchip.value_B [13] ^ \mchip.value_A [13]);
	assign _1260_ = \mchip.value_B [12] ^ \mchip.value_A [12];
	assign _1261_ = _1259_ & ~_1260_;
	assign _1262_ = ~(\mchip.value_B [10] ^ \mchip.value_A [10]);
	assign _1263_ = ~(\mchip.value_B [11] ^ \mchip.value_A [11]);
	assign _1264_ = _1263_ & _1262_;
	assign _1265_ = ~(_1264_ & _1261_);
	assign _1266_ = \mchip.value_B [14] & \mchip.value_A [14];
	assign _1267_ = ~(_1266_ | _1258_);
	assign _1268_ = _1267_ | _1265_;
	assign _1269_ = \mchip.value_B [9] | ~\mchip.value_A [9];
	assign _1270_ = \mchip.value_B [8] | ~\mchip.value_A [8];
	assign _1272_ = ~(\mchip.value_A [9] | \mchip.value_B [9]);
	assign _1273_ = _1272_ | _2678_;
	assign _1274_ = _1273_ & ~_1270_;
	assign _1275_ = _1269_ & ~_1274_;
	assign _1276_ = \mchip.value_A [8] ^ \mchip.value_B [8];
	assign _1277_ = _1273_ & ~_1276_;
	assign _1278_ = \mchip.value_B [7] | ~\mchip.value_A [7];
	assign _1279_ = ~(\mchip.value_A [7] ^ \mchip.value_B [7]);
	assign _1280_ = \mchip.value_B [6] | ~\mchip.value_A [6];
	assign _1281_ = _1279_ & ~_1280_;
	assign _1282_ = _1278_ & ~_1281_;
	assign _1283_ = \mchip.value_A [6] ^ \mchip.value_B [6];
	assign _1284_ = _1279_ & ~_1283_;
	assign _1285_ = \mchip.value_B [5] | ~\mchip.value_A [5];
	assign _1286_ = \mchip.value_A [4] & ~\mchip.value_B [4];
	assign _1287_ = \mchip.value_B [5] ^ \mchip.value_A [5];
	assign _1288_ = _1286_ & ~_1287_;
	assign _1289_ = _1285_ & ~_1288_;
	assign _1290_ = _1284_ & ~_1289_;
	assign _1291_ = _1282_ & ~_1290_;
	assign _1292_ = \mchip.value_A [4] ^ \mchip.value_B [4];
	assign _1293_ = _1292_ | _1287_;
	assign _1294_ = _1284_ & ~_1293_;
	assign _1295_ = \mchip.value_B [3] | ~\mchip.value_A [3];
	assign _1296_ = ~(\mchip.value_A [3] ^ \mchip.value_B [3]);
	assign _1297_ = \mchip.value_B [2] | ~\mchip.value_A [2];
	assign _1298_ = _1296_ & ~_1297_;
	assign _1299_ = _1295_ & ~_1298_;
	assign _1300_ = \mchip.value_B [2] ^ \mchip.value_A [2];
	assign _1301_ = _1296_ & ~_1300_;
	assign _1303_ = \mchip.value_B [1] | ~\mchip.value_A [1];
	assign _1304_ = ~(\mchip.value_B [1] ^ \mchip.value_A [1]);
	assign _1305_ = \mchip.value_B [0] & ~\mchip.value_A [0];
	assign _1306_ = _1304_ & ~_1305_;
	assign _1307_ = _1303_ & ~_1306_;
	assign _1308_ = _1301_ & ~_1307_;
	assign _1309_ = _1299_ & ~_1308_;
	assign _1310_ = _1294_ & ~_1309_;
	assign _1311_ = _1291_ & ~_1310_;
	assign _1312_ = _1277_ & ~_1311_;
	assign _1313_ = _1275_ & ~_1312_;
	assign _1314_ = (_1313_ ? \mchip.value_B [11] : \mchip.value_A [11]);
	assign _1315_ = (_1268_ ? \mchip.value_A [11] : _1314_);
	assign _1316_ = \mchip.value_B [14] | ~\mchip.value_A [14];
	assign _1317_ = \mchip.value_B [13] | ~\mchip.value_A [13];
	assign _1318_ = \mchip.value_B [12] | ~\mchip.value_A [12];
	assign _1319_ = _1259_ & ~_1318_;
	assign _1320_ = _1317_ & ~_1319_;
	assign _1321_ = \mchip.value_B [11] | ~\mchip.value_A [11];
	assign _1322_ = \mchip.value_B [10] & ~\mchip.value_A [10];
	assign _1324_ = _1263_ & ~_1322_;
	assign _1325_ = _1321_ & ~_1324_;
	assign _1326_ = _1261_ & ~_1325_;
	assign _1327_ = _1326_ | ~_1320_;
	assign _1328_ = _1327_ & ~_1267_;
	assign _1329_ = _1316_ & ~_1328_;
	assign _1330_ = (_1329_ ? \mchip.value_B [11] : _1315_);
	assign _1331_ = (_1313_ ? \mchip.value_B [10] : \mchip.value_A [10]);
	assign _1332_ = (_1268_ ? \mchip.value_A [10] : _1331_);
	assign _1333_ = (_1329_ ? \mchip.value_B [10] : _1332_);
	assign _1335_ = _1333_ | _1330_;
	assign _1336_ = (_1313_ ? \mchip.value_B [13] : \mchip.value_A [13]);
	assign _1337_ = (_1268_ ? \mchip.value_A [13] : _1336_);
	assign _1338_ = (_1329_ ? \mchip.value_B [13] : _1337_);
	assign _1339_ = (_1313_ ? \mchip.value_B [12] : \mchip.value_A [12]);
	assign _1340_ = (_1268_ ? \mchip.value_A [12] : _1339_);
	assign _1341_ = (_1329_ ? \mchip.value_B [12] : _1340_);
	assign _1342_ = _1341_ | _1338_;
	assign _1343_ = _1342_ | _1335_;
	assign _1344_ = _1258_ & ~_1343_;
	assign _1345_ = ~(_1344_ & _1333_);
	assign _1346_ = _1330_ & ~_1345_;
	assign _1347_ = ~(_1341_ & _1338_);
	assign _1348_ = _1346_ & ~_1347_;
	assign _1349_ = _1348_ ^ _1258_;
	assign _1350_ = ~_1341_;
	assign _1351_ = _1346_ & ~_1350_;
	assign _1352_ = ~(_1351_ ^ _1338_);
	assign _1353_ = _1352_ | _1349_;
	assign _1354_ = _1346_ ^ _1341_;
	assign _1355_ = ~(_1345_ ^ _1330_);
	assign _1356_ = ~(_1355_ & _1354_);
	assign _1357_ = _1356_ | _1353_;
	assign _1358_ = ~(_1344_ ^ _1333_);
	assign _1359_ = _1358_ & ~_1357_;
	assign _1360_ = (_1313_ ? \mchip.value_A [13] : \mchip.value_B [13]);
	assign _1361_ = (_1268_ ? \mchip.value_B [13] : _1360_);
	assign _1362_ = (_1329_ ? \mchip.value_A [13] : _1361_);
	assign _1363_ = (_1313_ ? \mchip.value_A [12] : \mchip.value_B [12]);
	assign _1364_ = (_1268_ ? \mchip.value_B [12] : _1363_);
	assign _1365_ = (_1329_ ? \mchip.value_A [12] : _1364_);
	assign _1366_ = _1365_ | _1362_;
	assign _1367_ = (_1313_ ? \mchip.value_A [10] : \mchip.value_B [10]);
	assign _1368_ = (_1268_ ? \mchip.value_B [10] : _1367_);
	assign _1369_ = (_1329_ ? \mchip.value_A [10] : _1368_);
	assign _1370_ = (_1313_ ? \mchip.value_A [11] : \mchip.value_B [11]);
	assign _1371_ = (_1268_ ? \mchip.value_B [11] : _1370_);
	assign _1372_ = (_1329_ ? \mchip.value_A [11] : _1371_);
	assign _1373_ = _1372_ | _1369_;
	assign _1374_ = _1373_ | _1366_;
	assign _1375_ = ~(_1374_ | _1266_);
	assign _1376_ = ~_1365_;
	assign _1377_ = ~_1372_;
	assign _1378_ = _1374_ | _1266_;
	assign _1379_ = _1369_ & ~_1378_;
	assign _1380_ = _1379_ & ~_1377_;
	assign _1381_ = _1380_ & ~_1376_;
	assign _1382_ = ~(_1381_ ^ _1362_);
	assign _1383_ = _1382_ & ~_1352_;
	assign _1384_ = _1380_ ^ _1376_;
	assign _1385_ = _1384_ & _1354_;
	assign _1386_ = _1382_ ^ _1352_;
	assign _1387_ = _1385_ & ~_1386_;
	assign _1388_ = _1387_ | _1383_;
	assign _1389_ = _1379_ ^ _1377_;
	assign _1390_ = ~(_1389_ & _1355_);
	assign _1391_ = _1389_ ^ _1355_;
	assign _1392_ = _1378_ ^ _1369_;
	assign _1393_ = _1358_ & ~_1392_;
	assign _1394_ = _1391_ & ~_1393_;
	assign _1395_ = _1390_ & ~_1394_;
	assign _1396_ = _1384_ ^ _1354_;
	assign _1397_ = _1396_ & ~_1386_;
	assign _1398_ = _1397_ & ~_1395_;
	assign _1399_ = _1398_ | _1388_;
	assign _1400_ = ~(_1365_ & _1362_);
	assign _1401_ = _1380_ & ~_1400_;
	assign _1402_ = _1401_ ^ _1266_;
	assign _1403_ = _1402_ ^ _1349_;
	assign _1404_ = _1403_ ^ _1399_;
	assign _1405_ = _1396_ & ~_1395_;
	assign _1406_ = _1405_ | _1385_;
	assign _1407_ = ~(_1382_ ^ _1352_);
	assign _1408_ = _1407_ ^ _1406_;
	assign _1409_ = ~(_1395_ ^ _1396_);
	assign _1410_ = _1409_ | _1408_;
	assign _1411_ = ~(_1393_ ^ _1391_);
	assign _1412_ = ~(_1392_ ^ _1358_);
	assign _1413_ = ~_1412_;
	assign _1414_ = _1413_ | _1411_;
	assign _1415_ = _1414_ | _1410_;
	assign _1416_ = ~(_1415_ | _1404_);
	assign _1417_ = _1416_ & ~_1375_;
	assign _1418_ = _1412_ | _1411_;
	assign _1419_ = ~(_1418_ | _1410_);
	assign _1420_ = _1419_ & ~_1404_;
	assign _1421_ = _1420_ & ~_1375_;
	assign _1422_ = ~\mchip.value_A [9];
	assign _1423_ = ~\mchip.value_B [9];
	assign _1424_ = (_1268_ ? _1423_ : _2997_);
	assign _1425_ = (_1329_ ? _1422_ : _1424_);
	assign _1426_ = _1416_ & ~_1425_;
	assign _1427_ = ~(_1426_ | _1421_);
	assign _1428_ = ~_1409_;
	assign _1429_ = _1428_ | _1408_;
	assign _1430_ = ~(_1413_ & _1411_);
	assign _1431_ = _1430_ | _1429_;
	assign _1432_ = ~(_1431_ | _1404_);
	assign _1433_ = _1386_ ^ _1406_;
	assign _1434_ = _1433_ | _1409_;
	assign _1435_ = _1434_ | _1414_;
	assign _1436_ = ~(_1435_ | _1404_);
	assign _1437_ = _1436_ | _1432_;
	assign _1438_ = _1434_ | _1418_;
	assign _1439_ = ~(_1438_ | _1404_);
	assign _1440_ = ~(_1412_ & _1411_);
	assign _1441_ = _1440_ | _1434_;
	assign _1442_ = ~(_1441_ | _1404_);
	assign _1443_ = _1442_ | _1439_;
	assign _1444_ = ~(_1443_ | _1437_);
	assign _1445_ = _1430_ | _1410_;
	assign _1446_ = ~(_1445_ | _1404_);
	assign _1447_ = _1429_ | _1414_;
	assign _1448_ = ~(_1447_ | _1404_);
	assign _1449_ = _1448_ | _1446_;
	assign _1450_ = _1429_ | _1418_;
	assign _1451_ = ~(_1450_ | _1404_);
	assign _1452_ = _1440_ | _1429_;
	assign _1453_ = ~(_1452_ | _1404_);
	assign _1454_ = _1453_ | _1451_;
	assign _1456_ = _1454_ | _1449_;
	assign _1457_ = _1444_ & ~_1456_;
	assign _1458_ = _1440_ | _1410_;
	assign _1459_ = ~(_1458_ | _1404_);
	assign _1460_ = _1459_ | _1420_;
	assign _1461_ = _1460_ | _1416_;
	assign _1462_ = _1457_ & ~_1461_;
	assign _1463_ = ~(_1462_ | _1427_);
	assign _1464_ = _1375_ | ~_1459_;
	assign _1465_ = _1420_ & ~_1425_;
	assign _1467_ = _1464_ & ~_1465_;
	assign _1468_ = ~\mchip.value_A [8];
	assign _1469_ = ~\mchip.value_B [8];
	assign _1470_ = (_1313_ ? _1468_ : _1469_);
	assign _1471_ = (_1268_ ? _1469_ : _1470_);
	assign _1472_ = (_1329_ ? _1468_ : _1471_);
	assign _1473_ = _1416_ & ~_1472_;
	assign _1474_ = _1467_ & ~_1473_;
	assign _1475_ = ~(_1474_ | _1462_);
	assign _1476_ = _1475_ | _1463_;
	assign _1478_ = _1375_ | ~_1439_;
	assign _1479_ = _1432_ & ~_1472_;
	assign _1480_ = ~_1425_;
	assign _1481_ = _1436_ & _1480_;
	assign _1482_ = _1481_ | _1479_;
	assign _1483_ = _1478_ & ~_1482_;
	assign _1484_ = ~\mchip.value_A [4];
	assign _1485_ = ~\mchip.value_B [4];
	assign _1486_ = (_1313_ ? _1484_ : _1485_);
	assign _1487_ = (_1268_ ? _1485_ : _1486_);
	assign _1489_ = (_1329_ ? _1484_ : _1487_);
	assign _1490_ = _1446_ & ~_1489_;
	assign _1491_ = ~\mchip.value_A [5];
	assign _1492_ = ~\mchip.value_B [5];
	assign _1493_ = (_1313_ ? _1491_ : _1492_);
	assign _1494_ = (_1268_ ? _1492_ : _1493_);
	assign _1495_ = (_1329_ ? _1491_ : _1494_);
	assign _1496_ = _1448_ & ~_1495_;
	assign _1497_ = _1496_ | _1490_;
	assign _1498_ = ~\mchip.value_A [6];
	assign _1500_ = ~\mchip.value_B [6];
	assign _1501_ = (_1313_ ? _1498_ : _1500_);
	assign _1502_ = (_1268_ ? _1500_ : _1501_);
	assign _1503_ = (_1329_ ? _1498_ : _1502_);
	assign _1504_ = _1451_ & ~_1503_;
	assign _1505_ = ~\mchip.value_A [7];
	assign _1506_ = ~\mchip.value_B [7];
	assign _1507_ = (_1313_ ? _1505_ : _1506_);
	assign _1508_ = (_1268_ ? _1506_ : _1507_);
	assign _1509_ = (_1329_ ? _1505_ : _1508_);
	assign _1511_ = _1453_ & ~_1509_;
	assign _1512_ = _1511_ | _1504_;
	assign _1513_ = _1512_ | _1497_;
	assign _1514_ = _1483_ & ~_1513_;
	assign _1515_ = ~\mchip.value_A [1];
	assign _1516_ = ~\mchip.value_B [1];
	assign _1517_ = (_1313_ ? _1515_ : _1516_);
	assign _1518_ = (_1268_ ? _1516_ : _1517_);
	assign _1519_ = (_1329_ ? _1515_ : _1518_);
	assign _1520_ = _1416_ & ~_1519_;
	assign _1522_ = ~\mchip.value_A [2];
	assign _1523_ = ~\mchip.value_B [2];
	assign _1524_ = (_1313_ ? _1522_ : _1523_);
	assign _1525_ = (_1268_ ? _1523_ : _1524_);
	assign _1526_ = (_1329_ ? _1522_ : _1525_);
	assign _1527_ = _1420_ & ~_1526_;
	assign _1528_ = ~\mchip.value_A [3];
	assign _1529_ = ~\mchip.value_B [3];
	assign _1530_ = (_1313_ ? _1528_ : _1529_);
	assign _1531_ = (_1268_ ? _1529_ : _1530_);
	assign _1533_ = (_1329_ ? _1528_ : _1531_);
	assign _1534_ = _1459_ & ~_1533_;
	assign _1535_ = _1534_ | _1527_;
	assign _1536_ = _1535_ | _1520_;
	assign _1537_ = _1514_ & ~_1536_;
	assign _1538_ = _1537_ | _1462_;
	assign _1539_ = ~\mchip.value_A [0];
	assign _1540_ = ~\mchip.value_B [0];
	assign _1541_ = (_1313_ ? _1539_ : _1540_);
	assign _1542_ = (_1268_ ? _1540_ : _1541_);
	assign _1544_ = (_1329_ ? _1539_ : _1542_);
	assign _1545_ = _1544_ | ~_1416_;
	assign _1546_ = _1420_ & ~_1519_;
	assign _1547_ = _1459_ & ~_1526_;
	assign _1548_ = _1547_ | _1546_;
	assign _1549_ = _1545_ & ~_1548_;
	assign _1550_ = _1442_ & ~_1375_;
	assign _1551_ = _1439_ & _1480_;
	assign _1552_ = _1551_ | _1550_;
	assign _1553_ = _1432_ & ~_1509_;
	assign _1555_ = _1436_ & ~_1472_;
	assign _1556_ = _1555_ | _1553_;
	assign _1557_ = _1556_ | _1552_;
	assign _1558_ = _1446_ & ~_1533_;
	assign _1559_ = _1448_ & ~_1489_;
	assign _1560_ = _1559_ | _1558_;
	assign _1561_ = _1451_ & ~_1495_;
	assign _1562_ = _1453_ & ~_1503_;
	assign _1563_ = _1562_ | _1561_;
	assign _1564_ = _1563_ | _1560_;
	assign _1566_ = _1564_ | _1557_;
	assign _1567_ = _1549_ & ~_1566_;
	assign _1568_ = ~(_1567_ | _1462_);
	assign _1569_ = _1538_ & ~_1568_;
	assign _1570_ = _1375_ | ~_1436_;
	assign _1571_ = _1432_ & _1480_;
	assign _1572_ = _1570_ & ~_1571_;
	assign _1573_ = _1446_ & ~_1495_;
	assign _1574_ = _1448_ & ~_1503_;
	assign _1575_ = _1574_ | _1573_;
	assign _1577_ = _1451_ & ~_1509_;
	assign _1578_ = _1453_ & ~_1472_;
	assign _1579_ = _1578_ | _1577_;
	assign _1580_ = _1579_ | _1575_;
	assign _1581_ = _1572_ & ~_1580_;
	assign _1582_ = _1416_ & ~_1526_;
	assign _1583_ = _1420_ & ~_1533_;
	assign _1584_ = _1459_ & ~_1489_;
	assign _1585_ = _1584_ | _1583_;
	assign _1586_ = _1585_ | _1582_;
	assign _1588_ = _1581_ & ~_1586_;
	assign _1589_ = ~(_1588_ | _1462_);
	assign _1590_ = _1375_ | ~_1432_;
	assign _1591_ = _1446_ & ~_1503_;
	assign _1592_ = _1448_ & ~_1509_;
	assign _1593_ = _1592_ | _1591_;
	assign _1594_ = _1451_ & ~_1472_;
	assign _1595_ = _1453_ & _1480_;
	assign _1596_ = _1595_ | _1594_;
	assign _1597_ = _1596_ | _1593_;
	assign _1599_ = _1590_ & ~_1597_;
	assign _1600_ = _1416_ & ~_1533_;
	assign _1601_ = _1420_ & ~_1489_;
	assign _1602_ = _1459_ & ~_1495_;
	assign _1603_ = _1602_ | _1601_;
	assign _1604_ = _1603_ | _1600_;
	assign _1605_ = _1599_ & ~_1604_;
	assign _1606_ = ~(_1605_ | _1462_);
	assign _1607_ = _1606_ | _1589_;
	assign _1608_ = _1569_ & ~_1607_;
	assign _1610_ = _1375_ | ~_1448_;
	assign _1611_ = _1446_ & _1480_;
	assign _1612_ = _1610_ & ~_1611_;
	assign _1613_ = _1416_ & ~_1503_;
	assign _1614_ = _1420_ & ~_1509_;
	assign _1615_ = _1459_ & ~_1472_;
	assign _1616_ = _1615_ | _1614_;
	assign _1617_ = _1616_ | _1613_;
	assign _1618_ = _1612_ & ~_1617_;
	assign _1619_ = ~(_1618_ | _1462_);
	assign _1621_ = _1375_ | ~_1446_;
	assign _1622_ = _1416_ & ~_1509_;
	assign _1623_ = _1420_ & ~_1472_;
	assign _1624_ = _1459_ & _1480_;
	assign _1625_ = _1624_ | _1623_;
	assign _1626_ = _1625_ | _1622_;
	assign _1627_ = _1621_ & ~_1626_;
	assign _1628_ = ~(_1627_ | _1462_);
	assign _1629_ = _1628_ | _1619_;
	assign _1630_ = _1375_ | ~_1453_;
	assign _1632_ = _1451_ & _1480_;
	assign _1633_ = _1630_ & ~_1632_;
	assign _1634_ = _1446_ & ~_1509_;
	assign _1635_ = _1448_ & ~_1472_;
	assign _1636_ = _1635_ | _1634_;
	assign _1637_ = _1633_ & ~_1636_;
	assign _1638_ = _1416_ & ~_1489_;
	assign _1639_ = _1420_ & ~_1495_;
	assign _1640_ = _1459_ & ~_1503_;
	assign _1641_ = _1640_ | _1639_;
	assign _1643_ = _1641_ | _1638_;
	assign _1644_ = _1637_ & ~_1643_;
	assign _1645_ = ~(_1644_ | _1462_);
	assign _1646_ = _1375_ | ~_1451_;
	assign _1647_ = _1446_ & ~_1472_;
	assign _1648_ = _1448_ & _1480_;
	assign _1649_ = _1648_ | _1647_;
	assign _1650_ = _1646_ & ~_1649_;
	assign _1651_ = _1416_ & ~_1495_;
	assign _1652_ = _1420_ & ~_1503_;
	assign _1654_ = _1459_ & ~_1509_;
	assign _1655_ = _1654_ | _1652_;
	assign _1656_ = _1655_ | _1651_;
	assign _1657_ = _1650_ & ~_1656_;
	assign _1658_ = ~(_1657_ | _1462_);
	assign _1659_ = _1658_ | _1645_;
	assign _1660_ = _1659_ | _1629_;
	assign _1661_ = _1660_ | ~_1608_;
	assign _1662_ = _1661_ | _1476_;
	assign _1663_ = _1417_ ^ _1662_;
	assign _1665_ = (_1257_ ? _1417_ : _1663_);
	assign _1666_ = _1665_ & ~_1344_;
	assign _1667_ = _1665_ ^ _1344_;
	assign _1668_ = ~_1667_;
	assign _1669_ = (_1268_ ? _1422_ : _1272_);
	assign _1670_ = (_1329_ ? _1423_ : _1669_);
	assign _1671_ = ~_1670_;
	assign _1672_ = _1661_ | _1475_;
	assign _1673_ = _1672_ ^ _1463_;
	assign _1674_ = (_1257_ ? _1463_ : _1673_);
	assign _1676_ = ~(_1674_ & _1671_);
	assign _1677_ = _1674_ ^ _1671_;
	assign _1678_ = (_1313_ ? _1469_ : _1468_);
	assign _1679_ = (_1268_ ? _1468_ : _1678_);
	assign _1680_ = (_1329_ ? _1469_ : _1679_);
	assign _1681_ = _1661_ ^ _1475_;
	assign _1682_ = (_1257_ ? _1475_ : _1681_);
	assign _1683_ = _1680_ | ~_1682_;
	assign _1684_ = _1677_ & ~_1683_;
	assign _1685_ = _1676_ & ~_1684_;
	assign _1687_ = ~(_1682_ ^ _1680_);
	assign _1688_ = ~_1687_;
	assign _1689_ = _1677_ & ~_1688_;
	assign _1690_ = (_1313_ ? \mchip.value_B [7] : \mchip.value_A [7]);
	assign _1691_ = (_1268_ ? \mchip.value_A [7] : _1690_);
	assign _1692_ = (_1329_ ? \mchip.value_B [7] : _1691_);
	assign _1693_ = _1608_ & ~_1659_;
	assign _1694_ = _1693_ & ~_1619_;
	assign _1695_ = ~(_1694_ ^ _1628_);
	assign _1696_ = (_1257_ ? _1628_ : _1695_);
	assign _1698_ = ~(_1696_ & _1692_);
	assign _1699_ = _1696_ ^ _1692_;
	assign _1700_ = (_1313_ ? _1500_ : _1498_);
	assign _1701_ = (_1268_ ? _1498_ : _1700_);
	assign _1702_ = (_1329_ ? _1500_ : _1701_);
	assign _1703_ = ~(_1693_ ^ _1619_);
	assign _1704_ = (_1257_ ? _1619_ : _1703_);
	assign _1705_ = _1702_ | ~_1704_;
	assign _1706_ = _1699_ & ~_1705_;
	assign _1707_ = _1698_ & ~_1706_;
	assign _1709_ = _1704_ ^ _1702_;
	assign _1710_ = _1699_ & ~_1709_;
	assign _1711_ = (_1313_ ? _1492_ : _1491_);
	assign _1712_ = (_1268_ ? _1491_ : _1711_);
	assign _1713_ = (_1329_ ? _1492_ : _1712_);
	assign _1714_ = _1608_ & ~_1645_;
	assign _1715_ = ~(_1714_ ^ _1658_);
	assign _1716_ = (_1257_ ? _1658_ : _1715_);
	assign _1717_ = _1713_ | ~_1716_;
	assign _1718_ = ~(_1716_ ^ _1713_);
	assign _1720_ = (_1313_ ? _1485_ : _1484_);
	assign _1721_ = (_1268_ ? _1484_ : _1720_);
	assign _1722_ = (_1329_ ? _1485_ : _1721_);
	assign _1723_ = ~(_1645_ ^ _1608_);
	assign _1724_ = (_1257_ ? _1645_ : _1723_);
	assign _1725_ = _1722_ | ~_1724_;
	assign _1726_ = _1718_ & ~_1725_;
	assign _1727_ = _1717_ & ~_1726_;
	assign _1728_ = _1710_ & ~_1727_;
	assign _1729_ = _1707_ & ~_1728_;
	assign _1731_ = _1724_ ^ _1722_;
	assign _1732_ = _1718_ & ~_1731_;
	assign _1733_ = _1732_ & _1710_;
	assign _1734_ = (_1313_ ? _1529_ : _1528_);
	assign _1735_ = (_1268_ ? _1528_ : _1734_);
	assign _1736_ = (_1329_ ? _1529_ : _1735_);
	assign _1737_ = _1569_ & ~_1589_;
	assign _1738_ = ~(_1737_ ^ _1606_);
	assign _1739_ = (_1257_ ? _1606_ : _1738_);
	assign _1740_ = _1736_ | ~_1739_;
	assign _1742_ = ~(_1739_ ^ _1736_);
	assign _1743_ = (_1313_ ? _1523_ : _1522_);
	assign _1744_ = (_1268_ ? _1522_ : _1743_);
	assign _1745_ = (_1329_ ? _1523_ : _1744_);
	assign _1746_ = ~(_1589_ ^ _1569_);
	assign _1747_ = (_1257_ ? _1589_ : _1746_);
	assign _1748_ = _1745_ | ~_1747_;
	assign _1749_ = _1742_ & ~_1748_;
	assign _1750_ = _1740_ & ~_1749_;
	assign _1751_ = _1747_ ^ _1745_;
	assign _1753_ = _1742_ & ~_1751_;
	assign _1754_ = (_1313_ ? _1516_ : _1515_);
	assign _1755_ = (_1268_ ? _1515_ : _1754_);
	assign _1756_ = (_1329_ ? _1516_ : _1755_);
	assign _1757_ = ~(_1537_ | _1462_);
	assign _1758_ = ~(_1568_ ^ _1538_);
	assign _1759_ = (_1257_ ? _1757_ : _1758_);
	assign _1760_ = _1756_ | ~_1759_;
	assign _1761_ = (_1313_ ? _1540_ : _1539_);
	assign _1762_ = (_1268_ ? _1539_ : _1761_);
	assign _1764_ = (_1329_ ? _1540_ : _1762_);
	assign _1765_ = _1568_ & ~_1764_;
	assign _1766_ = _1759_ ^ _1756_;
	assign _1767_ = _1765_ & ~_1766_;
	assign _1768_ = _1760_ & ~_1767_;
	assign _1769_ = _1753_ & ~_1768_;
	assign _1770_ = _1750_ & ~_1769_;
	assign _1771_ = _1733_ & ~_1770_;
	assign _1772_ = _1729_ & ~_1771_;
	assign _1773_ = _1689_ & ~_1772_;
	assign _1775_ = _1685_ & ~_1773_;
	assign _1776_ = _1668_ & ~_1775_;
	assign _1777_ = ~(_1776_ | _1666_);
	assign _1778_ = _1777_ | ~_1359_;
	assign _1779_ = _1257_ & ~_1778_;
	assign _1780_ = ~(_1779_ | _2441_);
	assign _1781_ = _1764_ ^ _1568_;
	assign _1782_ = ~_1781_;
	assign _1783_ = ~_1709_;
	assign _1784_ = _1732_ & ~_1770_;
	assign _1786_ = _1727_ & ~_1784_;
	assign _1787_ = _1783_ & ~_1786_;
	assign _1788_ = _1705_ & ~_1787_;
	assign _1789_ = ~(_1788_ ^ _1699_);
	assign _1790_ = _1786_ ^ _1709_;
	assign _1791_ = _1790_ & ~_1789_;
	assign _1792_ = _1687_ & ~_1772_;
	assign _1793_ = _1683_ & ~_1792_;
	assign _1794_ = ~(_1793_ ^ _1677_);
	assign _1795_ = _1772_ ^ _1687_;
	assign _1797_ = ~_1795_;
	assign _1798_ = _1797_ | _1794_;
	assign _1799_ = _1791_ & ~_1798_;
	assign _1800_ = _1775_ ^ _1667_;
	assign _1801_ = _1799_ & ~_1800_;
	assign _1802_ = ~(_1770_ | _1731_);
	assign _1803_ = _1725_ & ~_1802_;
	assign _1804_ = ~(_1803_ ^ _1718_);
	assign _1805_ = _1804_ & ~_1790_;
	assign _1806_ = _1797_ | _1789_;
	assign _1808_ = _1805_ & ~_1806_;
	assign _1809_ = _1800_ | _1794_;
	assign _1810_ = _1808_ & ~_1809_;
	assign _1811_ = _1810_ | _1801_;
	assign _1812_ = _1790_ | _1789_;
	assign _1813_ = _1770_ ^ _1731_;
	assign _1814_ = _1813_ & ~_1804_;
	assign _1815_ = _1814_ & ~_1812_;
	assign _1816_ = _1800_ | _1798_;
	assign _1817_ = _1815_ & ~_1816_;
	assign _1819_ = ~(_1768_ | _1751_);
	assign _1820_ = _1748_ & ~_1819_;
	assign _1821_ = ~(_1820_ ^ _1742_);
	assign _1822_ = _1821_ & ~_1813_;
	assign _1823_ = _1804_ | _1790_;
	assign _1824_ = _1822_ & ~_1823_;
	assign _1825_ = _1809_ | _1806_;
	assign _1826_ = _1824_ & ~_1825_;
	assign _1827_ = _1826_ | _1817_;
	assign _1828_ = _1827_ | _1811_;
	assign _1830_ = _1768_ ^ _1751_;
	assign _1831_ = ~(_1766_ ^ _1765_);
	assign _1832_ = _1830_ | ~_1831_;
	assign _1833_ = _1821_ | _1813_;
	assign _1834_ = _1833_ | _1832_;
	assign _1835_ = _1823_ | _1806_;
	assign _1836_ = _1835_ | _1834_;
	assign _1837_ = ~(_1836_ | _1809_);
	assign _1838_ = ~_1800_;
	assign _1839_ = _1812_ | _1798_;
	assign _1841_ = _1813_ | _1804_;
	assign _1842_ = ~_1830_;
	assign _1843_ = _1842_ | _1821_;
	assign _1844_ = _1843_ | _1841_;
	assign _1845_ = _1844_ | _1839_;
	assign _1846_ = _1838_ & ~_1845_;
	assign _1847_ = _1846_ | _1837_;
	assign _1848_ = _1847_ | _1827_;
	assign _1849_ = _1795_ | _1794_;
	assign _1850_ = _1838_ & ~_1849_;
	assign _1852_ = _1789_ & ~_1797_;
	assign _1853_ = _1852_ & ~_1809_;
	assign _1854_ = _1853_ | _1850_;
	assign _1855_ = _1854_ | _1811_;
	assign _1856_ = _1855_ | _1848_;
	assign _1857_ = ~(_1856_ | _1809_);
	assign _1858_ = _1828_ & ~_1857_;
	assign _1859_ = _1857_ | _1847_;
	assign _1860_ = _1859_ | _1858_;
	assign _1861_ = _1800_ | ~_1794_;
	assign _1863_ = _1853_ | _1810_;
	assign _1864_ = _1837_ | _1826_;
	assign _1865_ = _1864_ | _1863_;
	assign _1866_ = _1861_ & ~_1865_;
	assign _1867_ = ~(_1866_ | _1857_);
	assign _1868_ = _1854_ | _1827_;
	assign _1869_ = ~(_1868_ | _1857_);
	assign _1870_ = _1867_ | ~_1869_;
	assign _1871_ = _1870_ | _1860_;
	assign _1872_ = _1871_ | ~_1782_;
	assign _1874_ = _1434_ | _1430_;
	assign _1875_ = _1874_ | _1404_;
	assign _1876_ = ~(_1875_ | _1375_);
	assign _1877_ = _1439_ & ~_1472_;
	assign _1878_ = _1442_ & _1480_;
	assign _1879_ = _1878_ | _1877_;
	assign _1880_ = ~(_1879_ | _1876_);
	assign _1881_ = _1451_ & ~_1489_;
	assign _1882_ = _1453_ & ~_1495_;
	assign _1883_ = _1882_ | _1881_;
	assign _1885_ = _1432_ & ~_1503_;
	assign _1886_ = _1436_ & ~_1509_;
	assign _1887_ = _1886_ | _1885_;
	assign _1888_ = _1887_ | _1883_;
	assign _1889_ = _1880_ & ~_1888_;
	assign _1890_ = _1420_ & ~_1544_;
	assign _1891_ = _1459_ & ~_1519_;
	assign _1892_ = _1891_ | _1890_;
	assign _1893_ = _1446_ & ~_1526_;
	assign _1894_ = _1448_ & ~_1533_;
	assign _1896_ = _1894_ | _1893_;
	assign _1897_ = _1896_ | _1892_;
	assign _1898_ = _1889_ & ~_1897_;
	assign _1899_ = _1447_ | ~_1404_;
	assign _1900_ = _1404_ & ~_1450_;
	assign _1901_ = _1899_ & ~_1900_;
	assign _1902_ = _1458_ | ~_1404_;
	assign _1903_ = _1445_ | ~_1404_;
	assign _1904_ = ~(_1903_ & _1902_);
	assign _1905_ = _1901_ & ~_1904_;
	assign _1907_ = _1433_ | _1428_;
	assign _1908_ = _1907_ | _1418_;
	assign _1909_ = _1908_ | _1404_;
	assign _1910_ = _1907_ | _1440_;
	assign _1911_ = _1910_ | _1404_;
	assign _1912_ = ~(_1911_ & _1909_);
	assign _1913_ = ~_1415_;
	assign _1914_ = ~(_1907_ | _1430_);
	assign _1915_ = (_1404_ ? _1913_ : _1914_);
	assign _1916_ = _1404_ & _1419_;
	assign _1918_ = _1916_ | _1915_;
	assign _1919_ = _1918_ | _1912_;
	assign _1920_ = _1905_ & ~_1919_;
	assign _1921_ = _1454_ | _1437_;
	assign _1922_ = _1907_ | _1414_;
	assign _1923_ = _1922_ | _1404_;
	assign _1924_ = ~(_1923_ & _1875_);
	assign _1925_ = _1924_ | _1443_;
	assign _1926_ = _1925_ | _1921_;
	assign _1927_ = _1920_ & ~_1926_;
	assign _1929_ = _1460_ | _1449_;
	assign _1930_ = _1927_ & ~_1929_;
	assign _1931_ = ~(_1930_ | _1898_);
	assign _1932_ = ~(_1869_ & _1867_);
	assign _1933_ = _1932_ | _1860_;
	assign _1934_ = _1931_ & ~_1933_;
	assign _1935_ = _1872_ & ~_1934_;
	assign _1936_ = _1923_ | _1375_;
	assign _1937_ = _1480_ & ~_1875_;
	assign _1938_ = _1936_ & ~_1937_;
	assign _1940_ = _1439_ & ~_1509_;
	assign _1941_ = _1442_ & ~_1472_;
	assign _1942_ = _1941_ | _1940_;
	assign _1943_ = _1938_ & ~_1942_;
	assign _1944_ = _1451_ & ~_1533_;
	assign _1945_ = _1453_ & ~_1489_;
	assign _1946_ = _1945_ | _1944_;
	assign _1947_ = _1432_ & ~_1495_;
	assign _1948_ = _1436_ & ~_1503_;
	assign _1949_ = _1948_ | _1947_;
	assign _1951_ = _1949_ | _1946_;
	assign _1952_ = _1943_ & ~_1951_;
	assign _1953_ = _1459_ & ~_1544_;
	assign _1954_ = _1446_ & ~_1519_;
	assign _1955_ = _1448_ & ~_1526_;
	assign _1956_ = _1955_ | _1954_;
	assign _1957_ = _1956_ | _1953_;
	assign _1958_ = _1952_ & ~_1957_;
	assign _1959_ = ~(_1958_ | _1930_);
	assign _1960_ = _1869_ | _1867_;
	assign _1962_ = _1960_ | _1860_;
	assign _1963_ = _1959_ & ~_1962_;
	assign _1964_ = _1909_ | _1375_;
	assign _1965_ = _1451_ & ~_1526_;
	assign _1966_ = _1453_ & ~_1533_;
	assign _1967_ = _1966_ | _1965_;
	assign _1968_ = _1432_ & ~_1489_;
	assign _1969_ = _1436_ & ~_1495_;
	assign _1970_ = _1969_ | _1968_;
	assign _1971_ = _1970_ | _1967_;
	assign _1973_ = _1439_ & ~_1503_;
	assign _1974_ = _1442_ & ~_1509_;
	assign _1975_ = _1974_ | _1973_;
	assign _1976_ = ~(_1875_ | _1472_);
	assign _1977_ = _1480_ & ~_1923_;
	assign _1978_ = _1977_ | _1976_;
	assign _1979_ = _1978_ | _1975_;
	assign _1980_ = _1979_ | _1971_;
	assign _1981_ = _1964_ & ~_1980_;
	assign _1982_ = _1446_ & ~_1544_;
	assign _1984_ = _1448_ & ~_1519_;
	assign _1985_ = _1984_ | _1982_;
	assign _1986_ = _1981_ & ~_1985_;
	assign _1987_ = ~(_1986_ | _1930_);
	assign _1988_ = _1869_ | ~_1867_;
	assign _1989_ = _1988_ | _1860_;
	assign _1990_ = _1987_ & ~_1989_;
	assign _1991_ = _1990_ | _1963_;
	assign _1992_ = _1911_ | _1375_;
	assign _1993_ = _1480_ & ~_1909_;
	assign _1995_ = _1992_ & ~_1993_;
	assign _1996_ = _1451_ & ~_1519_;
	assign _1997_ = _1453_ & ~_1526_;
	assign _1998_ = _1997_ | _1996_;
	assign _1999_ = _1432_ & ~_1533_;
	assign _2000_ = _1436_ & ~_1489_;
	assign _2001_ = _2000_ | _1999_;
	assign _2002_ = _2001_ | _1998_;
	assign _2003_ = _1439_ & ~_1495_;
	assign _2004_ = _1442_ & ~_1503_;
	assign _2006_ = _2004_ | _2003_;
	assign _2007_ = ~(_1875_ | _1509_);
	assign _2008_ = ~(_1923_ | _1472_);
	assign _2009_ = _2008_ | _2007_;
	assign _2010_ = _2009_ | _2006_;
	assign _2011_ = _2010_ | _2002_;
	assign _2012_ = _1995_ & ~_2011_;
	assign _2013_ = _1448_ & ~_1544_;
	assign _2014_ = _2012_ & ~_2013_;
	assign _2015_ = ~(_2014_ | _1930_);
	assign _2017_ = ~(_1857_ | _1847_);
	assign _2018_ = ~(_2017_ & _1858_);
	assign _2019_ = _2018_ | _1870_;
	assign _2020_ = _2015_ & ~_2019_;
	assign _2021_ = _2018_ | _1932_;
	assign _2022_ = ~(_1915_ & _1378_);
	assign _2023_ = ~(_1909_ | _1472_);
	assign _2024_ = _1480_ & ~_1911_;
	assign _2025_ = _2024_ | _2023_;
	assign _2026_ = _2022_ & ~_2025_;
	assign _2028_ = _1451_ & ~_1544_;
	assign _2029_ = _1453_ & ~_1519_;
	assign _2030_ = _2029_ | _2028_;
	assign _2031_ = _1432_ & ~_1526_;
	assign _2032_ = _1436_ & ~_1533_;
	assign _2033_ = _2032_ | _2031_;
	assign _2034_ = _2033_ | _2030_;
	assign _2035_ = _1439_ & ~_1489_;
	assign _2036_ = _1442_ & ~_1495_;
	assign _2037_ = _2036_ | _2035_;
	assign _2039_ = ~(_1875_ | _1503_);
	assign _2040_ = ~(_1923_ | _1509_);
	assign _2041_ = _2040_ | _2039_;
	assign _2042_ = _2041_ | _2037_;
	assign _2043_ = _2042_ | _2034_;
	assign _2044_ = _2026_ & ~_2043_;
	assign _2045_ = ~(_2044_ | _1930_);
	assign _2046_ = _2045_ & ~_2021_;
	assign _2047_ = _2046_ | _2020_;
	assign _2048_ = _2047_ | _1991_;
	assign _2050_ = _2018_ | _1960_;
	assign _2051_ = ~(_1916_ & _1378_);
	assign _2052_ = _1915_ & ~_1425_;
	assign _2053_ = _2051_ & ~_2052_;
	assign _2054_ = ~(_1909_ | _1509_);
	assign _2055_ = ~(_1911_ | _1472_);
	assign _2056_ = _2055_ | _2054_;
	assign _2057_ = _2053_ & ~_2056_;
	assign _2058_ = _1453_ & ~_1544_;
	assign _2059_ = _1432_ & ~_1519_;
	assign _2061_ = _1436_ & ~_1526_;
	assign _2062_ = _2061_ | _2059_;
	assign _2063_ = _2062_ | _2058_;
	assign _2064_ = _1439_ & ~_1533_;
	assign _2065_ = _1442_ & ~_1489_;
	assign _2066_ = _2065_ | _2064_;
	assign _2067_ = ~(_1875_ | _1495_);
	assign _2068_ = ~(_1923_ | _1503_);
	assign _2069_ = _2068_ | _2067_;
	assign _2070_ = _2069_ | _2066_;
	assign _2072_ = _2070_ | _2063_;
	assign _2073_ = _2057_ & ~_2072_;
	assign _2074_ = _2073_ | _1930_;
	assign _2075_ = ~(_2074_ | _2050_);
	assign _2076_ = _2018_ | _1988_;
	assign _2077_ = _1902_ | _1375_;
	assign _2078_ = ~(_1909_ | _1503_);
	assign _2079_ = ~(_1911_ | _1509_);
	assign _2080_ = _2079_ | _2078_;
	assign _2081_ = _1915_ & ~_1472_;
	assign _2083_ = _1916_ & ~_1425_;
	assign _2084_ = _2083_ | _2081_;
	assign _2085_ = _2084_ | _2080_;
	assign _2086_ = _2077_ & ~_2085_;
	assign _2087_ = _1432_ & ~_1544_;
	assign _2088_ = _1436_ & ~_1519_;
	assign _2089_ = _2088_ | _2087_;
	assign _2090_ = _1439_ & ~_1526_;
	assign _2091_ = _1442_ & ~_1533_;
	assign _2092_ = _2091_ | _2090_;
	assign _2094_ = ~(_1875_ | _1489_);
	assign _2095_ = ~(_1923_ | _1495_);
	assign _2096_ = _2095_ | _2094_;
	assign _2097_ = _2096_ | _2092_;
	assign _2098_ = _2097_ | _2089_;
	assign _2099_ = _2086_ & ~_2098_;
	assign _2100_ = _2099_ | _1930_;
	assign _2101_ = ~(_2100_ | _2076_);
	assign _2102_ = _2101_ | _2075_;
	assign _2103_ = _2017_ | _1858_;
	assign _2105_ = _2103_ | _1870_;
	assign _2106_ = _1903_ | _1375_;
	assign _2107_ = _1480_ & ~_1902_;
	assign _2108_ = _2106_ & ~_2107_;
	assign _2109_ = ~(_1909_ | _1495_);
	assign _2110_ = ~(_1911_ | _1503_);
	assign _2111_ = _2110_ | _2109_;
	assign _2112_ = _1915_ & ~_1509_;
	assign _2113_ = _1916_ & ~_1472_;
	assign _2114_ = _2113_ | _2112_;
	assign _2116_ = _2114_ | _2111_;
	assign _2117_ = _2108_ & ~_2116_;
	assign _2118_ = _1436_ & ~_1544_;
	assign _2119_ = _1439_ & ~_1519_;
	assign _2120_ = _1442_ & ~_1526_;
	assign _2121_ = _2120_ | _2119_;
	assign _2122_ = ~(_1875_ | _1533_);
	assign _2123_ = ~(_1923_ | _1489_);
	assign _2124_ = _2123_ | _2122_;
	assign _2125_ = _2124_ | _2121_;
	assign _2127_ = _2125_ | _2118_;
	assign _2128_ = _2117_ & ~_2127_;
	assign _2129_ = _2128_ | _1930_;
	assign _2130_ = ~(_2129_ | _2105_);
	assign _2131_ = _1899_ | _1375_;
	assign _2132_ = ~(_1902_ | _1472_);
	assign _2133_ = _1480_ & ~_1903_;
	assign _2134_ = _2133_ | _2132_;
	assign _2135_ = _2131_ & ~_2134_;
	assign _2136_ = ~(_1909_ | _1489_);
	assign _2138_ = ~(_1911_ | _1495_);
	assign _2139_ = _2138_ | _2136_;
	assign _2140_ = _1915_ & ~_1503_;
	assign _2141_ = _1916_ & ~_1509_;
	assign _2142_ = _2141_ | _2140_;
	assign _2143_ = _2142_ | _2139_;
	assign _2144_ = _2135_ & ~_2143_;
	assign _2145_ = _1439_ & ~_1544_;
	assign _2146_ = _1442_ & ~_1519_;
	assign _2147_ = _2146_ | _2145_;
	assign _2149_ = ~(_1875_ | _1526_);
	assign _2150_ = ~(_1923_ | _1533_);
	assign _2151_ = _2150_ | _2149_;
	assign _2152_ = _2151_ | _2147_;
	assign _2153_ = _2144_ & ~_2152_;
	assign _2154_ = ~(_2153_ | _1930_);
	assign _2155_ = _2103_ | _1932_;
	assign _2156_ = _2154_ & ~_2155_;
	assign _2157_ = _2156_ | _2130_;
	assign _2158_ = _2157_ | _2102_;
	assign _2160_ = _2158_ | _2048_;
	assign _2161_ = _1935_ & ~_2160_;
	assign _2162_ = _2155_ & _2105_;
	assign _2163_ = ~(_2076_ & _2050_);
	assign _2164_ = _2162_ & ~_2163_;
	assign _2165_ = ~(_1989_ & _1962_);
	assign _2166_ = ~(_2021_ & _2019_);
	assign _2167_ = _2166_ | _2165_;
	assign _2168_ = _2164_ & ~_2167_;
	assign _2169_ = ~(_1933_ & _1871_);
	assign _2171_ = _2168_ & ~_2169_;
	assign _2172_ = _1544_ | ~_1442_;
	assign _2173_ = ~(_1875_ | _1519_);
	assign _2174_ = ~(_1923_ | _1526_);
	assign _2175_ = _2174_ | _2173_;
	assign _2176_ = _2172_ & ~_2175_;
	assign _2177_ = ~(_1909_ | _1533_);
	assign _2178_ = ~(_1911_ | _1489_);
	assign _2179_ = _2178_ | _2177_;
	assign _2180_ = _1915_ & ~_1495_;
	assign _2182_ = _1916_ & ~_1503_;
	assign _2183_ = _2182_ | _2180_;
	assign _2184_ = _2183_ | _2179_;
	assign _2185_ = ~(_1902_ | _1509_);
	assign _2186_ = ~(_1903_ | _1472_);
	assign _2187_ = _2186_ | _2185_;
	assign _2188_ = _1480_ & ~_1899_;
	assign _2189_ = _1900_ & ~_1375_;
	assign _2190_ = _2189_ | _2188_;
	assign _2191_ = _2190_ | _2187_;
	assign _2193_ = _2191_ | _2184_;
	assign _2194_ = _2176_ & ~_2193_;
	assign _2195_ = _2194_ | _1930_;
	assign _2196_ = (_2171_ ? _2195_ : _2161_);
	assign _2197_ = ~(_1859_ & _1352_);
	assign _2198_ = _1859_ ^ _1352_;
	assign _2199_ = ~_1354_;
	assign _2200_ = ~(_1858_ & _2199_);
	assign _2201_ = _2198_ & ~_2200_;
	assign _2202_ = _2197_ & ~_2201_;
	assign _2204_ = _1858_ ^ _1354_;
	assign _2205_ = _2198_ & ~_2204_;
	assign _2206_ = _1869_ | _1355_;
	assign _2207_ = _1869_ ^ _1355_;
	assign _2208_ = ~(_1867_ | _1358_);
	assign _2209_ = _2207_ & ~_2208_;
	assign _2210_ = _2206_ & ~_2209_;
	assign _2211_ = _2205_ & ~_2210_;
	assign _2212_ = _2202_ & ~_2211_;
	assign _2213_ = _1349_ & ~_2212_;
	assign _2215_ = ~_2207_;
	assign _2216_ = _1867_ & _1358_;
	assign _2217_ = _2216_ | _2208_;
	assign _2218_ = _2217_ | _2215_;
	assign _2219_ = _2218_ | ~_2205_;
	assign _2220_ = _1349_ & ~_2219_;
	assign _2221_ = _2213_ & ~_2220_;
	assign _2222_ = _2221_ | _2196_;
	assign _2223_ = ~_1831_;
	assign _2224_ = (_1777_ ? _1781_ : _2223_);
	assign _2226_ = (_1257_ ? _2224_ : _2222_);
	assign _2227_ = ~(_1382_ & _1384_);
	assign _2228_ = ~(_1392_ & _1389_);
	assign _2229_ = ~(_2228_ | _2227_);
	assign _2230_ = _2229_ & ~_1402_;
	assign _2231_ = ~(_1472_ & _1425_);
	assign _2232_ = ~(_1509_ & _1503_);
	assign _2233_ = ~(_1495_ & _1489_);
	assign _2234_ = _2233_ | _2232_;
	assign _2235_ = ~(_1533_ & _1526_);
	assign _2237_ = ~(_1544_ & _1519_);
	assign _2238_ = _2237_ | _2235_;
	assign _2239_ = _2238_ | _2234_;
	assign _2240_ = _2239_ | _2231_;
	assign _2241_ = _2230_ & ~_2240_;
	assign _2242_ = (_2241_ ? _1764_ : _2226_);
	assign _2243_ = _1780_ & ~_2242_;
	assign _0055_ = (io_in[8] ? _2243_ : _1256_);
	assign _2244_ = ~_0307_;
	assign _2245_ = ~(_0351_ ^ _0286_);
	assign _2247_ = (_0358_ ? _2245_ : _1134_);
	assign _2248_ = _1223_ | _0881_;
	assign _2249_ = _0950_ & ~_1214_;
	assign _2250_ = _0843_ & ~_1217_;
	assign _2251_ = _2250_ | _2249_;
	assign _2252_ = _2248_ & ~_2251_;
	assign _2253_ = _1068_ & ~_1196_;
	assign _2254_ = _0981_ & ~_1201_;
	assign _2255_ = _2254_ | _2253_;
	assign _2256_ = _1013_ & ~_1206_;
	assign _2258_ = _0914_ & ~_1209_;
	assign _2259_ = _2258_ | _2256_;
	assign _2260_ = _2259_ | _2255_;
	assign _2261_ = _2252_ & ~_2260_;
	assign _2262_ = _1115_ & ~_1185_;
	assign _2263_ = ~_1041_;
	assign _2264_ = _1191_ & ~_2263_;
	assign _2265_ = _2264_ | _2262_;
	assign _2266_ = _2261_ & ~_2265_;
	assign _2267_ = _2266_ | _1242_;
	assign _2269_ = (_1252_ ? _1188_ : _2267_);
	assign _2270_ = (_0359_ ? _2247_ : _2269_);
	assign _2271_ = (_2137_ ? _2270_ : _2244_);
	assign _2272_ = _1132_ & ~_2271_;
	assign _2273_ = _2155_ | _2129_;
	assign _2274_ = ~(_2105_ | _2100_);
	assign _2275_ = _2273_ & ~_2274_;
	assign _2276_ = _2045_ & ~_2050_;
	assign _2277_ = ~(_2076_ | _2074_);
	assign _2278_ = _2277_ | _2276_;
	assign _2280_ = _2275_ & ~_2278_;
	assign _2281_ = _1931_ & ~_1962_;
	assign _2282_ = _1959_ & ~_1989_;
	assign _2283_ = _2282_ | _2281_;
	assign _2284_ = _1987_ & ~_2019_;
	assign _2285_ = _2015_ & ~_2021_;
	assign _2286_ = _2285_ | _2284_;
	assign _2287_ = _2286_ | _2283_;
	assign _2288_ = _2280_ & ~_2287_;
	assign _2289_ = _1831_ & ~_1871_;
	assign _2291_ = _1782_ & ~_1933_;
	assign _2292_ = _2291_ | _2289_;
	assign _2293_ = _2292_ | ~_2288_;
	assign _2294_ = (_2171_ ? _2154_ : _2293_);
	assign _2295_ = _2221_ | ~_2294_;
	assign _2296_ = (_1777_ ? _2223_ : _1842_);
	assign _2297_ = (_1257_ ? _2296_ : _2295_);
	assign _2298_ = (_2241_ ? _1756_ : _2297_);
	assign _2299_ = _1780_ & ~_2298_;
	assign _0062_ = (io_in[8] ? _2299_ : _2272_);
	assign _2301_ = ~_0284_;
	assign _2302_ = ~(_0351_ & _0286_);
	assign _2303_ = _2302_ ^ _0265_;
	assign _2304_ = (_0358_ ? _2303_ : _2245_);
	assign _2305_ = _1217_ | _0881_;
	assign _2306_ = _0843_ & ~_1214_;
	assign _2307_ = _2305_ & ~_2306_;
	assign _2308_ = _0981_ & ~_1196_;
	assign _2309_ = _1013_ & ~_1201_;
	assign _2310_ = _2309_ | _2308_;
	assign _2312_ = _0914_ & ~_1206_;
	assign _2313_ = _0950_ & ~_1209_;
	assign _2314_ = _2313_ | _2312_;
	assign _2315_ = _2314_ | _2310_;
	assign _2316_ = _2307_ & ~_2315_;
	assign _2317_ = _1041_ & ~_1185_;
	assign _2318_ = ~_1068_;
	assign _2319_ = _1191_ & ~_2318_;
	assign _2320_ = _2319_ | _2317_;
	assign _2321_ = _2316_ & ~_2320_;
	assign _2323_ = _2321_ | _1242_;
	assign _2324_ = (_1252_ ? _2263_ : _2323_);
	assign _2325_ = (_0359_ ? _2304_ : _2324_);
	assign _2326_ = (_2137_ ? _2325_ : _2301_);
	assign _2327_ = _1132_ & ~_2326_;
	assign _2328_ = _2155_ | _2100_;
	assign _2329_ = ~(_2105_ | _2074_);
	assign _2330_ = _2328_ & ~_2329_;
	assign _2331_ = _2015_ & ~_2050_;
	assign _2332_ = _2045_ & ~_2076_;
	assign _2334_ = _2332_ | _2331_;
	assign _2335_ = _2330_ & ~_2334_;
	assign _2336_ = _1782_ & ~_1962_;
	assign _2337_ = _1931_ & ~_1989_;
	assign _2338_ = _2337_ | _2336_;
	assign _2339_ = _1959_ & ~_2019_;
	assign _2340_ = _1987_ & ~_2021_;
	assign _2341_ = _2340_ | _2339_;
	assign _2342_ = _2341_ | _2338_;
	assign _2343_ = _2335_ & ~_2342_;
	assign _2345_ = _1830_ & ~_1871_;
	assign _2346_ = _1831_ & ~_1933_;
	assign _2347_ = _2346_ | _2345_;
	assign _2348_ = _2343_ & ~_2347_;
	assign _2349_ = (_2171_ ? _2129_ : _2348_);
	assign _2350_ = _2349_ | _2221_;
	assign _2351_ = ~_1821_;
	assign _2352_ = (_1777_ ? _1842_ : _2351_);
	assign _2353_ = (_1257_ ? _2352_ : _2350_);
	assign _2354_ = (_2241_ ? _1745_ : _2353_);
	assign _2356_ = _1780_ & ~_2354_;
	assign _0063_ = (io_in[8] ? _2356_ : _2327_);
	assign _2357_ = ~_0262_;
	assign _2358_ = ~_0245_;
	assign _2359_ = ~(_0352_ ^ _2358_);
	assign _2360_ = (_0358_ ? _2359_ : _2303_);
	assign _2361_ = _1214_ | _0881_;
	assign _2362_ = _1013_ & ~_1196_;
	assign _2363_ = _0914_ & ~_1201_;
	assign _2364_ = _2363_ | _2362_;
	assign _2366_ = _0950_ & ~_1206_;
	assign _2367_ = _0843_ & ~_1209_;
	assign _2368_ = _2367_ | _2366_;
	assign _2369_ = _2368_ | _2364_;
	assign _2370_ = _2361_ & ~_2369_;
	assign _2371_ = _1068_ & ~_1185_;
	assign _2372_ = ~_0981_;
	assign _2373_ = _1191_ & ~_2372_;
	assign _2374_ = _2373_ | _2371_;
	assign _2375_ = _2370_ & ~_2374_;
	assign _2377_ = _2375_ | _1242_;
	assign _2378_ = (_1252_ ? _2318_ : _2377_);
	assign _2379_ = (_0359_ ? _2360_ : _2378_);
	assign _2380_ = (_2137_ ? _2379_ : _2357_);
	assign _2381_ = _1132_ & ~_2380_;
	assign _2382_ = _2155_ | _2074_;
	assign _2383_ = _2045_ & ~_2105_;
	assign _2384_ = _2382_ & ~_2383_;
	assign _2385_ = _1987_ & ~_2050_;
	assign _2386_ = _2015_ & ~_2076_;
	assign _2388_ = _2386_ | _2385_;
	assign _2389_ = _2384_ & ~_2388_;
	assign _2390_ = _1831_ & ~_1962_;
	assign _2391_ = _1782_ & ~_1989_;
	assign _2392_ = _2391_ | _2390_;
	assign _2393_ = _1931_ & ~_2019_;
	assign _2394_ = _1959_ & ~_2021_;
	assign _2395_ = _2394_ | _2393_;
	assign _2396_ = _2395_ | _2392_;
	assign _2397_ = _2389_ & ~_2396_;
	assign _2399_ = _1821_ & ~_1871_;
	assign _2400_ = _1830_ & ~_1933_;
	assign _2401_ = _2400_ | _2399_;
	assign _2402_ = _2397_ & ~_2401_;
	assign _2403_ = (_2171_ ? _2100_ : _2402_);
	assign _2404_ = _2403_ | _2221_;
	assign _2405_ = ~_1813_;
	assign _2406_ = (_1777_ ? _2351_ : _2405_);
	assign _2407_ = (_1257_ ? _2406_ : _2404_);
	assign _2408_ = (_2241_ ? _1736_ : _2407_);
	assign _2410_ = _1780_ & ~_2408_;
	assign _0064_ = (io_in[8] ? _2410_ : _2381_);
	assign _2411_ = ~_0242_;
	assign _2412_ = _0352_ | _2358_;
	assign _2413_ = _2412_ ^ _0227_;
	assign _2414_ = (_0358_ ? _2413_ : _2359_);
	assign _2415_ = _1209_ | _0881_;
	assign _2416_ = _0843_ & ~_1206_;
	assign _2417_ = _2415_ & ~_2416_;
	assign _2418_ = _0914_ & ~_1196_;
	assign _2420_ = _0950_ & ~_1201_;
	assign _2421_ = _2420_ | _2418_;
	assign _2422_ = _2417_ & ~_2421_;
	assign _2423_ = _0981_ & ~_1185_;
	assign _2424_ = ~_1013_;
	assign _2425_ = _1191_ & ~_2424_;
	assign _2426_ = _2425_ | _2423_;
	assign _2427_ = _2422_ & ~_2426_;
	assign _2428_ = _2427_ | _1242_;
	assign _2429_ = (_1252_ ? _2372_ : _2428_);
	assign _2431_ = (_0359_ ? _2414_ : _2429_);
	assign _2432_ = (_2137_ ? _2431_ : _2411_);
	assign _2433_ = _1132_ & ~_2432_;
	assign _2434_ = ~_2045_;
	assign _2435_ = _2155_ | _2434_;
	assign _2436_ = _2015_ & ~_2105_;
	assign _2437_ = _2435_ & ~_2436_;
	assign _2438_ = _1959_ & ~_2050_;
	assign _2439_ = _1987_ & ~_2076_;
	assign _2440_ = _2439_ | _2438_;
	assign _2442_ = _2437_ & ~_2440_;
	assign _2443_ = _1830_ & ~_1962_;
	assign _2444_ = _1831_ & ~_1989_;
	assign _2445_ = _2444_ | _2443_;
	assign _2446_ = _1782_ & ~_2019_;
	assign _2447_ = _1931_ & ~_2021_;
	assign _2448_ = _2447_ | _2446_;
	assign _2449_ = _2448_ | _2445_;
	assign _2450_ = _2442_ & ~_2449_;
	assign _2451_ = _1813_ & ~_1871_;
	assign _2453_ = _1821_ & ~_1933_;
	assign _2454_ = _2453_ | _2451_;
	assign _2455_ = _2450_ & ~_2454_;
	assign _2456_ = (_2171_ ? _2074_ : _2455_);
	assign _2457_ = _2456_ | _2221_;
	assign _2458_ = ~_1804_;
	assign _2459_ = (_1777_ ? _2405_ : _2458_);
	assign _2460_ = (_1257_ ? _2459_ : _2457_);
	assign _2461_ = (_2241_ ? _1722_ : _2460_);
	assign _2462_ = _1780_ & ~_2461_;
	assign _0065_ = (io_in[8] ? _2462_ : _2433_);
	assign _2464_ = ~_0219_;
	assign _2465_ = ~(_0352_ | _0343_);
	assign _2466_ = _2465_ ^ _0341_;
	assign _2467_ = (_0358_ ? _2466_ : _2413_);
	assign _2468_ = _1206_ | _0881_;
	assign _2469_ = _0950_ & ~_1196_;
	assign _2470_ = _0843_ & ~_1201_;
	assign _2471_ = _2470_ | _2469_;
	assign _2472_ = _2468_ & ~_2471_;
	assign _2474_ = _1013_ & ~_1185_;
	assign _2475_ = ~_0914_;
	assign _2476_ = _1191_ & ~_2475_;
	assign _2477_ = _2476_ | _2474_;
	assign _2478_ = _2472_ & ~_2477_;
	assign _2479_ = _2478_ | _1242_;
	assign _2480_ = (_1252_ ? _2424_ : _2479_);
	assign _2481_ = (_0359_ ? _2467_ : _2480_);
	assign _2482_ = (_2137_ ? _2481_ : _2464_);
	assign _2483_ = _1132_ & ~_2482_;
	assign _2485_ = _2155_ | ~_2015_;
	assign _2486_ = _1987_ & ~_2105_;
	assign _2487_ = _2485_ & ~_2486_;
	assign _2488_ = _1931_ & ~_2050_;
	assign _2489_ = _1959_ & ~_2076_;
	assign _2490_ = _2489_ | _2488_;
	assign _2491_ = _2487_ & ~_2490_;
	assign _2492_ = _1821_ & ~_1962_;
	assign _2493_ = _1830_ & ~_1989_;
	assign _2494_ = _2493_ | _2492_;
	assign _2496_ = _1831_ & ~_2019_;
	assign _2497_ = _1782_ & ~_2021_;
	assign _2498_ = _2497_ | _2496_;
	assign _2499_ = _2498_ | _2494_;
	assign _2500_ = _2491_ & ~_2499_;
	assign _2501_ = _1804_ & ~_1871_;
	assign _2502_ = _1813_ & ~_1933_;
	assign _2503_ = _2502_ | _2501_;
	assign _2504_ = _2500_ & ~_2503_;
	assign _2505_ = (_2171_ ? _2434_ : _2504_);
	assign _2507_ = _2505_ | _2221_;
	assign _2508_ = ~_1790_;
	assign _2509_ = (_1777_ ? _2458_ : _2508_);
	assign _2510_ = (_1257_ ? _2509_ : _2507_);
	assign _2511_ = (_2241_ ? _1713_ : _2510_);
	assign _2512_ = _1780_ & ~_2511_;
	assign _0066_ = (io_in[8] ? _2512_ : _2483_);
	assign _2513_ = ~_0204_;
	assign _2514_ = ~(_2465_ & _0206_);
	assign _2515_ = _2514_ ^ _0193_;
	assign _2517_ = (_0358_ ? _2515_ : _2466_);
	assign _2518_ = _1201_ | _0881_;
	assign _2519_ = _0843_ & ~_1196_;
	assign _2520_ = _2518_ & ~_2519_;
	assign _2521_ = _0914_ & ~_1185_;
	assign _2522_ = ~_0950_;
	assign _2523_ = _1191_ & ~_2522_;
	assign _2524_ = _2523_ | _2521_;
	assign _2525_ = _2520_ & ~_2524_;
	assign _2526_ = _2525_ | _1242_;
	assign _2528_ = (_1252_ ? _2475_ : _2526_);
	assign _2529_ = (_0359_ ? _2517_ : _2528_);
	assign _2530_ = (_2137_ ? _2529_ : _2513_);
	assign _2531_ = _1132_ & ~_2530_;
	assign _2532_ = _2155_ | ~_1987_;
	assign _2533_ = _1959_ & ~_2105_;
	assign _2534_ = _2532_ & ~_2533_;
	assign _2535_ = _1782_ & ~_2050_;
	assign _2536_ = _1931_ & ~_2076_;
	assign _2537_ = _2536_ | _2535_;
	assign _2539_ = _2534_ & ~_2537_;
	assign _2540_ = _1813_ & ~_1962_;
	assign _2541_ = _1821_ & ~_1989_;
	assign _2542_ = _2541_ | _2540_;
	assign _2543_ = _1830_ & ~_2019_;
	assign _2544_ = _1831_ & ~_2021_;
	assign _2545_ = _2544_ | _2543_;
	assign _2546_ = _2545_ | _2542_;
	assign _2547_ = _2539_ & ~_2546_;
	assign _2548_ = _1790_ & ~_1871_;
	assign _2550_ = _1804_ & ~_1933_;
	assign _2551_ = _2550_ | _2548_;
	assign _2552_ = _2551_ | ~_2547_;
	assign _2553_ = (_2171_ ? _2015_ : _2552_);
	assign _2554_ = _2221_ | ~_2553_;
	assign _2555_ = ~_1789_;
	assign _2556_ = (_1777_ ? _2508_ : _2555_);
	assign _2557_ = (_1257_ ? _2556_ : _2554_);
	assign _2558_ = (_2241_ ? _1702_ : _2557_);
	assign _2559_ = _1780_ & ~_2558_;
	assign _0067_ = (io_in[8] ? _2559_ : _2531_);
	assign _2561_ = ~_0190_;
	assign _2562_ = ~(_0353_ ^ _0181_);
	assign _2563_ = (_0358_ ? _2562_ : _2515_);
	assign _2564_ = _1196_ | _0881_;
	assign _2565_ = _0950_ & ~_1185_;
	assign _2566_ = ~_0843_;
	assign _2567_ = _1191_ & ~_2566_;
	assign _2568_ = _2567_ | _2565_;
	assign _2569_ = _2564_ & ~_2568_;
	assign _2571_ = _2569_ | _1242_;
	assign _2572_ = (_1252_ ? _2522_ : _2571_);
	assign _2573_ = (_0359_ ? _2563_ : _2572_);
	assign _2574_ = (_2137_ ? _2573_ : _2561_);
	assign _2575_ = _1132_ & ~_2574_;
	assign _2576_ = ~_1692_;
	assign _2577_ = _2155_ | ~_1959_;
	assign _2578_ = _1931_ & ~_2105_;
	assign _2579_ = _2577_ & ~_2578_;
	assign _2580_ = _1831_ & ~_2050_;
	assign _2582_ = _1782_ & ~_2076_;
	assign _2583_ = _2582_ | _2580_;
	assign _2584_ = _2579_ & ~_2583_;
	assign _2585_ = _1804_ & ~_1962_;
	assign _2586_ = _1813_ & ~_1989_;
	assign _2587_ = _2586_ | _2585_;
	assign _2588_ = _1821_ & ~_2019_;
	assign _2589_ = _1830_ & ~_2021_;
	assign _2590_ = _2589_ | _2588_;
	assign _2591_ = _2590_ | _2587_;
	assign _2593_ = _2584_ & ~_2591_;
	assign _2594_ = _1789_ & ~_1871_;
	assign _2595_ = _1790_ & ~_1933_;
	assign _2596_ = _2595_ | _2594_;
	assign _2597_ = _2596_ | ~_2593_;
	assign _2598_ = (_2171_ ? _1987_ : _2597_);
	assign _2599_ = _2221_ | ~_2598_;
	assign _2600_ = (_1777_ ? _2555_ : _1795_);
	assign _2601_ = (_1257_ ? _2600_ : _2599_);
	assign _2602_ = (_2241_ ? _2576_ : _2601_);
	assign _2604_ = _1780_ & ~_2602_;
	assign _0068_ = (io_in[8] ? _2604_ : _2575_);
	assign _2605_ = ~_0179_;
	assign _2606_ = ~(_0353_ & _0181_);
	assign _2607_ = _2606_ ^ _0171_;
	assign _2608_ = (_0358_ ? _2607_ : _2562_);
	assign _2609_ = _0881_ | ~_1191_;
	assign _2610_ = _0843_ & ~_1185_;
	assign _2611_ = _2609_ & ~_2610_;
	assign _2612_ = _2611_ | _1242_;
	assign _2614_ = (_1252_ ? _2566_ : _2612_);
	assign _2615_ = (_0359_ ? _2608_ : _2614_);
	assign _2616_ = (_2137_ ? _2615_ : _2605_);
	assign _2617_ = _1132_ & ~_2616_;
	assign _2618_ = _2155_ | ~_1931_;
	assign _2619_ = _1782_ & ~_2105_;
	assign _2620_ = _2618_ & ~_2619_;
	assign _2621_ = _1830_ & ~_2050_;
	assign _2622_ = _1831_ & ~_2076_;
	assign _2623_ = _2622_ | _2621_;
	assign _2625_ = _2620_ & ~_2623_;
	assign _2626_ = _1790_ & ~_1962_;
	assign _2627_ = _1804_ & ~_1989_;
	assign _2628_ = _2627_ | _2626_;
	assign _2629_ = _1813_ & ~_2019_;
	assign _2630_ = _1821_ & ~_2021_;
	assign _2631_ = _2630_ | _2629_;
	assign _2632_ = _2631_ | _2628_;
	assign _2633_ = _2625_ & ~_2632_;
	assign _2634_ = _1797_ & ~_1871_;
	assign _2636_ = _1789_ & ~_1933_;
	assign _2637_ = _2636_ | _2634_;
	assign _2638_ = _2637_ | ~_2633_;
	assign _2639_ = (_2171_ ? _1959_ : _2638_);
	assign _2640_ = _2221_ | ~_2639_;
	assign _2641_ = ~_1794_;
	assign _2642_ = (_1777_ ? _1795_ : _2641_);
	assign _2643_ = (_1257_ ? _2642_ : _2640_);
	assign _2644_ = (_2241_ ? _1680_ : _2643_);
	assign _2645_ = _1780_ & ~_2644_;
	assign _0069_ = (io_in[8] ? _2645_ : _2617_);
	assign _2647_ = ~_0165_;
	assign _2648_ = (_0358_ ? _0356_ : _2607_);
	assign _2649_ = _1185_ | _0881_;
	assign _2650_ = (_1252_ ? _0881_ : _2649_);
	assign _2651_ = (_0359_ ? _2648_ : _2650_);
	assign _2652_ = (_2137_ ? _2651_ : _2647_);
	assign _2653_ = _1132_ & ~_2652_;
	assign _2654_ = _2155_ | ~_1782_;
	assign _2655_ = _1831_ & ~_2105_;
	assign _2657_ = _2654_ & ~_2655_;
	assign _2658_ = _1821_ & ~_2050_;
	assign _2659_ = _1830_ & ~_2076_;
	assign _2660_ = _2659_ | _2658_;
	assign _2661_ = _2657_ & ~_2660_;
	assign _2662_ = _1789_ & ~_1962_;
	assign _2663_ = _1790_ & ~_1989_;
	assign _2664_ = _2663_ | _2662_;
	assign _2665_ = _1804_ & ~_2019_;
	assign _2666_ = _1813_ & ~_2021_;
	assign _2668_ = _2666_ | _2665_;
	assign _2669_ = _2668_ | _2664_;
	assign _2670_ = _2661_ & ~_2669_;
	assign _2671_ = _1794_ & ~_1871_;
	assign _2672_ = _1797_ & ~_1933_;
	assign _2673_ = _2672_ | _2671_;
	assign _2674_ = _2673_ | ~_2670_;
	assign _2675_ = (_2171_ ? _1931_ : _2674_);
	assign _2676_ = _2221_ | ~_2675_;
	assign _2677_ = (_1777_ ? _2641_ : _1838_);
	assign _2679_ = (_1257_ ? _2677_ : _2676_);
	assign _2680_ = (_2241_ ? _1670_ : _2679_);
	assign _2681_ = _1780_ & ~_2680_;
	assign _0070_ = (io_in[8] ? _2681_ : _2653_);
	assign _2682_ = _1131_ | ~_2137_;
	assign _2683_ = _1252_ & ~_2682_;
	assign _2684_ = ~(_1157_ | _0359_);
	assign _2685_ = _0358_ ^ _0087_;
	assign _2686_ = ~(_2685_ ^ _2684_);
	assign _2687_ = _2686_ ^ _0359_;
	assign _2689_ = _2452_ & ~_2687_;
	assign _2690_ = _2683_ & ~_2689_;
	assign _2691_ = ~(_2103_ | _1960_);
	assign _2692_ = ~(_2691_ | _2221_);
	assign _2693_ = _2692_ & _2217_;
	assign _2694_ = _2241_ | _1777_;
	assign _2695_ = _2694_ | ~_1257_;
	assign _2696_ = ~(_2243_ ^ _1782_);
	assign _2697_ = _2299_ ^ _1831_;
	assign _2698_ = _2696_ & ~_2697_;
	assign _2700_ = _2410_ ^ _1821_;
	assign _2701_ = _2356_ ^ _1830_;
	assign _2702_ = _2701_ | _2700_;
	assign _2703_ = _2698_ & ~_2702_;
	assign _2704_ = _2604_ ^ _1789_;
	assign _2705_ = _2559_ ^ _1790_;
	assign _2706_ = _2705_ | _2704_;
	assign _2707_ = _2512_ ^ _1804_;
	assign _2708_ = _2462_ ^ _1813_;
	assign _2709_ = _2708_ | _2707_;
	assign _2711_ = _2709_ | _2706_;
	assign _2712_ = _2703_ & ~_2711_;
	assign _2713_ = _2681_ ^ _1794_;
	assign _2714_ = _2645_ ^ _1797_;
	assign _2715_ = _2714_ | _2713_;
	assign _2716_ = _2715_ | _1800_;
	assign _2717_ = _2712_ & ~_2716_;
	assign _2718_ = _2717_ ^ _1358_;
	assign _2719_ = _2718_ ^ _2695_;
	assign _2720_ = (_1257_ ? _2719_ : _2693_);
	assign _2722_ = _2720_ | ~_1780_;
	assign _0056_ = (io_in[8] ? _2722_ : _2690_);
	assign _2723_ = ~(_2686_ | _0359_);
	assign _2724_ = _0358_ & ~_0088_;
	assign _2725_ = _2685_ & _2684_;
	assign _2726_ = ~(_2725_ | _2724_);
	assign _2727_ = ~(_1145_ | _0359_);
	assign _2728_ = _2727_ ^ _0086_;
	assign _2729_ = _2728_ ^ _2726_;
	assign _2730_ = ~(_2729_ ^ _2723_);
	assign _2732_ = _2452_ & ~_2730_;
	assign _2733_ = _2683_ & ~_2732_;
	assign _2734_ = _2216_ ^ _2207_;
	assign _2735_ = _2692_ & ~_2734_;
	assign _2736_ = ~(_2718_ | _2695_);
	assign _2737_ = _1345_ ^ _1330_;
	assign _2738_ = _2717_ & _1358_;
	assign _2739_ = _2738_ ^ _2737_;
	assign _2740_ = ~(_2739_ ^ _2736_);
	assign _2741_ = (_1257_ ? _2740_ : _2735_);
	assign _2743_ = _2741_ | ~_1780_;
	assign _0057_ = (io_in[8] ? _2743_ : _2733_);
	assign _2744_ = _2723_ & ~_2729_;
	assign _2745_ = _2728_ & ~_2726_;
	assign _2746_ = _2745_ | _2744_;
	assign _2747_ = _2727_ & _0086_;
	assign _2748_ = ~(_1138_ | _0359_);
	assign _2749_ = _2748_ ^ _0085_;
	assign _2750_ = _2749_ ^ _2747_;
	assign _2751_ = _2750_ ^ _2746_;
	assign _2753_ = _2452_ & ~_2751_;
	assign _2754_ = _2683_ & ~_2753_;
	assign _2755_ = _2216_ | ~_2207_;
	assign _2756_ = _1869_ & ~_2737_;
	assign _2757_ = _2755_ & ~_2756_;
	assign _2758_ = ~(_2757_ ^ _2204_);
	assign _2759_ = _2692_ & ~_2758_;
	assign _2760_ = _2737_ & ~_2738_;
	assign _2761_ = _2736_ & ~_2739_;
	assign _2762_ = _2761_ | _2760_;
	assign _2764_ = _2737_ ^ _1354_;
	assign _2765_ = _2764_ ^ _2762_;
	assign _2766_ = (_1257_ ? _2765_ : _2759_);
	assign _2767_ = _2766_ | ~_1780_;
	assign _0058_ = (io_in[8] ? _2767_ : _2754_);
	assign _2768_ = _2749_ & _2747_;
	assign _2769_ = _2750_ & _2746_;
	assign _2770_ = _2769_ | _2768_;
	assign _2771_ = _2748_ & _0085_;
	assign _2772_ = ~(_1167_ | _0359_);
	assign _2774_ = _2772_ ^ _0084_;
	assign _2775_ = _2774_ ^ _2771_;
	assign _2776_ = _2775_ ^ _2770_;
	assign _2777_ = _2452_ & ~_2776_;
	assign _2778_ = _2683_ & ~_2777_;
	assign _2779_ = _2757_ | _2204_;
	assign _2780_ = _1354_ & ~_1858_;
	assign _2781_ = _2779_ & ~_2780_;
	assign _2782_ = _2781_ ^ _2198_;
	assign _2783_ = _2692_ & ~_2782_;
	assign _2785_ = _1355_ & ~_1354_;
	assign _2786_ = _2764_ & _2762_;
	assign _2787_ = _2786_ | _2785_;
	assign _2788_ = _1354_ ^ _1352_;
	assign _2789_ = _2788_ ^ _2787_;
	assign _2790_ = (_1257_ ? _2789_ : _2783_);
	assign _2791_ = _2790_ | ~_1780_;
	assign _0059_ = (io_in[8] ? _2791_ : _2778_);
	assign _2792_ = _2774_ & _2771_;
	assign _2793_ = _2775_ & _2768_;
	assign _2795_ = _2793_ | _2792_;
	assign _2796_ = ~(_2775_ & _2750_);
	assign _2797_ = _2746_ & ~_2796_;
	assign _2798_ = _2797_ | _2795_;
	assign _2799_ = _2772_ & _0084_;
	assign _2800_ = ~(_1182_ | _0359_);
	assign _2801_ = _2800_ ^ _0102_;
	assign _2802_ = _2801_ ^ _2799_;
	assign _2803_ = _2802_ ^ _2798_;
	assign _2804_ = _2452_ & ~_2803_;
	assign _2806_ = _2683_ & ~_2804_;
	assign _2807_ = _1859_ | _1352_;
	assign _2808_ = _2780_ & _2198_;
	assign _2809_ = _2807_ & ~_2808_;
	assign _2810_ = _2205_ & ~_2757_;
	assign _2811_ = _2809_ & ~_2810_;
	assign _2812_ = _2811_ ^ _1349_;
	assign _2813_ = _2692_ & ~_2812_;
	assign _2814_ = _1352_ & ~_2199_;
	assign _2815_ = _2788_ & _2785_;
	assign _2817_ = _2815_ | _2814_;
	assign _2818_ = ~(_2788_ & _2764_);
	assign _2819_ = _2762_ & ~_2818_;
	assign _2820_ = _2819_ | _2817_;
	assign _2821_ = ~(_1352_ ^ _1349_);
	assign _2822_ = _2821_ ^ _2820_;
	assign _2823_ = (_1257_ ? _2822_ : _2813_);
	assign _2824_ = _2823_ | ~_1780_;
	assign _0060_ = (io_in[8] ? _2824_ : _2806_);
	assign _2825_ = \mchip.value_A [15] ^ \mchip.value_B [15];
	assign _2827_ = (_1313_ ? \mchip.value_B [15] : \mchip.value_A [15]);
	assign _2828_ = (_1268_ ? \mchip.value_A [15] : _2827_);
	assign _2829_ = (_1329_ ? \mchip.value_B [15] : _2828_);
	assign _0061_ = (io_in[8] ? _2829_ : _2825_);
	assign _2830_ = _2419_ | _2387_;
	assign _2831_ = _2246_ & ~_2279_;
	assign \mchip.temp_valid_add  = _2830_ & ~_2831_;
	assign _2832_ = ~\mchip.j [1];
	assign _2833_ = ~(\mchip.j [1] | \mchip.j [2]);
	assign _2834_ = _2833_ ^ \mchip.j [3];
	assign _2836_ = ~(\mchip.j [1] ^ \mchip.j [2]);
	assign _2837_ = _2836_ | _2834_;
	assign _2838_ = \mchip.j [1] & ~_2837_;
	assign _2839_ = \mchip.j [3] | \mchip.j [2];
	assign _2840_ = _2832_ & ~_2839_;
	assign _2841_ = _2840_ ^ \mchip.j [4];
	assign _2842_ = _2838_ & ~_2841_;
	assign _2843_ = _2840_ & ~\mchip.j [4];
	assign _2844_ = ~(_2843_ ^ \mchip.j [5]);
	assign _2845_ = _2844_ ^ _2842_;
	assign _2847_ = ~\mchip.j [30];
	assign _2848_ = \mchip.j [5] | \mchip.j [4];
	assign _2849_ = _2848_ | \mchip.j [30];
	assign _2850_ = _2840_ & ~_2849_;
	assign _2851_ = _2847_ & ~_2850_;
	assign _2852_ = _2840_ & ~_2848_;
	assign _2853_ = _2847_ & ~_2852_;
	assign _2854_ = _2841_ | ~_2844_;
	assign _2855_ = _2854_ | ~_2853_;
	assign _2856_ = _2838_ & ~_2855_;
	assign _2858_ = _2851_ & ~_2856_;
	assign _2859_ = _2858_ ^ _2845_;
	assign _2861_ = _2850_ ^ \mchip.j [30];
	assign _2862_ = _2856_ & ~_2861_;
	assign _2863_ = _2862_ ^ _2851_;
	assign _2864_ = _2863_ ^ _2845_;
	assign _2865_ = ~(_2861_ ^ _2856_);
	assign _2866_ = _2865_ ^ _2845_;
	assign _2867_ = _2838_ & ~_2854_;
	assign _2868_ = _2852_ ^ \mchip.j [30];
	assign _2869_ = _2867_ & ~_2868_;
	assign _2870_ = _2869_ ^ _2853_;
	assign _2872_ = _2870_ ^ _2845_;
	assign _2873_ = ~(_2868_ ^ _2867_);
	assign _2874_ = _2873_ ^ _2845_;
	assign _2875_ = _2874_ | _2872_;
	assign _2876_ = _2875_ | _2866_;
	assign _2877_ = _2876_ | _2864_;
	assign _2878_ = _2877_ | _2859_;
	assign _2879_ = _2878_ | _2859_;
	assign _2880_ = _2879_ | _2859_;
	assign _2881_ = _2880_ | _2859_;
	assign _2883_ = _2881_ | _2859_;
	assign _2884_ = _2883_ | _2859_;
	assign _2885_ = _2884_ | _2859_;
	assign _2886_ = _2885_ | _2859_;
	assign _2887_ = _2886_ | _2859_;
	assign _2888_ = _2887_ | _2859_;
	assign _2889_ = _2888_ | _2859_;
	assign _2890_ = _2889_ | _2859_;
	assign _2891_ = _2890_ | _2859_;
	assign _2892_ = _2891_ | _2859_;
	assign _2894_ = _2892_ | _2859_;
	assign _2895_ = _2894_ | _2859_;
	assign _2896_ = _2895_ | _2859_;
	assign _2897_ = _2896_ | _2859_;
	assign _2898_ = _2897_ | ~io_in[7];
	assign _2899_ = ~(_2898_ | _2845_);
	assign _2900_ = _2897_ | ~io_in[5];
	assign _2901_ = ~(_2900_ | _2845_);
	assign _2902_ = ~_2845_;
	assign _2903_ = _2897_ | ~io_in[4];
	assign _2905_ = _2902_ & ~_2903_;
	assign _2906_ = (\mchip.j [1] ? _2905_ : _2901_);
	assign _2907_ = (\mchip.j [1] ? _2906_ : _2899_);
	assign _2908_ = _2836_ ^ \mchip.j [1];
	assign _2909_ = ~_2908_;
	assign _2910_ = _2907_ & ~_2909_;
	assign _2911_ = \mchip.j [3] ^ \mchip.j [2];
	assign _2912_ = _2910_ & ~_2911_;
	assign _2913_ = _2841_ ^ _2838_;
	assign _2914_ = ~_2913_;
	assign _2916_ = _2912_ & ~_2914_;
	assign _2917_ = ~_2911_;
	assign _2918_ = _2897_ | _2845_;
	assign _2919_ = _2918_ | \mchip.j [1];
	assign _2920_ = \mchip.j [1] & ~_2918_;
	assign _2921_ = _2919_ & ~_2920_;
	assign _2922_ = _2921_ | _2909_;
	assign _2923_ = _2922_ | ~_2917_;
	assign _2924_ = ~(_2923_ | _2914_);
	assign _2925_ = \mchip.tmp_input_B [0] & ~_2924_;
	assign _0026_ = _2925_ | _2916_;
	assign _2927_ = ~(_2901_ & \mchip.j [1]);
	assign _2928_ = _2927_ | _2909_;
	assign _2929_ = _2917_ & ~_2928_;
	assign _2930_ = _2903_ | _2902_;
	assign _2931_ = _2930_ | \mchip.j [1];
	assign _2932_ = _2931_ | _2908_;
	assign _2933_ = _2911_ & ~_2932_;
	assign _2934_ = (_2913_ ? _2929_ : _2933_);
	assign _2935_ = ~(_2920_ & _2908_);
	assign _2937_ = _2917_ & ~_2935_;
	assign _2938_ = _2897_ | _2902_;
	assign _2939_ = _2938_ | \mchip.j [1];
	assign _2940_ = _2939_ | ~_2909_;
	assign _2941_ = ~(_2940_ | _2917_);
	assign _2942_ = (_2913_ ? _2937_ : _2941_);
	assign _2943_ = \mchip.tmp_input_B [1] & ~_2942_;
	assign _0033_ = _2943_ | _2934_;
	assign _2944_ = _2897_ | ~io_in[6];
	assign _2945_ = ~(_2944_ | _2845_);
	assign _2947_ = (\mchip.j [1] ? _2945_ : _2899_);
	assign _2948_ = ~(_2947_ & \mchip.j [1]);
	assign _2949_ = _2948_ | _2909_;
	assign _2950_ = _2917_ & ~_2949_;
	assign _2951_ = _2900_ | ~_2845_;
	assign _2952_ = (\mchip.j [1] ? _2930_ : _2951_);
	assign _2953_ = _2952_ | \mchip.j [1];
	assign _2954_ = _2953_ | ~_2909_;
	assign _2955_ = ~(_2954_ | _2917_);
	assign _2956_ = (_2913_ ? _2950_ : _2955_);
	assign _2958_ = \mchip.tmp_input_B [2] & ~_2942_;
	assign _0034_ = _2958_ | _2956_;
	assign _2959_ = ~(_2899_ & \mchip.j [1]);
	assign _2960_ = _2959_ | _2909_;
	assign _2961_ = _2917_ & ~_2960_;
	assign _2962_ = _2944_ | ~_2845_;
	assign _2963_ = (\mchip.j [1] ? _2951_ : _2962_);
	assign _2964_ = (\mchip.j [1] ? _2931_ : _2963_);
	assign _2965_ = _2964_ | _2908_;
	assign _2966_ = _2911_ & ~_2965_;
	assign _2968_ = (_2913_ ? _2961_ : _2966_);
	assign _2969_ = \mchip.tmp_input_B [3] & ~_2942_;
	assign _0035_ = _2969_ | _2968_;
	assign _2970_ = _2898_ | ~_2845_;
	assign _2971_ = (\mchip.j [1] ? _2962_ : _2970_);
	assign _2972_ = (\mchip.j [1] ? _2952_ : _2971_);
	assign _2973_ = _2972_ | ~_2909_;
	assign _2974_ = _2973_ | _2917_;
	assign _2975_ = _2914_ & ~_2974_;
	assign _2976_ = _2938_ | _2832_;
	assign _2978_ = _2976_ & _2939_;
	assign _2979_ = _2978_ | ~_2909_;
	assign _2980_ = _2979_ | _2917_;
	assign _2981_ = _2914_ & ~_2980_;
	assign _2982_ = \mchip.tmp_input_B [4] & ~_2981_;
	assign _0036_ = _2982_ | _2975_;
	assign _2983_ = _2963_ | _2832_;
	assign _2984_ = (_2908_ ? _2931_ : _2983_);
	assign _2985_ = _2984_ | _2917_;
	assign _2986_ = _2914_ & ~_2985_;
	assign _2988_ = (_2908_ ? _2939_ : _2976_);
	assign _2989_ = _2988_ | _2917_;
	assign _2990_ = _2914_ & ~_2989_;
	assign _2991_ = \mchip.tmp_input_B [5] & ~_2990_;
	assign _0037_ = _2991_ | _2986_;
	assign _2992_ = _2962_ | _2832_;
	assign _2993_ = (_2908_ ? _2953_ : _2992_);
	assign _2994_ = _2993_ | _2917_;
	assign _2995_ = _2914_ & ~_2994_;
	assign _2996_ = \mchip.tmp_input_B [6] & ~_2990_;
	assign _0038_ = _2996_ | _2995_;
	assign _2998_ = _2970_ | _2832_;
	assign _2999_ = (_2908_ ? _2964_ : _2998_);
	assign _3000_ = _2999_ | _2917_;
	assign _3001_ = _2914_ & ~_3000_;
	assign _3002_ = \mchip.tmp_input_B [7] & ~_2990_;
	assign _0039_ = _3002_ | _3001_;
	assign _3003_ = _2972_ | _2909_;
	assign _3004_ = _3003_ | _2917_;
	assign _3005_ = _2914_ & ~_3004_;
	assign _3007_ = _2978_ | _2909_;
	assign _3008_ = _3007_ | _2917_;
	assign _3009_ = _2914_ & ~_3008_;
	assign _3010_ = \mchip.tmp_input_B [8] & ~_3009_;
	assign _0040_ = _3010_ | _3005_;
	assign _3011_ = _2983_ | _2909_;
	assign _3012_ = (_2911_ ? _3011_ : _2932_);
	assign _3013_ = _2914_ & ~_3012_;
	assign _3014_ = _2976_ | _2909_;
	assign _3015_ = (_2911_ ? _3014_ : _2940_);
	assign _3017_ = _2914_ & ~_3015_;
	assign _3018_ = \mchip.tmp_input_B [9] & ~_3017_;
	assign _0041_ = _3018_ | _3013_;
	assign _3019_ = _2992_ | _2909_;
	assign _3020_ = (_2911_ ? _3019_ : _2954_);
	assign _3021_ = _2914_ & ~_3020_;
	assign _3022_ = \mchip.tmp_input_B [10] & ~_3017_;
	assign _0027_ = _3022_ | _3021_;
	assign _3023_ = _2998_ | _2909_;
	assign _3024_ = (_2911_ ? _3023_ : _2965_);
	assign _3026_ = _2914_ & ~_3024_;
	assign _3027_ = \mchip.tmp_input_B [11] & ~_3017_;
	assign _0028_ = _3027_ | _3026_;
	assign _3028_ = _2973_ | ~_2917_;
	assign _3029_ = _2914_ & ~_3028_;
	assign _3030_ = _2979_ | ~_2917_;
	assign _3031_ = _2914_ & ~_3030_;
	assign _3032_ = \mchip.tmp_input_B [12] & ~_3031_;
	assign _0029_ = _3032_ | _3029_;
	assign _3033_ = _2984_ | ~_2917_;
	assign _3035_ = _2914_ & ~_3033_;
	assign _3036_ = _2988_ | ~_2917_;
	assign _3037_ = _2914_ & ~_3036_;
	assign _3038_ = \mchip.tmp_input_B [13] & ~_3037_;
	assign _0030_ = _3038_ | _3035_;
	assign _3039_ = _2993_ | ~_2917_;
	assign _3040_ = _2914_ & ~_3039_;
	assign _3041_ = \mchip.tmp_input_B [14] & ~_3037_;
	assign _0031_ = _3041_ | _3040_;
	assign _3042_ = _2999_ | ~_2917_;
	assign _3044_ = _2914_ & ~_3042_;
	assign _3045_ = \mchip.tmp_input_B [15] & ~_3037_;
	assign _0032_ = _3045_ | _3044_;
	assign _3046_ = _2897_ | ~io_in[3];
	assign _3047_ = _3046_ | _2845_;
	assign _3048_ = _2897_ | ~io_in[1];
	assign _3049_ = _3048_ | _2845_;
	assign _3050_ = _2897_ | ~io_in[0];
	assign _3051_ = _3050_ | _2845_;
	assign _3052_ = (\mchip.j [1] ? _3051_ : _3049_);
	assign _3054_ = (\mchip.j [1] ? _3052_ : _3047_);
	assign _3055_ = _3054_ | _2909_;
	assign _3056_ = _3055_ | _2911_;
	assign _3057_ = _2913_ & ~_3056_;
	assign _3058_ = \mchip.tmp_input_A [0] & ~_2924_;
	assign _0010_ = _3058_ | _3057_;
	assign _3059_ = _3049_ | _2832_;
	assign _3060_ = _3059_ | _2909_;
	assign _3061_ = _2917_ & ~_3060_;
	assign _3062_ = _3050_ | _2902_;
	assign _3064_ = _3062_ | \mchip.j [1];
	assign _3065_ = _3064_ | _2908_;
	assign _3066_ = _2911_ & ~_3065_;
	assign _3067_ = (_2913_ ? _3061_ : _3066_);
	assign _3068_ = \mchip.tmp_input_A [1] & ~_2942_;
	assign _0017_ = _3068_ | _3067_;
	assign _3069_ = _2897_ | ~io_in[2];
	assign _3070_ = _3069_ | _2845_;
	assign _3071_ = (\mchip.j [1] ? _3070_ : _3047_);
	assign _3072_ = _3071_ | _2832_;
	assign _3074_ = _3072_ | _2909_;
	assign _3075_ = _2917_ & ~_3074_;
	assign _3076_ = _3048_ | _2902_;
	assign _3077_ = (\mchip.j [1] ? _3062_ : _3076_);
	assign _3078_ = _3077_ | \mchip.j [1];
	assign _3079_ = _3078_ | ~_2909_;
	assign _3080_ = ~(_3079_ | _2917_);
	assign _3081_ = (_2913_ ? _3075_ : _3080_);
	assign _3082_ = \mchip.tmp_input_A [2] & ~_2942_;
	assign _0018_ = _3082_ | _3081_;
	assign _3084_ = _3047_ | _2832_;
	assign _3085_ = _3084_ | _2909_;
	assign _3086_ = _2917_ & ~_3085_;
	assign _3087_ = _3069_ | ~_2845_;
	assign _3088_ = (\mchip.j [1] ? _3076_ : _3087_);
	assign _3089_ = (\mchip.j [1] ? _3064_ : _3088_);
	assign _3090_ = _3089_ | _2908_;
	assign _3091_ = _2911_ & ~_3090_;
	assign _3092_ = (_2913_ ? _3086_ : _3091_);
	assign _3093_ = \mchip.tmp_input_A [3] & ~_2942_;
	assign _0019_ = _3093_ | _3092_;
	assign _3095_ = _3046_ | _2902_;
	assign _3096_ = (\mchip.j [1] ? _3087_ : _3095_);
	assign _3097_ = (\mchip.j [1] ? _3077_ : _3096_);
	assign _3098_ = _3097_ | ~_2909_;
	assign _3099_ = _3098_ | _2917_;
	assign _3100_ = _2914_ & ~_3099_;
	assign _3101_ = \mchip.tmp_input_A [4] & ~_2981_;
	assign _0020_ = _3101_ | _3100_;
	assign _3102_ = _3088_ | _2832_;
	assign _3104_ = (_2908_ ? _3064_ : _3102_);
	assign _3105_ = _3104_ | _2917_;
	assign _3106_ = _2914_ & ~_3105_;
	assign _3107_ = \mchip.tmp_input_A [5] & ~_2990_;
	assign _0021_ = _3107_ | _3106_;
	assign _3108_ = _3087_ | _2832_;
	assign _3109_ = (_2908_ ? _3078_ : _3108_);
	assign _3110_ = _3109_ | _2917_;
	assign _3111_ = _2914_ & ~_3110_;
	assign _3112_ = \mchip.tmp_input_A [6] & ~_2990_;
	assign _0022_ = _3112_ | _3111_;
	assign _3114_ = _3095_ | _2832_;
	assign _3115_ = (_2908_ ? _3089_ : _3114_);
	assign _3116_ = _3115_ | _2917_;
	assign _3117_ = _2914_ & ~_3116_;
	assign _3118_ = \mchip.tmp_input_A [7] & ~_2990_;
	assign _0023_ = _3118_ | _3117_;
	assign _3119_ = _3097_ | _2909_;
	assign _3120_ = _3119_ | _2917_;
	assign _3121_ = _2914_ & ~_3120_;
	assign _3123_ = \mchip.tmp_input_A [8] & ~_3009_;
	assign _0024_ = _3123_ | _3121_;
	assign _3124_ = _3102_ | _2909_;
	assign _3125_ = (_2911_ ? _3124_ : _3065_);
	assign _3126_ = _2914_ & ~_3125_;
	assign _3127_ = \mchip.tmp_input_A [9] & ~_3017_;
	assign _0025_ = _3127_ | _3126_;
	assign _3128_ = _3108_ | _2909_;
	assign _3129_ = (_2911_ ? _3128_ : _3079_);
	assign _3130_ = _2914_ & ~_3129_;
	assign _3132_ = \mchip.tmp_input_A [10] & ~_3017_;
	assign _0011_ = _3132_ | _3130_;
	assign _3133_ = _3114_ | _2909_;
	assign _3134_ = (_2911_ ? _3133_ : _3090_);
	assign _3135_ = _2914_ & ~_3134_;
	assign _3136_ = \mchip.tmp_input_A [11] & ~_3017_;
	assign _0012_ = _3136_ | _3135_;
	assign _3137_ = _3098_ | ~_2917_;
	assign _3138_ = _2914_ & ~_3137_;
	assign _3139_ = \mchip.tmp_input_A [12] & ~_3031_;
	assign _0013_ = _3139_ | _3138_;
	assign _3141_ = _3104_ | ~_2917_;
	assign _3142_ = _2914_ & ~_3141_;
	assign _3143_ = \mchip.tmp_input_A [13] & ~_3037_;
	assign _0014_ = _3143_ | _3142_;
	assign _3144_ = _3109_ | ~_2917_;
	assign _3145_ = _2914_ & ~_3144_;
	assign _3146_ = \mchip.tmp_input_A [14] & ~_3037_;
	assign _0015_ = _3146_ | _3145_;
	assign _3147_ = _3115_ | _2911_;
	assign _3149_ = _2914_ & ~_3147_;
	assign _3150_ = \mchip.tmp_input_A [15] & ~_3037_;
	assign _0016_ = _3150_ | _3149_;
	assign _3758_[2] = _0942_ ^ \mchip.count [2];
	assign _3151_ = _0942_ & ~\mchip.count [2];
	assign _3758_[3] = _3151_ ^ \mchip.count [3];
	reg \mchip.io_out_reg[8] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.io_out_reg[8]  <= 1'h0;
		else if (_0009_)
			\mchip.io_out_reg[8]  <= _0042_;
	assign \mchip.io_out [8] = \mchip.io_out_reg[8] ;
	always @(posedge io_in[12])
		if (_0007_)
			\mchip.value_B [0] <= \mchip.tmp_input_B [0];
	always @(posedge io_in[12])
		if (_0007_)
			\mchip.value_B [1] <= \mchip.tmp_input_B [1];
	always @(posedge io_in[12])
		if (_0007_)
			\mchip.value_B [2] <= \mchip.tmp_input_B [2];
	always @(posedge io_in[12])
		if (_0007_)
			\mchip.value_B [3] <= \mchip.tmp_input_B [3];
	always @(posedge io_in[12])
		if (_0007_)
			\mchip.value_B [4] <= \mchip.tmp_input_B [4];
	always @(posedge io_in[12])
		if (_0007_)
			\mchip.value_B [5] <= \mchip.tmp_input_B [5];
	always @(posedge io_in[12])
		if (_0007_)
			\mchip.value_B [6] <= \mchip.tmp_input_B [6];
	always @(posedge io_in[12])
		if (_0007_)
			\mchip.value_B [7] <= \mchip.tmp_input_B [7];
	always @(posedge io_in[12])
		if (_0007_)
			\mchip.value_B [8] <= \mchip.tmp_input_B [8];
	always @(posedge io_in[12])
		if (_0007_)
			\mchip.value_B [9] <= \mchip.tmp_input_B [9];
	always @(posedge io_in[12])
		if (_0007_)
			\mchip.value_B [10] <= \mchip.tmp_input_B [10];
	always @(posedge io_in[12])
		if (_0007_)
			\mchip.value_B [11] <= \mchip.tmp_input_B [11];
	always @(posedge io_in[12])
		if (_0007_)
			\mchip.value_B [12] <= \mchip.tmp_input_B [12];
	always @(posedge io_in[12])
		if (_0007_)
			\mchip.value_B [13] <= \mchip.tmp_input_B [13];
	always @(posedge io_in[12])
		if (_0007_)
			\mchip.value_B [14] <= \mchip.tmp_input_B [14];
	always @(posedge io_in[12])
		if (_0007_)
			\mchip.value_B [15] <= \mchip.tmp_input_B [15];
	always @(posedge io_in[12]) \mchip.i [0] <= _0000_;
	always @(posedge io_in[12]) \mchip.i [1] <= _0001_;
	always @(posedge io_in[12]) \mchip.i [2] <= _0002_;
	always @(posedge io_in[12]) \mchip.i [3] <= _0003_;
	reg \mchip.j_reg[1] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.j_reg[1]  <= 1'h0;
		else if (_0004_)
			\mchip.j_reg[1]  <= 1'h1;
	assign \mchip.j [1] = \mchip.j_reg[1] ;
	reg \mchip.j_reg[2] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.j_reg[2]  <= 1'h0;
		else if (_0004_)
			\mchip.j_reg[2]  <= _3757_[0];
	assign \mchip.j [2] = \mchip.j_reg[2] ;
	reg \mchip.j_reg[3] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.j_reg[3]  <= 1'h0;
		else if (_0004_)
			\mchip.j_reg[3]  <= _3758_[1];
	assign \mchip.j [3] = \mchip.j_reg[3] ;
	reg \mchip.j_reg[4] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.j_reg[4]  <= 1'h0;
		else if (_0004_)
			\mchip.j_reg[4]  <= _3758_[2];
	assign \mchip.j [4] = \mchip.j_reg[4] ;
	reg \mchip.j_reg[5] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.j_reg[5]  <= 1'h0;
		else if (_0004_)
			\mchip.j_reg[5]  <= _3758_[3];
	assign \mchip.j [5] = \mchip.j_reg[5] ;
	reg \mchip.j_reg[30] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.j_reg[30]  <= 1'h0;
		else if (_0004_)
			\mchip.j_reg[30]  <= _3758_[4];
	assign \mchip.j [30] = \mchip.j_reg[30] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.count [0] <= 1'h1;
		else if (_0005_)
			\mchip.count [0] <= _0051_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.count [1] <= 1'h0;
		else if (_0005_)
			\mchip.count [1] <= _0052_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.count [2] <= 1'h0;
		else if (_0005_)
			\mchip.count [2] <= _0053_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.count [3] <= 1'h0;
		else if (_0005_)
			\mchip.count [3] <= _0054_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.valid  <= 1'h0;
		else if (_0006_)
			\mchip.valid  <= \mchip.temp_valid_add ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.result [0] <= 1'h0;
		else if (_0006_)
			\mchip.result [0] <= _0055_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.result [1] <= 1'h0;
		else if (_0006_)
			\mchip.result [1] <= _0062_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.result [2] <= 1'h0;
		else if (_0006_)
			\mchip.result [2] <= _0063_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.result [3] <= 1'h0;
		else if (_0006_)
			\mchip.result [3] <= _0064_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.result [4] <= 1'h0;
		else if (_0006_)
			\mchip.result [4] <= _0065_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.result [5] <= 1'h0;
		else if (_0006_)
			\mchip.result [5] <= _0066_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.result [6] <= 1'h0;
		else if (_0006_)
			\mchip.result [6] <= _0067_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.result [7] <= 1'h0;
		else if (_0006_)
			\mchip.result [7] <= _0068_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.result [8] <= 1'h0;
		else if (_0006_)
			\mchip.result [8] <= _0069_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.result [9] <= 1'h0;
		else if (_0006_)
			\mchip.result [9] <= _0070_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.result [10] <= 1'h0;
		else if (_0006_)
			\mchip.result [10] <= _0056_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.result [11] <= 1'h0;
		else if (_0006_)
			\mchip.result [11] <= _0057_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.result [12] <= 1'h0;
		else if (_0006_)
			\mchip.result [12] <= _0058_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.result [13] <= 1'h0;
		else if (_0006_)
			\mchip.result [13] <= _0059_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.result [14] <= 1'h0;
		else if (_0006_)
			\mchip.result [14] <= _0060_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.result [15] <= 1'h0;
		else if (_0006_)
			\mchip.result [15] <= _0061_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.tmp_input_B [0] <= 1'h0;
		else if (_0004_)
			\mchip.tmp_input_B [0] <= _0026_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.tmp_input_B [1] <= 1'h0;
		else if (_0004_)
			\mchip.tmp_input_B [1] <= _0033_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.tmp_input_B [2] <= 1'h0;
		else if (_0004_)
			\mchip.tmp_input_B [2] <= _0034_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.tmp_input_B [3] <= 1'h0;
		else if (_0004_)
			\mchip.tmp_input_B [3] <= _0035_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.tmp_input_B [4] <= 1'h0;
		else if (_0004_)
			\mchip.tmp_input_B [4] <= _0036_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.tmp_input_B [5] <= 1'h0;
		else if (_0004_)
			\mchip.tmp_input_B [5] <= _0037_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.tmp_input_B [6] <= 1'h0;
		else if (_0004_)
			\mchip.tmp_input_B [6] <= _0038_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.tmp_input_B [7] <= 1'h0;
		else if (_0004_)
			\mchip.tmp_input_B [7] <= _0039_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.tmp_input_B [8] <= 1'h0;
		else if (_0004_)
			\mchip.tmp_input_B [8] <= _0040_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.tmp_input_B [9] <= 1'h0;
		else if (_0004_)
			\mchip.tmp_input_B [9] <= _0041_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.tmp_input_B [10] <= 1'h0;
		else if (_0004_)
			\mchip.tmp_input_B [10] <= _0027_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.tmp_input_B [11] <= 1'h0;
		else if (_0004_)
			\mchip.tmp_input_B [11] <= _0028_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.tmp_input_B [12] <= 1'h0;
		else if (_0004_)
			\mchip.tmp_input_B [12] <= _0029_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.tmp_input_B [13] <= 1'h0;
		else if (_0004_)
			\mchip.tmp_input_B [13] <= _0030_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.tmp_input_B [14] <= 1'h0;
		else if (_0004_)
			\mchip.tmp_input_B [14] <= _0031_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.tmp_input_B [15] <= 1'h0;
		else if (_0004_)
			\mchip.tmp_input_B [15] <= _0032_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.tmp_input_A [0] <= 1'h0;
		else if (_0004_)
			\mchip.tmp_input_A [0] <= _0010_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.tmp_input_A [1] <= 1'h0;
		else if (_0004_)
			\mchip.tmp_input_A [1] <= _0017_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.tmp_input_A [2] <= 1'h0;
		else if (_0004_)
			\mchip.tmp_input_A [2] <= _0018_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.tmp_input_A [3] <= 1'h0;
		else if (_0004_)
			\mchip.tmp_input_A [3] <= _0019_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.tmp_input_A [4] <= 1'h0;
		else if (_0004_)
			\mchip.tmp_input_A [4] <= _0020_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.tmp_input_A [5] <= 1'h0;
		else if (_0004_)
			\mchip.tmp_input_A [5] <= _0021_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.tmp_input_A [6] <= 1'h0;
		else if (_0004_)
			\mchip.tmp_input_A [6] <= _0022_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.tmp_input_A [7] <= 1'h0;
		else if (_0004_)
			\mchip.tmp_input_A [7] <= _0023_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.tmp_input_A [8] <= 1'h0;
		else if (_0004_)
			\mchip.tmp_input_A [8] <= _0024_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.tmp_input_A [9] <= 1'h0;
		else if (_0004_)
			\mchip.tmp_input_A [9] <= _0025_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.tmp_input_A [10] <= 1'h0;
		else if (_0004_)
			\mchip.tmp_input_A [10] <= _0011_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.tmp_input_A [11] <= 1'h0;
		else if (_0004_)
			\mchip.tmp_input_A [11] <= _0012_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.tmp_input_A [12] <= 1'h0;
		else if (_0004_)
			\mchip.tmp_input_A [12] <= _0013_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.tmp_input_A [13] <= 1'h0;
		else if (_0004_)
			\mchip.tmp_input_A [13] <= _0014_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.tmp_input_A [14] <= 1'h0;
		else if (_0004_)
			\mchip.tmp_input_A [14] <= _0015_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.tmp_input_A [15] <= 1'h0;
		else if (_0004_)
			\mchip.tmp_input_A [15] <= _0016_;
	always @(posedge io_in[12])
		if (_0007_)
			\mchip.value_A [0] <= \mchip.tmp_input_A [0];
	always @(posedge io_in[12])
		if (_0007_)
			\mchip.value_A [1] <= \mchip.tmp_input_A [1];
	always @(posedge io_in[12])
		if (_0007_)
			\mchip.value_A [2] <= \mchip.tmp_input_A [2];
	always @(posedge io_in[12])
		if (_0007_)
			\mchip.value_A [3] <= \mchip.tmp_input_A [3];
	always @(posedge io_in[12])
		if (_0007_)
			\mchip.value_A [4] <= \mchip.tmp_input_A [4];
	always @(posedge io_in[12])
		if (_0007_)
			\mchip.value_A [5] <= \mchip.tmp_input_A [5];
	always @(posedge io_in[12])
		if (_0007_)
			\mchip.value_A [6] <= \mchip.tmp_input_A [6];
	always @(posedge io_in[12])
		if (_0007_)
			\mchip.value_A [7] <= \mchip.tmp_input_A [7];
	always @(posedge io_in[12])
		if (_0007_)
			\mchip.value_A [8] <= \mchip.tmp_input_A [8];
	always @(posedge io_in[12])
		if (_0007_)
			\mchip.value_A [9] <= \mchip.tmp_input_A [9];
	always @(posedge io_in[12])
		if (_0007_)
			\mchip.value_A [10] <= \mchip.tmp_input_A [10];
	always @(posedge io_in[12])
		if (_0007_)
			\mchip.value_A [11] <= \mchip.tmp_input_A [11];
	always @(posedge io_in[12])
		if (_0007_)
			\mchip.value_A [12] <= \mchip.tmp_input_A [12];
	always @(posedge io_in[12])
		if (_0007_)
			\mchip.value_A [13] <= \mchip.tmp_input_A [13];
	always @(posedge io_in[12])
		if (_0007_)
			\mchip.value_A [14] <= \mchip.tmp_input_A [14];
	always @(posedge io_in[12])
		if (_0007_)
			\mchip.value_A [15] <= \mchip.tmp_input_A [15];
	reg \mchip.io_out_reg[0] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.io_out_reg[0]  <= 1'h0;
		else if (_0008_)
			\mchip.io_out_reg[0]  <= _0043_;
	assign \mchip.io_out [0] = \mchip.io_out_reg[0] ;
	reg \mchip.io_out_reg[1] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.io_out_reg[1]  <= 1'h0;
		else if (_0008_)
			\mchip.io_out_reg[1]  <= _0044_;
	assign \mchip.io_out [1] = \mchip.io_out_reg[1] ;
	reg \mchip.io_out_reg[2] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.io_out_reg[2]  <= 1'h0;
		else if (_0008_)
			\mchip.io_out_reg[2]  <= _0045_;
	assign \mchip.io_out [2] = \mchip.io_out_reg[2] ;
	reg \mchip.io_out_reg[3] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.io_out_reg[3]  <= 1'h0;
		else if (_0008_)
			\mchip.io_out_reg[3]  <= _0046_;
	assign \mchip.io_out [3] = \mchip.io_out_reg[3] ;
	reg \mchip.io_out_reg[4] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.io_out_reg[4]  <= 1'h0;
		else if (_0008_)
			\mchip.io_out_reg[4]  <= _0047_;
	assign \mchip.io_out [4] = \mchip.io_out_reg[4] ;
	reg \mchip.io_out_reg[5] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.io_out_reg[5]  <= 1'h0;
		else if (_0008_)
			\mchip.io_out_reg[5]  <= _0048_;
	assign \mchip.io_out [5] = \mchip.io_out_reg[5] ;
	reg \mchip.io_out_reg[6] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.io_out_reg[6]  <= 1'h0;
		else if (_0008_)
			\mchip.io_out_reg[6]  <= _0049_;
	assign \mchip.io_out [6] = \mchip.io_out_reg[6] ;
	reg \mchip.io_out_reg[7] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.io_out_reg[7]  <= 1'h0;
		else if (_0008_)
			\mchip.io_out_reg[7]  <= _0050_;
	assign \mchip.io_out [7] = \mchip.io_out_reg[7] ;
	assign _3757_[3:1] = \mchip.count [3:1];
	assign _3758_[0] = _3757_[0];
	assign io_out = {5'h00, \mchip.io_out [8:0]};
	assign \mchip.clock  = io_in[12];
	assign \mchip.inst_add.add_valid  = \mchip.temp_valid_add ;
	assign \mchip.inst_add.input_a  = \mchip.value_A ;
	assign \mchip.inst_add.input_b  = \mchip.value_B ;
	assign \mchip.inst_add.temp_3  = 5'h00;
	assign \mchip.inst_mul.expo_1_temp  = \mchip.value_A [14:10];
	assign \mchip.inst_mul.expo_2_temp  = \mchip.value_B [14:10];
	assign \mchip.inst_mul.frac_1  = \mchip.value_A [9:0];
	assign \mchip.inst_mul.frac_2  = \mchip.value_B [9:0];
	assign \mchip.inst_mul.input_a  = \mchip.value_A ;
	assign \mchip.inst_mul.input_b  = \mchip.value_B ;
	assign \mchip.inst_mul.mul_valid  = \mchip.temp_valid_add ;
	assign \mchip.inst_mul.sign_1  = \mchip.value_A [15];
	assign \mchip.inst_mul.sign_2  = \mchip.value_B [15];
	assign \mchip.inst_mul.temp_f_1  = {1'h0, \mchip.value_A [9:0], 10'h000};
	assign \mchip.inst_mul.temp_f_2  = {1'h0, \mchip.value_B [9:0]};
	assign \mchip.inst_mul.temp_value[0]  = 21'h000000;
	assign \mchip.inst_mul.temp_value[10]  = 21'h000000;
	assign \mchip.inst_mul.temp_value[1]  = 21'h000000;
	assign \mchip.inst_mul.temp_value[2]  = 21'h000000;
	assign \mchip.inst_mul.temp_value[3]  = 21'h000000;
	assign \mchip.inst_mul.temp_value[4]  = 21'h000000;
	assign \mchip.inst_mul.temp_value[5]  = 21'h000000;
	assign \mchip.inst_mul.temp_value[6]  = 21'h000000;
	assign \mchip.inst_mul.temp_value[7]  = 21'h000000;
	assign \mchip.inst_mul.temp_value[8]  = 21'h000000;
	assign \mchip.inst_mul.temp_value[9]  = 21'h000000;
	assign \mchip.io_in  = io_in[11:0];
	assign \mchip.io_out [11:9] = 3'h0;
	assign {\mchip.j [31], \mchip.j [29:6], \mchip.j [0]} = {\mchip.j [30], \mchip.j [30], \mchip.j [30], \mchip.j [30], \mchip.j [30], \mchip.j [30], \mchip.j [30], \mchip.j [30], \mchip.j [30], \mchip.j [30], \mchip.j [30], \mchip.j [30], \mchip.j [30], \mchip.j [30], \mchip.j [30], \mchip.j [30], \mchip.j [30], \mchip.j [30], \mchip.j [30], \mchip.j [30], \mchip.j [30], \mchip.j [30], \mchip.j [30], \mchip.j [30], \mchip.j [30], \mchip.j [1]};
	assign \mchip.reset  = io_in[13];
	assign \mchip.select  = io_in[8];
	assign \mchip.temp_valid_mul  = \mchip.temp_valid_add ;
endmodule
module d28_gvenkata_ucpu (
	io_in,
	io_out
);
	wire [3:0] _0000_;
	wire [7:0] _0001_;
	wire _0002_;
	wire _0003_;
	wire _0004_;
	wire _0005_;
	wire _0006_;
	wire _0007_;
	wire _0008_;
	wire _0009_;
	wire _0010_;
	wire _0011_;
	wire _0012_;
	wire _0013_;
	wire _0014_;
	wire _0015_;
	wire _0016_;
	wire _0017_;
	wire _0018_;
	wire _0019_;
	wire _0020_;
	wire _0021_;
	wire _0022_;
	wire _0023_;
	wire _0024_;
	wire _0025_;
	wire _0026_;
	wire _0027_;
	wire _0028_;
	wire _0029_;
	wire _0030_;
	wire _0031_;
	wire _0032_;
	wire _0033_;
	wire _0034_;
	wire _0035_;
	wire _0036_;
	wire _0037_;
	wire _0038_;
	wire _0039_;
	wire _0040_;
	wire _0041_;
	wire _0042_;
	wire _0043_;
	wire _0044_;
	wire _0045_;
	wire _0046_;
	wire _0047_;
	wire _0048_;
	wire _0049_;
	wire _0050_;
	wire _0051_;
	wire _0052_;
	wire _0053_;
	wire _0054_;
	wire _0055_;
	wire _0056_;
	wire _0057_;
	wire _0058_;
	wire _0059_;
	wire _0060_;
	wire _0061_;
	wire _0062_;
	wire _0063_;
	wire _0064_;
	wire _0065_;
	wire _0066_;
	wire _0067_;
	wire _0068_;
	wire _0069_;
	wire _0070_;
	wire _0071_;
	wire _0072_;
	wire _0073_;
	wire _0074_;
	wire _0075_;
	wire _0076_;
	wire _0077_;
	wire _0078_;
	wire _0079_;
	wire _0080_;
	wire _0081_;
	wire _0082_;
	wire _0083_;
	wire _0084_;
	wire _0085_;
	wire _0086_;
	wire _0087_;
	wire _0088_;
	wire _0089_;
	wire _0090_;
	wire _0091_;
	wire _0092_;
	wire _0093_;
	wire _0094_;
	wire _0095_;
	wire _0096_;
	wire _0097_;
	wire _0098_;
	wire _0099_;
	wire _0100_;
	wire _0101_;
	wire _0102_;
	wire _0103_;
	wire _0104_;
	wire _0105_;
	wire _0106_;
	wire _0107_;
	wire _0108_;
	wire _0109_;
	wire _0110_;
	wire _0111_;
	wire _0112_;
	wire _0113_;
	wire _0114_;
	wire _0115_;
	wire _0116_;
	wire _0117_;
	wire _0118_;
	wire _0119_;
	wire _0120_;
	wire _0121_;
	wire _0122_;
	wire _0123_;
	wire _0124_;
	wire _0125_;
	wire _0126_;
	wire _0127_;
	wire _0128_;
	wire _0129_;
	wire _0130_;
	wire _0131_;
	wire _0132_;
	wire _0133_;
	wire _0134_;
	wire _0135_;
	wire _0136_;
	wire _0137_;
	wire _0138_;
	wire _0139_;
	wire _0140_;
	wire _0141_;
	wire _0142_;
	wire _0143_;
	wire _0144_;
	wire _0145_;
	wire _0146_;
	wire _0147_;
	wire _0148_;
	wire _0149_;
	wire _0150_;
	wire _0151_;
	wire _0152_;
	wire _0153_;
	wire _0154_;
	wire _0155_;
	wire _0156_;
	wire _0157_;
	wire _0158_;
	wire _0159_;
	wire _0160_;
	wire _0161_;
	wire _0162_;
	wire _0163_;
	wire _0164_;
	wire _0165_;
	wire _0166_;
	wire _0167_;
	wire _0168_;
	wire _0169_;
	wire _0170_;
	wire _0171_;
	wire _0172_;
	wire _0173_;
	wire _0174_;
	wire _0175_;
	wire _0176_;
	wire _0177_;
	wire _0178_;
	wire _0179_;
	wire _0180_;
	wire _0181_;
	wire _0182_;
	wire _0183_;
	wire _0184_;
	wire _0185_;
	wire _0186_;
	wire _0187_;
	wire _0188_;
	wire _0189_;
	wire _0190_;
	wire _0191_;
	wire _0192_;
	wire _0193_;
	wire _0194_;
	wire _0195_;
	wire _0196_;
	wire _0197_;
	wire _0198_;
	wire _0199_;
	wire _0200_;
	wire _0201_;
	wire _0202_;
	wire _0203_;
	wire _0204_;
	wire _0205_;
	wire _0206_;
	wire _0207_;
	wire _0208_;
	wire _0209_;
	wire _0210_;
	wire _0211_;
	wire _0212_;
	wire _0213_;
	wire _0214_;
	wire _0215_;
	wire _0216_;
	wire _0217_;
	wire _0218_;
	wire _0219_;
	wire _0220_;
	wire _0221_;
	wire _0222_;
	wire _0223_;
	wire _0224_;
	wire _0225_;
	wire _0226_;
	wire _0227_;
	wire _0228_;
	wire _0229_;
	wire _0230_;
	wire _0231_;
	wire _0232_;
	wire _0233_;
	wire _0234_;
	wire _0235_;
	wire _0236_;
	wire _0237_;
	wire _0238_;
	wire _0239_;
	wire _0240_;
	wire _0241_;
	wire _0242_;
	wire _0243_;
	wire _0244_;
	wire _0245_;
	wire _0246_;
	wire _0247_;
	wire _0248_;
	wire _0249_;
	wire _0250_;
	wire _0251_;
	wire _0252_;
	wire _0253_;
	wire _0254_;
	wire _0255_;
	wire _0256_;
	wire _0257_;
	wire _0258_;
	wire _0259_;
	wire _0260_;
	wire _0261_;
	wire _0262_;
	wire _0263_;
	wire _0264_;
	wire _0265_;
	wire _0266_;
	wire _0267_;
	wire _0268_;
	wire _0269_;
	wire _0270_;
	wire _0271_;
	wire _0272_;
	wire _0273_;
	wire _0274_;
	wire _0275_;
	wire _0276_;
	wire _0277_;
	wire _0278_;
	wire _0279_;
	wire _0280_;
	wire _0281_;
	wire _0282_;
	wire _0283_;
	wire _0284_;
	wire _0285_;
	wire _0286_;
	wire _0287_;
	wire _0288_;
	wire _0289_;
	wire _0290_;
	wire _0291_;
	wire _0292_;
	wire _0293_;
	wire _0294_;
	wire _0295_;
	wire _0296_;
	wire _0297_;
	wire _0298_;
	wire _0299_;
	wire _0300_;
	wire _0301_;
	wire _0302_;
	wire _0303_;
	wire _0304_;
	wire _0305_;
	wire _0306_;
	wire _0307_;
	wire _0308_;
	wire _0309_;
	wire _0310_;
	wire _0311_;
	wire _0312_;
	wire _0313_;
	wire _0314_;
	wire _0315_;
	wire _0316_;
	wire _0317_;
	wire _0318_;
	wire _0319_;
	wire _0320_;
	wire _0321_;
	wire _0322_;
	wire _0323_;
	wire _0324_;
	wire _0325_;
	wire _0326_;
	wire _0327_;
	wire _0328_;
	wire _0329_;
	wire _0330_;
	wire _0331_;
	wire _0332_;
	wire _0333_;
	wire _0334_;
	wire _0335_;
	wire _0336_;
	wire _0337_;
	wire _0338_;
	wire _0339_;
	wire _0340_;
	wire _0341_;
	wire _0342_;
	wire _0343_;
	wire _0344_;
	wire _0345_;
	wire _0346_;
	wire _0347_;
	wire _0348_;
	wire _0349_;
	wire _0350_;
	wire _0351_;
	wire _0352_;
	wire _0353_;
	wire _0354_;
	wire _0355_;
	wire _0356_;
	wire _0357_;
	wire _0358_;
	wire _0359_;
	wire _0360_;
	wire _0361_;
	wire _0362_;
	wire _0363_;
	wire _0364_;
	wire _0365_;
	wire _0366_;
	wire _0367_;
	wire _0368_;
	wire _0369_;
	wire _0370_;
	wire _0371_;
	wire _0372_;
	wire _0373_;
	wire _0374_;
	wire _0375_;
	wire _0376_;
	wire _0377_;
	wire _0378_;
	wire _0379_;
	wire _0380_;
	wire _0381_;
	wire _0382_;
	wire _0383_;
	wire _0384_;
	wire _0385_;
	wire _0386_;
	wire _0387_;
	wire _0388_;
	wire _0389_;
	wire _0390_;
	wire _0391_;
	wire _0392_;
	wire _0393_;
	wire _0394_;
	wire _0395_;
	wire _0396_;
	wire _0397_;
	wire _0398_;
	wire _0399_;
	wire _0400_;
	wire _0401_;
	wire _0402_;
	wire _0403_;
	wire _0404_;
	wire _0405_;
	wire _0406_;
	wire _0407_;
	wire _0408_;
	wire _0409_;
	wire _0410_;
	wire _0411_;
	wire _0412_;
	wire _0413_;
	wire _0414_;
	wire _0415_;
	wire _0416_;
	wire _0417_;
	wire _0418_;
	wire _0419_;
	wire _0420_;
	wire _0421_;
	wire _0422_;
	wire _0423_;
	wire _0424_;
	wire _0425_;
	wire _0426_;
	wire _0427_;
	wire _0428_;
	wire _0429_;
	wire _0430_;
	wire _0431_;
	wire _0432_;
	wire _0433_;
	wire _0434_;
	wire _0435_;
	wire _0436_;
	wire _0437_;
	wire _0438_;
	wire _0439_;
	wire _0440_;
	wire _0441_;
	wire _0442_;
	wire _0443_;
	wire _0444_;
	wire _0445_;
	wire _0446_;
	wire _0447_;
	wire _0448_;
	wire _0449_;
	wire _0450_;
	wire _0451_;
	wire _0452_;
	wire _0453_;
	wire _0454_;
	wire _0455_;
	wire _0456_;
	wire _0457_;
	wire _0458_;
	wire _0459_;
	wire _0460_;
	wire _0461_;
	wire _0462_;
	wire _0463_;
	wire _0464_;
	wire _0465_;
	wire _0466_;
	wire _0467_;
	wire _0468_;
	wire _0469_;
	wire _0470_;
	wire _0471_;
	wire _0472_;
	wire _0473_;
	wire _0474_;
	wire _0475_;
	wire _0476_;
	wire _0477_;
	wire _0478_;
	wire _0479_;
	wire _0480_;
	wire _0481_;
	wire _0482_;
	wire _0483_;
	wire _0484_;
	wire _0485_;
	wire _0486_;
	wire _0487_;
	wire _0488_;
	wire _0489_;
	wire _0490_;
	wire _0491_;
	wire _0492_;
	wire _0493_;
	wire _0494_;
	wire _0495_;
	wire _0496_;
	wire _0497_;
	wire _0498_;
	wire _0499_;
	wire _0500_;
	wire _0501_;
	wire _0502_;
	wire _0503_;
	wire _0504_;
	wire _0505_;
	wire _0506_;
	wire _0507_;
	wire _0508_;
	wire _0509_;
	wire _0510_;
	wire _0511_;
	wire _0512_;
	wire _0513_;
	wire _0514_;
	wire _0515_;
	wire _0516_;
	wire _0517_;
	wire _0518_;
	wire _0519_;
	wire _0520_;
	wire _0521_;
	wire _0522_;
	wire _0523_;
	wire _0524_;
	wire _0525_;
	wire _0526_;
	wire _0527_;
	wire _0528_;
	wire _0529_;
	wire _0530_;
	wire _0531_;
	wire _0532_;
	wire _0533_;
	wire _0534_;
	wire _0535_;
	wire _0536_;
	wire _0537_;
	wire _0538_;
	wire _0539_;
	wire _0540_;
	wire _0541_;
	wire _0542_;
	wire _0543_;
	wire _0544_;
	wire _0545_;
	wire _0546_;
	wire _0547_;
	wire _0548_;
	wire _0549_;
	wire _0550_;
	wire _0551_;
	wire _0552_;
	wire _0553_;
	wire _0554_;
	wire _0555_;
	wire _0556_;
	wire _0557_;
	wire _0558_;
	wire _0559_;
	wire _0560_;
	wire _0561_;
	wire _0562_;
	wire _0563_;
	wire _0564_;
	wire _0565_;
	wire _0566_;
	wire _0567_;
	wire _0568_;
	wire _0569_;
	wire _0570_;
	wire _0571_;
	wire _0572_;
	wire _0573_;
	wire _0574_;
	wire _0575_;
	wire _0576_;
	wire _0577_;
	wire _0578_;
	wire _0579_;
	wire _0580_;
	wire _0581_;
	wire _0582_;
	wire _0583_;
	wire _0584_;
	wire _0585_;
	wire _0586_;
	wire _0587_;
	wire _0588_;
	wire _0589_;
	wire _0590_;
	wire _0591_;
	wire _0592_;
	wire _0593_;
	wire _0594_;
	wire _0595_;
	wire _0596_;
	wire _0597_;
	wire _0598_;
	wire _0599_;
	wire _0600_;
	wire _0601_;
	wire _0602_;
	wire _0603_;
	wire _0604_;
	wire _0605_;
	wire _0606_;
	wire _0607_;
	wire _0608_;
	wire _0609_;
	wire _0610_;
	wire _0611_;
	wire _0612_;
	wire _0613_;
	wire _0614_;
	wire _0615_;
	wire _0616_;
	wire _0617_;
	wire _0618_;
	wire _0619_;
	wire _0620_;
	wire _0621_;
	wire _0622_;
	wire _0623_;
	wire _0624_;
	wire _0625_;
	wire _0626_;
	wire _0627_;
	wire _0628_;
	wire _0629_;
	wire _0630_;
	wire _0631_;
	wire _0632_;
	wire _0633_;
	wire _0634_;
	wire _0635_;
	wire _0636_;
	wire _0637_;
	wire _0638_;
	wire _0639_;
	wire _0640_;
	wire _0641_;
	wire _0642_;
	wire _0643_;
	wire _0644_;
	wire _0645_;
	wire _0646_;
	wire _0647_;
	wire _0648_;
	wire _0649_;
	wire _0650_;
	wire _0651_;
	wire _0652_;
	wire _0653_;
	wire _0654_;
	wire _0655_;
	wire _0656_;
	wire _0657_;
	wire _0658_;
	wire _0659_;
	wire _0660_;
	wire _0661_;
	wire _0662_;
	wire _0663_;
	wire _0664_;
	wire _0665_;
	wire _0666_;
	wire _0667_;
	wire _0668_;
	wire _0669_;
	wire _0670_;
	wire _0671_;
	wire _0672_;
	wire _0673_;
	wire _0674_;
	wire _0675_;
	wire _0676_;
	wire _0677_;
	wire _0678_;
	wire _0679_;
	wire _0680_;
	wire _0681_;
	wire _0682_;
	wire _0683_;
	wire _0684_;
	wire _0685_;
	wire _0686_;
	wire _0687_;
	wire _0688_;
	wire _0689_;
	wire _0690_;
	wire _0691_;
	wire _0692_;
	wire _0693_;
	wire _0694_;
	wire _0695_;
	wire _0696_;
	wire _0697_;
	wire _0698_;
	wire _0699_;
	wire _0700_;
	wire _0701_;
	wire _0702_;
	wire _0703_;
	wire _0704_;
	wire _0705_;
	wire _0706_;
	wire _0707_;
	wire _0708_;
	wire _0709_;
	wire _0710_;
	wire _0711_;
	wire _0712_;
	wire _0713_;
	wire _0714_;
	wire _0715_;
	wire _0716_;
	wire _0717_;
	wire _0718_;
	wire _0719_;
	wire _0720_;
	wire _0721_;
	wire _0722_;
	wire _0723_;
	wire _0724_;
	wire _0725_;
	wire _0726_;
	wire _0727_;
	wire _0728_;
	wire _0729_;
	wire _0730_;
	wire _0731_;
	wire _0732_;
	wire _0733_;
	wire _0734_;
	wire _0735_;
	wire _0736_;
	wire _0737_;
	wire _0738_;
	wire _0739_;
	wire _0740_;
	wire _0741_;
	wire _0742_;
	wire _0743_;
	wire _0744_;
	wire _0745_;
	wire _0746_;
	wire _0747_;
	wire _0748_;
	wire [3:0] _0749_;
	input wire [13:0] io_in;
	output wire [13:0] io_out;
	wire \mchip.clock ;
	wire [11:0] \mchip.io_in ;
	wire [11:0] \mchip.io_out ;
	wire [7:0] \mchip.micro_coded_cpu.A_reg ;
	wire \mchip.micro_coded_cpu.B_Reg ;
	wire [7:0] \mchip.micro_coded_cpu.B_reg ;
	wire \mchip.micro_coded_cpu.alu_en_A ;
	wire \mchip.micro_coded_cpu.alu_en_A_md ;
	wire \mchip.micro_coded_cpu.alu_en_B ;
	wire \mchip.micro_coded_cpu.alu_en_B_md ;
	wire [2:0] \mchip.micro_coded_cpu.alu_op ;
	wire [2:0] \mchip.micro_coded_cpu.alu_op_md ;
	wire [7:0] \mchip.micro_coded_cpu.alu_result ;
	wire [7:0] \mchip.micro_coded_cpu.alu_top.A_bus ;
	reg [7:0] \mchip.micro_coded_cpu.alu_top.A_reg ;
	wire [7:0] \mchip.micro_coded_cpu.alu_top.B_bus ;
	reg [7:0] \mchip.micro_coded_cpu.alu_top.B_reg ;
	wire [7:0] \mchip.micro_coded_cpu.alu_top.alu.A ;
	wire [7:0] \mchip.micro_coded_cpu.alu_top.alu.B ;
	wire \mchip.micro_coded_cpu.alu_top.alu.a_equal_b ;
	wire \mchip.micro_coded_cpu.alu_top.alu.a_greater_b ;
	wire [2:0] \mchip.micro_coded_cpu.alu_top.alu.alu_op ;
	wire [7:0] \mchip.micro_coded_cpu.alu_top.alu.alu_result ;
	wire [7:0] \mchip.micro_coded_cpu.alu_top.alu.alu_result_tmp ;
	wire \mchip.micro_coded_cpu.alu_top.alu.carry_in ;
	wire \mchip.micro_coded_cpu.alu_top.alu.equal ;
	wire \mchip.micro_coded_cpu.alu_top.alu.greater ;
	wire [7:0] \mchip.micro_coded_cpu.alu_top.alu.zero ;
	wire \mchip.micro_coded_cpu.alu_top.alu_en_A_reg ;
	wire \mchip.micro_coded_cpu.alu_top.alu_en_B_reg ;
	wire [2:0] \mchip.micro_coded_cpu.alu_top.alu_op ;
	reg [7:0] \mchip.micro_coded_cpu.alu_top.alu_result ;
	wire [7:0] \mchip.micro_coded_cpu.alu_top.alu_result_out ;
	wire \mchip.micro_coded_cpu.alu_top.carry_in ;
	wire \mchip.micro_coded_cpu.alu_top.cc_equal ;
	wire \mchip.micro_coded_cpu.alu_top.cc_equal_out ;
	wire \mchip.micro_coded_cpu.alu_top.cc_greater ;
	wire \mchip.micro_coded_cpu.alu_top.cc_greater_out ;
	wire [3:0] \mchip.micro_coded_cpu.alu_top.cpu_state ;
	wire \mchip.micro_coded_cpu.alu_top.sys_clk ;
	wire \mchip.micro_coded_cpu.alu_top.sys_reset ;
	wire [7:0] \mchip.micro_coded_cpu.branch_target_id ;
	wire \mchip.micro_coded_cpu.cc_equal ;
	wire \mchip.micro_coded_cpu.cc_greater ;
	wire [3:0] \mchip.micro_coded_cpu.cpu_fsm_top.cpu_state ;
	reg [4:0] \mchip.micro_coded_cpu.cpu_fsm_top.current_minst_1 ;
	reg [5:0] \mchip.micro_coded_cpu.cpu_fsm_top.fsm_assist ;
	wire \mchip.micro_coded_cpu.cpu_fsm_top.is_micro_nop ;
	wire \mchip.micro_coded_cpu.cpu_fsm_top.is_nop ;
	wire \mchip.micro_coded_cpu.cpu_fsm_top.sys_clk ;
	wire \mchip.micro_coded_cpu.cpu_fsm_top.sys_reset ;
	wire [3:0] \mchip.micro_coded_cpu.cpu_state ;
	wire [7:0] \mchip.micro_coded_cpu.imm ;
	wire [7:0] \mchip.micro_coded_cpu.imm_id ;
	wire [7:0] \mchip.micro_coded_cpu.imm_md ;
	wire \mchip.micro_coded_cpu.inst_addr_stream ;
	wire [3:0] \mchip.micro_coded_cpu.inst_to_bit.cpu_state ;
	wire [7:0] \mchip.micro_coded_cpu.inst_to_bit.inst_addr ;
	wire \mchip.micro_coded_cpu.inst_to_bit.inst_addr_stream ;
	wire \mchip.micro_coded_cpu.inst_to_bit.sys_clk ;
	wire \mchip.micro_coded_cpu.inst_to_bit.sys_reset ;
	wire [4:0] \mchip.micro_coded_cpu.inst_type ;
	wire \mchip.micro_coded_cpu.instr_in ;
	wire [31:0] \mchip.micro_coded_cpu.instr_reg ;
	wire \mchip.micro_coded_cpu.instr_reg_top.instr_in ;
	reg [31:0] \mchip.micro_coded_cpu.instr_reg_top.instr_reg ;
	wire \mchip.micro_coded_cpu.instr_reg_top.sys_clk ;
	wire \mchip.micro_coded_cpu.instr_reg_top.sys_reset ;
	wire [7:0] \mchip.micro_coded_cpu.ir_decode_top.branch_target_id ;
	wire [7:0] \mchip.micro_coded_cpu.ir_decode_top.imm_id ;
	wire [4:0] \mchip.micro_coded_cpu.ir_decode_top.inst_type ;
	wire [31:0] \mchip.micro_coded_cpu.ir_decode_top.instr_in ;
	wire \mchip.micro_coded_cpu.ir_decode_top.is_imm_active_id ;
	wire [3:0] \mchip.micro_coded_cpu.ir_decode_top.reg_dst_id ;
	wire [3:0] \mchip.micro_coded_cpu.ir_decode_top.reg_src_1_id ;
	wire [3:0] \mchip.micro_coded_cpu.ir_decode_top.reg_src_2_id ;
	wire \mchip.micro_coded_cpu.is_current_inst_nop ;
	wire \mchip.micro_coded_cpu.is_current_micro_inst_nop ;
	wire \mchip.micro_coded_cpu.is_imm_active ;
	wire \mchip.micro_coded_cpu.is_imm_active_id ;
	wire \mchip.micro_coded_cpu.is_imm_active_md ;
	wire \mchip.micro_coded_cpu.load_m_pc_en ;
	wire \mchip.micro_coded_cpu.load_pc_en ;
	wire [8:0] \mchip.micro_coded_cpu.m_inst_addr_offset ;
	wire [31:0] \mchip.micro_coded_cpu.m_inst_addr_offset_gen.instr_in ;
	wire [4:0] \mchip.micro_coded_cpu.m_inst_addr_offset_gen.instr_type ;
	wire [8:0] \mchip.micro_coded_cpu.m_inst_addr_offset_gen.m_inst_addr_base ;
	wire [8:0] \mchip.micro_coded_cpu.m_inst_addr_offset_gen.offset ;
	wire \mchip.micro_coded_cpu.m_inst_addr_stream ;
	wire \mchip.micro_coded_cpu.m_inst_decode_top.alu_en_A_md ;
	wire \mchip.micro_coded_cpu.m_inst_decode_top.alu_en_B_md ;
	wire [2:0] \mchip.micro_coded_cpu.m_inst_decode_top.alu_op_md ;
	wire [7:0] \mchip.micro_coded_cpu.m_inst_decode_top.imm_md ;
	wire \mchip.micro_coded_cpu.m_inst_decode_top.is_imm_active_md ;
	wire [9:0] \mchip.micro_coded_cpu.m_inst_decode_top.m_args ;
	wire [7:0] \mchip.micro_coded_cpu.m_inst_decode_top.mbranch_target_md ;
	wire [43:0] \mchip.micro_coded_cpu.m_inst_decode_top.minstr_in ;
	wire [2:0] \mchip.micro_coded_cpu.m_inst_decode_top.minstr_type ;
	wire [4:0] \mchip.micro_coded_cpu.m_inst_decode_top.reg_dst_md ;
	wire \mchip.micro_coded_cpu.m_inst_decode_top.reg_file_en_md ;
	wire \mchip.micro_coded_cpu.m_inst_decode_top.reg_file_rw_md ;
	wire [4:0] \mchip.micro_coded_cpu.m_inst_decode_top.reg_src_md ;
	wire [3:0] \mchip.micro_coded_cpu.m_inst_to_bit.cpu_state ;
	reg [3:0] \mchip.micro_coded_cpu.m_inst_to_bit.current_bit_index ;
	wire [8:0] \mchip.micro_coded_cpu.m_inst_to_bit.m_inst_addr ;
	wire \mchip.micro_coded_cpu.m_inst_to_bit.m_inst_addr_stream ;
	wire \mchip.micro_coded_cpu.m_inst_to_bit.sys_clk ;
	wire \mchip.micro_coded_cpu.m_inst_to_bit.sys_reset ;
	wire \mchip.micro_coded_cpu.m_instr_in ;
	wire [43:0] \mchip.micro_coded_cpu.m_instr_reg ;
	reg [43:0] \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg ;
	wire \mchip.micro_coded_cpu.m_instr_reg_top.minstr_in ;
	wire \mchip.micro_coded_cpu.m_instr_reg_top.sys_clk ;
	wire \mchip.micro_coded_cpu.m_instr_reg_top.sys_reset ;
	wire [7:0] \mchip.micro_coded_cpu.m_pc ;
	wire \mchip.micro_coded_cpu.m_pc_top.load_m_pc_en ;
	reg [7:0] \mchip.micro_coded_cpu.m_pc_top.m_pc ;
	wire [7:0] \mchip.micro_coded_cpu.m_pc_top.next_m_pc ;
	wire \mchip.micro_coded_cpu.m_pc_top.sys_clk ;
	wire \mchip.micro_coded_cpu.m_pc_top.sys_reset ;
	wire [7:0] \mchip.micro_coded_cpu.mbranch_target ;
	wire [7:0] \mchip.micro_coded_cpu.mbranch_target_md ;
	reg \mchip.micro_coded_cpu.mdecode_reg_top.alu_en_A ;
	wire \mchip.micro_coded_cpu.mdecode_reg_top.alu_en_A_md ;
	reg \mchip.micro_coded_cpu.mdecode_reg_top.alu_en_B ;
	wire \mchip.micro_coded_cpu.mdecode_reg_top.alu_en_B_md ;
	reg [2:0] \mchip.micro_coded_cpu.mdecode_reg_top.alu_op ;
	wire [2:0] \mchip.micro_coded_cpu.mdecode_reg_top.alu_op_md ;
	reg [7:0] \mchip.micro_coded_cpu.mdecode_reg_top.imm ;
	wire [7:0] \mchip.micro_coded_cpu.mdecode_reg_top.imm_md ;
	reg \mchip.micro_coded_cpu.mdecode_reg_top.is_imm_active ;
	wire \mchip.micro_coded_cpu.mdecode_reg_top.is_imm_active_md ;
	reg [7:0] \mchip.micro_coded_cpu.mdecode_reg_top.mbranch_target ;
	wire [7:0] \mchip.micro_coded_cpu.mdecode_reg_top.mbranch_target_md ;
	reg [4:0] \mchip.micro_coded_cpu.mdecode_reg_top.reg_dst ;
	wire [4:0] \mchip.micro_coded_cpu.mdecode_reg_top.reg_dst_md ;
	reg \mchip.micro_coded_cpu.mdecode_reg_top.reg_file_en ;
	wire \mchip.micro_coded_cpu.mdecode_reg_top.reg_file_en_md ;
	reg \mchip.micro_coded_cpu.mdecode_reg_top.reg_file_rw ;
	wire \mchip.micro_coded_cpu.mdecode_reg_top.reg_file_rw_md ;
	reg [4:0] \mchip.micro_coded_cpu.mdecode_reg_top.reg_src ;
	wire [4:0] \mchip.micro_coded_cpu.mdecode_reg_top.reg_src_md ;
	wire \mchip.micro_coded_cpu.mdecode_reg_top.sys_clk ;
	wire \mchip.micro_coded_cpu.mdecode_reg_top.sys_reset ;
	wire [2:0] \mchip.micro_coded_cpu.minstr_type ;
	wire [8:0] \mchip.micro_coded_cpu.mpc_offset ;
	wire [7:0] \mchip.micro_coded_cpu.next_m_pc ;
	wire [7:0] \mchip.micro_coded_cpu.pc ;
	wire \mchip.micro_coded_cpu.pc_top.load_pc_en ;
	wire [7:0] \mchip.micro_coded_cpu.pc_top.pc ;
	wire \mchip.micro_coded_cpu.pc_top.sys_clk ;
	wire \mchip.micro_coded_cpu.pc_top.sys_reset ;
	wire [4:0] \mchip.micro_coded_cpu.reg_dst ;
	wire [3:0] \mchip.micro_coded_cpu.reg_dst_id ;
	wire [4:0] \mchip.micro_coded_cpu.reg_dst_md ;
	wire \mchip.micro_coded_cpu.reg_file_en ;
	wire \mchip.micro_coded_cpu.reg_file_en_md ;
	wire [3:0] \mchip.micro_coded_cpu.reg_file_interface.cpu_state ;
	reg [7:0] \mchip.micro_coded_cpu.reg_file_interface.mreg_file[0] ;
	reg [7:0] \mchip.micro_coded_cpu.reg_file_interface.mreg_file[1] ;
	reg [7:0] \mchip.micro_coded_cpu.reg_file_interface.mreg_file[2] ;
	reg [7:0] \mchip.micro_coded_cpu.reg_file_interface.mreg_file[3] ;
	wire [3:0] \mchip.micro_coded_cpu.reg_file_interface.reg_dst ;
	wire \mchip.micro_coded_cpu.reg_file_interface.reg_file_en ;
	wire \mchip.micro_coded_cpu.reg_file_interface.reg_file_rw ;
	wire [7:0] \mchip.micro_coded_cpu.reg_file_interface.reg_rd_data ;
	reg [7:0] \mchip.micro_coded_cpu.reg_file_interface.reg_rd_data_out ;
	reg [1:0] \mchip.micro_coded_cpu.reg_file_interface.reg_sel_in ;
	reg [7:0] \mchip.micro_coded_cpu.reg_file_interface.reg_wr_data_in ;
	wire [7:0] \mchip.micro_coded_cpu.reg_file_interface.shared_write_bus ;
	wire \mchip.micro_coded_cpu.reg_file_interface.sys_clk ;
	wire \mchip.micro_coded_cpu.reg_file_interface.sys_reset ;
	wire \mchip.micro_coded_cpu.reg_file_rw ;
	wire \mchip.micro_coded_cpu.reg_file_rw_md ;
	wire [7:0] \mchip.micro_coded_cpu.reg_rd_data ;
	wire [4:0] \mchip.micro_coded_cpu.reg_src ;
	wire [3:0] \mchip.micro_coded_cpu.reg_src_1_id ;
	wire [3:0] \mchip.micro_coded_cpu.reg_src_2_id ;
	wire [7:0] \mchip.micro_coded_cpu.reg_src_dst_cmp_branch.A ;
	wire [7:0] \mchip.micro_coded_cpu.reg_src_dst_cmp_branch.B ;
	wire [7:0] \mchip.micro_coded_cpu.reg_src_dst_cmp_branch.alu_result ;
	wire \mchip.micro_coded_cpu.reg_src_dst_cmp_branch.cc_equal ;
	wire \mchip.micro_coded_cpu.reg_src_dst_cmp_branch.cc_greater ;
	wire [7:0] \mchip.micro_coded_cpu.reg_src_dst_cmp_branch.imm ;
	wire \mchip.micro_coded_cpu.reg_src_dst_cmp_branch.is_imm_active ;
	wire [4:0] \mchip.micro_coded_cpu.reg_src_dst_cmp_branch.reg_dst ;
	wire [4:0] \mchip.micro_coded_cpu.reg_src_md ;
	wire [7:0] \mchip.micro_coded_cpu.shared_mcpu_bus.alu_result ;
	wire \mchip.micro_coded_cpu.shared_mcpu_bus.cc_equal ;
	wire \mchip.micro_coded_cpu.shared_mcpu_bus.cc_greater ;
	wire [7:0] \mchip.micro_coded_cpu.shared_mcpu_bus.imm ;
	wire [7:0] \mchip.micro_coded_cpu.shared_mcpu_bus.m_pc ;
	wire [7:0] \mchip.micro_coded_cpu.shared_mcpu_bus.mbranch_target ;
	wire [2:0] \mchip.micro_coded_cpu.shared_mcpu_bus.minstr_type ;
	wire [4:0] \mchip.micro_coded_cpu.shared_mcpu_bus.reg_dst ;
	wire [7:0] \mchip.micro_coded_cpu.shared_mcpu_bus.reg_rd_data ;
	wire [4:0] \mchip.micro_coded_cpu.shared_mcpu_bus.reg_src ;
	wire [1:0] \mchip.micro_coded_cpu.shared_mcpu_bus.rs1 ;
	wire [1:0] \mchip.micro_coded_cpu.shared_mcpu_bus.rs2 ;
	wire [7:0] \mchip.micro_coded_cpu.shared_mcpu_bus.write_bus_out ;
	wire [7:0] \mchip.micro_coded_cpu.shared_write_bus ;
	wire \mchip.micro_coded_cpu.sys_clk ;
	wire \mchip.micro_coded_cpu.sys_reset ;
	wire \mchip.reset ;
	assign _0749_[0] = ~\mchip.micro_coded_cpu.m_inst_to_bit.current_bit_index [0];
	assign _0041_ = ~\mchip.micro_coded_cpu.cpu_fsm_top.cpu_state [2];
	assign _0042_ = \mchip.micro_coded_cpu.cpu_fsm_top.cpu_state [0] & \mchip.micro_coded_cpu.cpu_fsm_top.cpu_state [1];
	assign _0043_ = _0042_ & ~_0041_;
	assign _0044_ = _0043_ & ~\mchip.micro_coded_cpu.mdecode_reg_top.reg_file_rw ;
	assign _0045_ = ~\mchip.micro_coded_cpu.mdecode_reg_top.reg_file_en ;
	assign _0046_ = \mchip.micro_coded_cpu.cpu_fsm_top.cpu_state [1] & ~\mchip.micro_coded_cpu.cpu_fsm_top.cpu_state [0];
	assign _0047_ = _0046_ & ~_0041_;
	assign _0048_ = _0047_ | _0045_;
	assign _0003_ = _0044_ & ~_0048_;
	assign _0049_ = ~io_in[13];
	assign _0050_ = _0042_ & ~\mchip.micro_coded_cpu.cpu_fsm_top.cpu_state [2];
	assign _0008_ = ~(_0050_ & _0049_);
	assign _0051_ = \mchip.micro_coded_cpu.instr_reg_top.instr_reg [25] | ~\mchip.micro_coded_cpu.instr_reg_top.instr_reg [24];
	assign _0052_ = \mchip.micro_coded_cpu.instr_reg_top.instr_reg [23] | ~\mchip.micro_coded_cpu.instr_reg_top.instr_reg [22];
	assign _0053_ = ~(_0052_ | _0051_);
	assign _0054_ = ~(_0053_ & _0047_);
	assign _0005_ = \mchip.micro_coded_cpu.mdecode_reg_top.reg_file_en  & ~_0054_;
	assign _0055_ = \mchip.micro_coded_cpu.cpu_fsm_top.cpu_state [0] & ~\mchip.micro_coded_cpu.cpu_fsm_top.cpu_state [1];
	assign _0030_ = _0055_ & ~\mchip.micro_coded_cpu.cpu_fsm_top.cpu_state [2];
	assign _0056_ = ~(\mchip.micro_coded_cpu.cpu_fsm_top.cpu_state [0] | \mchip.micro_coded_cpu.cpu_fsm_top.cpu_state [1]);
	assign _0031_ = _0056_ & ~_0041_;
	assign _0057_ = ~_0030_;
	assign _0058_ = \mchip.micro_coded_cpu.cpu_fsm_top.fsm_assist [0] & \mchip.micro_coded_cpu.cpu_fsm_top.fsm_assist [1];
	assign _0059_ = ~(\mchip.micro_coded_cpu.cpu_fsm_top.fsm_assist [2] & \mchip.micro_coded_cpu.cpu_fsm_top.fsm_assist [3]);
	assign _0060_ = _0058_ & ~_0059_;
	assign _0061_ = \mchip.micro_coded_cpu.cpu_fsm_top.fsm_assist [5] | ~\mchip.micro_coded_cpu.cpu_fsm_top.fsm_assist [4];
	assign _0062_ = _0060_ & ~_0061_;
	assign _0063_ = _0062_ | _0057_;
	assign _0064_ = _0056_ & ~\mchip.micro_coded_cpu.cpu_fsm_top.cpu_state [2];
	assign _0065_ = ~_0064_;
	assign _0066_ = ~(\mchip.micro_coded_cpu.cpu_fsm_top.fsm_assist [5] | \mchip.micro_coded_cpu.cpu_fsm_top.fsm_assist [4]);
	assign _0067_ = \mchip.micro_coded_cpu.cpu_fsm_top.fsm_assist [2] & ~\mchip.micro_coded_cpu.cpu_fsm_top.fsm_assist [3];
	assign _0068_ = ~(_0067_ & _0058_);
	assign _0069_ = _0066_ & ~_0068_;
	assign _0070_ = (_0064_ ? _0069_ : _0063_);
	assign _0071_ = _0046_ & ~\mchip.micro_coded_cpu.cpu_fsm_top.cpu_state [2];
	assign _0072_ = ~(_0071_ | _0030_);
	assign _0073_ = \mchip.micro_coded_cpu.cpu_fsm_top.fsm_assist [2] | ~\mchip.micro_coded_cpu.cpu_fsm_top.fsm_assist [3];
	assign _0074_ = _0058_ & ~_0073_;
	assign _0075_ = \mchip.micro_coded_cpu.cpu_fsm_top.fsm_assist [4] | ~\mchip.micro_coded_cpu.cpu_fsm_top.fsm_assist [5];
	assign _0076_ = _0074_ & ~_0075_;
	assign _0077_ = _0076_ | ~_0031_;
	assign _0078_ = _0072_ & ~_0077_;
	assign _0079_ = _0064_ | _0050_;
	assign _0080_ = _0078_ & ~_0079_;
	assign _0081_ = ~_0050_;
	assign _0082_ = \mchip.micro_coded_cpu.cpu_fsm_top.fsm_assist [0] | \mchip.micro_coded_cpu.cpu_fsm_top.fsm_assist [1];
	assign _0083_ = _0082_ | _0073_;
	assign _0084_ = _0066_ & ~_0083_;
	assign _0085_ = ~(_0084_ | _0081_);
	assign _0086_ = ~(_0085_ & _0072_);
	assign _0087_ = _0065_ & ~_0086_;
	assign _0088_ = _0087_ | _0080_;
	assign _0089_ = _0070_ & ~_0088_;
	assign _0090_ = _0031_ | _0047_;
	assign _0091_ = _0072_ & ~_0090_;
	assign _0092_ = (\mchip.micro_coded_cpu.cpu_fsm_top.cpu_state [2] ? _0042_ : _0056_);
	assign _0093_ = (\mchip.micro_coded_cpu.cpu_fsm_top.cpu_state [2] ? _0055_ : _0042_);
	assign _0094_ = _0093_ | _0092_;
	assign _0095_ = _0091_ & ~_0094_;
	assign _0007_ = _0089_ & ~_0095_;
	assign _0096_ = (\mchip.micro_coded_cpu.cpu_fsm_top.cpu_state [2] ? _0056_ : _0042_);
	assign _0097_ = _0096_ | ~_0072_;
	assign _0002_ = _0097_ | _0064_;
	assign _0098_ = (\mchip.micro_coded_cpu.cpu_fsm_top.cpu_state [0] ? \mchip.micro_coded_cpu.cpu_fsm_top.cpu_state [2] : \mchip.micro_coded_cpu.cpu_fsm_top.cpu_state [1]);
	assign _0099_ = _0055_ & ~_0041_;
	assign _0100_ = _0099_ | ~_0043_;
	assign _0101_ = _0100_ | _0046_;
	assign _0006_ = _0098_ & ~_0101_;
	assign _0102_ = \mchip.micro_coded_cpu.instr_reg_top.instr_reg [22] | ~\mchip.micro_coded_cpu.instr_reg_top.instr_reg [23];
	assign _0103_ = ~(_0102_ | _0051_);
	assign _0104_ = ~(_0103_ & _0047_);
	assign _0004_ = \mchip.micro_coded_cpu.mdecode_reg_top.reg_file_en  & ~_0104_;
	assign _0105_ = ~(\mchip.micro_coded_cpu.mdecode_reg_top.alu_en_A  | \mchip.micro_coded_cpu.mdecode_reg_top.alu_en_B );
	assign _0011_ = _0043_ & ~_0105_;
	assign _0010_ = _0047_ & \mchip.micro_coded_cpu.mdecode_reg_top.alu_en_B ;
	assign _0009_ = _0047_ & \mchip.micro_coded_cpu.mdecode_reg_top.alu_en_A ;
	assign _0106_ = ~\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [43];
	assign _0107_ = ~(\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [41] & \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [42]);
	assign _0108_ = _0106_ & ~_0107_;
	assign _0109_ = \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [41] | ~\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [42];
	assign _0110_ = _0106_ & ~_0109_;
	assign _0111_ = \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [42] | ~\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [41];
	assign _0112_ = _0106_ & ~_0111_;
	assign _0113_ = _0112_ | _0110_;
	assign \mchip.micro_coded_cpu.mdecode_reg_top.is_imm_active_md  = _0113_ | _0108_;
	assign _0114_ = ~\mchip.micro_coded_cpu.instr_reg_top.instr_reg [28];
	assign _0115_ = ~\mchip.micro_coded_cpu.instr_reg_top.instr_reg [29];
	assign _0116_ = (_0030_ ? _0114_ : _0115_);
	assign _0117_ = _0049_ & ~_0116_;
	assign _0118_ = ~\mchip.micro_coded_cpu.instr_reg_top.instr_reg [26];
	assign _0119_ = ~\mchip.micro_coded_cpu.instr_reg_top.instr_reg [27];
	assign _0120_ = (_0030_ ? _0118_ : _0119_);
	assign _0121_ = _0049_ & ~_0120_;
	assign _0122_ = (_0030_ ? _0119_ : _0114_);
	assign _0123_ = _0049_ & ~_0122_;
	assign _0124_ = _0121_ & ~_0123_;
	assign _0125_ = _0124_ & ~_0117_;
	assign _0126_ = ~\mchip.micro_coded_cpu.instr_reg_top.instr_reg [30];
	assign _0127_ = (_0030_ ? _0115_ : _0126_);
	assign _0128_ = _0049_ & ~_0127_;
	assign _0129_ = _0125_ & ~_0128_;
	assign _0130_ = (_0030_ ? \mchip.micro_coded_cpu.instr_reg_top.instr_reg [30] : \mchip.micro_coded_cpu.instr_reg_top.instr_reg [31]);
	assign _0131_ = _0130_ & ~io_in[13];
	assign _0132_ = ~_0128_;
	assign _0133_ = ~_0117_;
	assign _0134_ = _0123_ & _0121_;
	assign _0135_ = (_0117_ ? _0134_ : _0124_);
	assign _0136_ = ~_0121_;
	assign _0137_ = _0121_ | ~_0123_;
	assign _0138_ = (_0117_ ? _0137_ : _0136_);
	assign _0139_ = (_0128_ ? _0138_ : _0135_);
	assign _0000_[0] = (_0131_ ? _0129_ : _0139_);
	assign _0140_ = _0123_ | _0117_;
	assign _0141_ = _0132_ & ~_0140_;
	assign _0142_ = _0123_ & _0117_;
	assign _0143_ = (_0121_ ? _0123_ : _0117_);
	assign _0144_ = (_0128_ ? _0143_ : _0142_);
	assign _0000_[1] = (_0131_ ? _0141_ : _0144_);
	assign _0145_ = _0137_ | _0117_;
	assign _0146_ = _0132_ & ~_0145_;
	assign _0147_ = ~(_0123_ | _0121_);
	assign _0148_ = _0147_ & ~_0117_;
	assign _0149_ = _0128_ & ~_0148_;
	assign _0000_[2] = (_0131_ ? _0146_ : _0149_);
	assign _0150_ = _0134_ | _0117_;
	assign _0151_ = _0132_ & ~_0150_;
	assign _0152_ = _0124_ & ~_0133_;
	assign _0153_ = _0147_ ^ _0117_;
	assign _0154_ = (_0128_ ? _0153_ : _0152_);
	assign _0000_[3] = (_0131_ ? _0151_ : _0154_);
	assign _0155_ = ~\mchip.micro_coded_cpu.m_pc_top.m_pc [0];
	assign _0156_ = ~(\mchip.micro_coded_cpu.mdecode_reg_top.reg_dst [1] & \mchip.micro_coded_cpu.mdecode_reg_top.reg_dst [0]);
	assign _0157_ = \mchip.micro_coded_cpu.mdecode_reg_top.reg_dst [3] | \mchip.micro_coded_cpu.mdecode_reg_top.reg_dst [2];
	assign _0158_ = _0157_ | _0156_;
	assign _0159_ = _0158_ | \mchip.micro_coded_cpu.mdecode_reg_top.reg_dst [4];
	assign _0160_ = ~\mchip.micro_coded_cpu.alu_top.A_reg [0];
	assign _0161_ = \mchip.micro_coded_cpu.mdecode_reg_top.reg_dst [0] | ~\mchip.micro_coded_cpu.mdecode_reg_top.reg_dst [1];
	assign _0162_ = _0161_ | _0157_;
	assign _0163_ = _0162_ | \mchip.micro_coded_cpu.mdecode_reg_top.reg_dst [4];
	assign _0164_ = ~\mchip.micro_coded_cpu.mdecode_reg_top.reg_dst [4];
	assign _0165_ = \mchip.micro_coded_cpu.mdecode_reg_top.reg_dst [2] | ~\mchip.micro_coded_cpu.mdecode_reg_top.reg_dst [3];
	assign _0166_ = \mchip.micro_coded_cpu.mdecode_reg_top.reg_dst [1] | \mchip.micro_coded_cpu.mdecode_reg_top.reg_dst [0];
	assign _0167_ = _0166_ | _0165_;
	assign _0168_ = _0164_ & ~_0167_;
	assign _0169_ = _0168_ & \mchip.micro_coded_cpu.mdecode_reg_top.is_imm_active ;
	assign _0170_ = (_0163_ ? _0169_ : \mchip.micro_coded_cpu.alu_top.alu_result [0]);
	assign _0171_ = \mchip.micro_coded_cpu.mdecode_reg_top.reg_dst [1] | ~\mchip.micro_coded_cpu.mdecode_reg_top.reg_dst [0];
	assign _0172_ = _0171_ | _0157_;
	assign _0173_ = _0164_ & ~_0172_;
	assign _0174_ = _0173_ | ~_0170_;
	assign _0175_ = _0166_ | _0157_;
	assign _0176_ = _0164_ & ~_0175_;
	assign _0177_ = (_0176_ ? _0160_ : _0174_);
	assign _0178_ = \mchip.micro_coded_cpu.mdecode_reg_top.reg_dst [3] | ~\mchip.micro_coded_cpu.mdecode_reg_top.reg_dst [2];
	assign _0179_ = _0178_ | _0166_;
	assign _0180_ = _0164_ & ~_0179_;
	assign _0181_ = _0180_ | _0177_;
	assign _0182_ = _0159_ & ~_0181_;
	assign _0183_ = ~(_0182_ ^ \mchip.micro_coded_cpu.mdecode_reg_top.imm [0]);
	assign _0184_ = ~\mchip.micro_coded_cpu.alu_top.A_reg [1];
	assign _0185_ = _0163_ | ~\mchip.micro_coded_cpu.alu_top.alu_result [1];
	assign _0186_ = _0185_ | _0173_;
	assign _0187_ = (_0176_ ? _0184_ : _0186_);
	assign _0188_ = _0187_ | _0180_;
	assign _0189_ = _0159_ & ~_0188_;
	assign _0190_ = _0189_ ^ \mchip.micro_coded_cpu.mdecode_reg_top.imm [1];
	assign _0191_ = _0183_ & ~_0190_;
	assign _0192_ = ~\mchip.micro_coded_cpu.alu_top.A_reg [3];
	assign _0193_ = ~\mchip.micro_coded_cpu.alu_top.alu_result [3];
	assign _0194_ = _0163_ | _0193_;
	assign _0195_ = _0194_ | _0173_;
	assign _0196_ = (_0176_ ? _0192_ : _0195_);
	assign _0197_ = _0196_ | _0180_;
	assign _0198_ = _0159_ & ~_0197_;
	assign _0199_ = _0198_ ^ \mchip.micro_coded_cpu.mdecode_reg_top.imm [3];
	assign _0200_ = ~\mchip.micro_coded_cpu.alu_top.A_reg [2];
	assign _0201_ = ~\mchip.micro_coded_cpu.alu_top.alu_result [2];
	assign _0202_ = _0163_ | _0201_;
	assign _0203_ = _0202_ | _0173_;
	assign _0204_ = (_0176_ ? _0200_ : _0203_);
	assign _0205_ = _0204_ | _0180_;
	assign _0206_ = _0159_ & ~_0205_;
	assign _0207_ = _0206_ ^ \mchip.micro_coded_cpu.mdecode_reg_top.imm [2];
	assign _0208_ = _0207_ | _0199_;
	assign _0209_ = _0191_ & ~_0208_;
	assign _0210_ = ~\mchip.micro_coded_cpu.alu_top.A_reg [7];
	assign _0211_ = ~\mchip.micro_coded_cpu.alu_top.alu_result [7];
	assign _0212_ = _0163_ | _0211_;
	assign _0213_ = _0212_ | _0173_;
	assign _0214_ = (_0176_ ? _0210_ : _0213_);
	assign _0215_ = _0214_ | _0180_;
	assign _0216_ = _0159_ & ~_0215_;
	assign _0217_ = _0216_ ^ \mchip.micro_coded_cpu.mdecode_reg_top.imm [7];
	assign _0218_ = ~\mchip.micro_coded_cpu.alu_top.A_reg [6];
	assign _0219_ = ~\mchip.micro_coded_cpu.alu_top.alu_result [6];
	assign _0220_ = _0163_ | _0219_;
	assign _0221_ = _0220_ | _0173_;
	assign _0222_ = (_0176_ ? _0218_ : _0221_);
	assign _0223_ = _0222_ | _0180_;
	assign _0224_ = _0159_ & ~_0223_;
	assign _0225_ = _0224_ ^ \mchip.micro_coded_cpu.mdecode_reg_top.imm [6];
	assign _0226_ = _0225_ | _0217_;
	assign _0227_ = ~\mchip.micro_coded_cpu.alu_top.A_reg [5];
	assign _0228_ = ~\mchip.micro_coded_cpu.alu_top.alu_result [5];
	assign _0229_ = _0163_ | _0228_;
	assign _0230_ = _0229_ | _0173_;
	assign _0231_ = (_0176_ ? _0227_ : _0230_);
	assign _0232_ = _0231_ | _0180_;
	assign _0233_ = _0159_ & ~_0232_;
	assign _0234_ = _0233_ ^ \mchip.micro_coded_cpu.mdecode_reg_top.imm [5];
	assign _0235_ = ~\mchip.micro_coded_cpu.alu_top.A_reg [4];
	assign _0236_ = ~\mchip.micro_coded_cpu.alu_top.alu_result [4];
	assign _0237_ = _0163_ | _0236_;
	assign _0238_ = _0237_ | _0173_;
	assign _0239_ = (_0176_ ? _0235_ : _0238_);
	assign _0240_ = _0239_ | _0180_;
	assign _0241_ = _0159_ & ~_0240_;
	assign _0242_ = _0241_ ^ \mchip.micro_coded_cpu.mdecode_reg_top.imm [4];
	assign _0243_ = _0242_ | _0234_;
	assign _0244_ = _0243_ | _0226_;
	assign _0245_ = _0244_ | ~_0209_;
	assign _0246_ = _0047_ & ~_0245_;
	assign _0247_ = (_0246_ ? \mchip.micro_coded_cpu.mdecode_reg_top.mbranch_target [0] : _0155_);
	assign \mchip.micro_coded_cpu.m_pc_top.next_m_pc [0] = _0247_ & ~_0071_;
	assign _0248_ = \mchip.micro_coded_cpu.m_pc_top.m_pc [1] ^ \mchip.micro_coded_cpu.m_pc_top.m_pc [0];
	assign _0249_ = (_0246_ ? \mchip.micro_coded_cpu.mdecode_reg_top.mbranch_target [1] : _0248_);
	assign \mchip.micro_coded_cpu.m_pc_top.next_m_pc [1] = _0249_ & ~_0071_;
	assign _0250_ = ~_0071_;
	assign _0251_ = ~\mchip.micro_coded_cpu.mdecode_reg_top.mbranch_target [2];
	assign _0252_ = ~\mchip.micro_coded_cpu.m_pc_top.m_pc [2];
	assign _0253_ = \mchip.micro_coded_cpu.m_pc_top.m_pc [1] & \mchip.micro_coded_cpu.m_pc_top.m_pc [0];
	assign _0254_ = _0253_ ^ _0252_;
	assign _0255_ = (_0246_ ? _0251_ : _0254_);
	assign \mchip.micro_coded_cpu.m_pc_top.next_m_pc [2] = _0250_ & ~_0255_;
	assign _0256_ = ~\mchip.micro_coded_cpu.mdecode_reg_top.mbranch_target [3];
	assign _0257_ = ~\mchip.micro_coded_cpu.m_pc_top.m_pc [3];
	assign _0258_ = _0253_ & ~_0252_;
	assign _0259_ = _0258_ ^ _0257_;
	assign _0260_ = (_0246_ ? _0256_ : _0259_);
	assign \mchip.micro_coded_cpu.m_pc_top.next_m_pc [3] = _0250_ & ~_0260_;
	assign _0261_ = ~\mchip.micro_coded_cpu.mdecode_reg_top.mbranch_target [4];
	assign _0262_ = ~\mchip.micro_coded_cpu.m_pc_top.m_pc [4];
	assign _0263_ = ~(\mchip.micro_coded_cpu.m_pc_top.m_pc [3] & \mchip.micro_coded_cpu.m_pc_top.m_pc [2]);
	assign _0264_ = _0253_ & ~_0263_;
	assign _0265_ = _0264_ ^ _0262_;
	assign _0266_ = (_0246_ ? _0261_ : _0265_);
	assign \mchip.micro_coded_cpu.m_pc_top.next_m_pc [4] = _0250_ & ~_0266_;
	assign _0267_ = ~\mchip.micro_coded_cpu.mdecode_reg_top.mbranch_target [5];
	assign _0268_ = ~\mchip.micro_coded_cpu.m_pc_top.m_pc [5];
	assign _0269_ = _0264_ & ~_0262_;
	assign _0270_ = _0269_ ^ _0268_;
	assign _0271_ = (_0246_ ? _0267_ : _0270_);
	assign \mchip.micro_coded_cpu.m_pc_top.next_m_pc [5] = _0250_ & ~_0271_;
	assign _0272_ = ~\mchip.micro_coded_cpu.mdecode_reg_top.mbranch_target [6];
	assign _0273_ = ~\mchip.micro_coded_cpu.m_pc_top.m_pc [6];
	assign _0274_ = ~(\mchip.micro_coded_cpu.m_pc_top.m_pc [5] & \mchip.micro_coded_cpu.m_pc_top.m_pc [4]);
	assign _0275_ = _0264_ & ~_0274_;
	assign _0276_ = _0275_ ^ _0273_;
	assign _0277_ = (_0246_ ? _0272_ : _0276_);
	assign \mchip.micro_coded_cpu.m_pc_top.next_m_pc [6] = _0250_ & ~_0277_;
	assign _0278_ = ~\mchip.micro_coded_cpu.mdecode_reg_top.mbranch_target [7];
	assign _0279_ = ~\mchip.micro_coded_cpu.m_pc_top.m_pc [7];
	assign _0280_ = _0275_ & ~_0273_;
	assign _0281_ = _0280_ ^ _0279_;
	assign _0282_ = (_0246_ ? _0278_ : _0281_);
	assign \mchip.micro_coded_cpu.m_pc_top.next_m_pc [7] = _0250_ & ~_0282_;
	assign _0283_ = _0099_ & ~_0031_;
	assign _0284_ = _0081_ & ~_0283_;
	assign _0285_ = _0250_ & ~_0284_;
	assign _0286_ = _0057_ & ~_0285_;
	assign _0023_ = _0286_ | _0064_;
	assign _0287_ = \mchip.micro_coded_cpu.cpu_fsm_top.current_minst_1 [0] & \mchip.micro_coded_cpu.cpu_fsm_top.current_minst_1 [1];
	assign _0288_ = ~(\mchip.micro_coded_cpu.cpu_fsm_top.current_minst_1 [2] & \mchip.micro_coded_cpu.cpu_fsm_top.current_minst_1 [3]);
	assign _0289_ = _0287_ & ~_0288_;
	assign _0290_ = _0289_ & \mchip.micro_coded_cpu.cpu_fsm_top.current_minst_1 [4];
	assign _0291_ = _0290_ & ~_0047_;
	assign _0292_ = _0291_ & ~_0099_;
	assign _0293_ = _0292_ | _0031_;
	assign _0294_ = _0081_ & ~_0293_;
	assign _0295_ = _0294_ | _0071_;
	assign _0296_ = _0057_ & ~_0295_;
	assign _0024_ = _0065_ & ~_0296_;
	assign _0297_ = _0099_ | _0047_;
	assign _0298_ = _0297_ | _0031_;
	assign _0299_ = _0081_ & ~_0298_;
	assign _0300_ = _0299_ | _0071_;
	assign _0301_ = _0300_ | _0030_;
	assign _0025_ = _0065_ & ~_0301_;
	assign _0302_ = (_0050_ ? _0084_ : _0076_);
	assign _0303_ = _0302_ | \mchip.micro_coded_cpu.cpu_fsm_top.fsm_assist [0];
	assign _0304_ = _0250_ & ~_0303_;
	assign _0305_ = ~(_0062_ | \mchip.micro_coded_cpu.cpu_fsm_top.fsm_assist [0]);
	assign _0306_ = (_0030_ ? _0305_ : _0304_);
	assign _0307_ = ~(_0069_ | \mchip.micro_coded_cpu.cpu_fsm_top.fsm_assist [0]);
	assign _0017_ = (_0064_ ? _0307_ : _0306_);
	assign _0308_ = _0058_ | ~_0082_;
	assign _0309_ = _0308_ | _0302_;
	assign _0310_ = _0250_ & ~_0309_;
	assign _0311_ = ~(_0308_ | _0062_);
	assign _0312_ = (_0030_ ? _0311_ : _0310_);
	assign _0313_ = ~(_0308_ | _0069_);
	assign _0018_ = (_0064_ ? _0313_ : _0312_);
	assign _0314_ = ~(_0058_ ^ \mchip.micro_coded_cpu.cpu_fsm_top.fsm_assist [2]);
	assign _0315_ = _0314_ | _0302_;
	assign _0316_ = _0250_ & ~_0315_;
	assign _0317_ = ~(_0314_ | _0062_);
	assign _0318_ = (_0030_ ? _0317_ : _0316_);
	assign _0319_ = ~(_0314_ | _0069_);
	assign _0019_ = (_0064_ ? _0319_ : _0318_);
	assign _0320_ = ~(_0058_ & \mchip.micro_coded_cpu.cpu_fsm_top.fsm_assist [2]);
	assign _0321_ = _0320_ ^ \mchip.micro_coded_cpu.cpu_fsm_top.fsm_assist [3];
	assign _0322_ = _0321_ | _0302_;
	assign _0323_ = _0250_ & ~_0322_;
	assign _0324_ = ~(_0321_ | _0062_);
	assign _0325_ = (_0030_ ? _0324_ : _0323_);
	assign _0326_ = ~(_0321_ | _0069_);
	assign _0020_ = (_0064_ ? _0326_ : _0325_);
	assign _0327_ = ~(_0060_ ^ \mchip.micro_coded_cpu.cpu_fsm_top.fsm_assist [4]);
	assign _0328_ = _0327_ | _0302_;
	assign _0329_ = _0250_ & ~_0328_;
	assign _0330_ = ~(_0327_ | _0062_);
	assign _0331_ = (_0030_ ? _0330_ : _0329_);
	assign _0332_ = ~(_0327_ | _0069_);
	assign _0021_ = (_0064_ ? _0332_ : _0331_);
	assign _0333_ = ~(_0060_ & \mchip.micro_coded_cpu.cpu_fsm_top.fsm_assist [4]);
	assign _0334_ = _0333_ ^ \mchip.micro_coded_cpu.cpu_fsm_top.fsm_assist [5];
	assign _0335_ = _0334_ | _0302_;
	assign _0336_ = _0250_ & ~_0335_;
	assign _0337_ = ~(_0334_ | _0062_);
	assign _0338_ = (_0030_ ? _0337_ : _0336_);
	assign _0339_ = ~(_0334_ | _0069_);
	assign _0022_ = (_0064_ ? _0339_ : _0338_);
	assign _0012_ = ~(_0290_ | \mchip.micro_coded_cpu.cpu_fsm_top.current_minst_1 [0]);
	assign _0013_ = \mchip.micro_coded_cpu.cpu_fsm_top.current_minst_1 [0] ^ \mchip.micro_coded_cpu.cpu_fsm_top.current_minst_1 [1];
	assign _0340_ = _0287_ ^ \mchip.micro_coded_cpu.cpu_fsm_top.current_minst_1 [2];
	assign _0014_ = _0340_ & ~_0290_;
	assign _0341_ = _0287_ & \mchip.micro_coded_cpu.cpu_fsm_top.current_minst_1 [2];
	assign _0342_ = _0341_ ^ \mchip.micro_coded_cpu.cpu_fsm_top.current_minst_1 [3];
	assign _0015_ = _0342_ & ~_0290_;
	assign _0016_ = _0289_ ^ \mchip.micro_coded_cpu.cpu_fsm_top.current_minst_1 [4];
	assign _0343_ = \mchip.micro_coded_cpu.mdecode_reg_top.reg_src [0] | ~\mchip.micro_coded_cpu.mdecode_reg_top.reg_src [1];
	assign _0344_ = ~(\mchip.micro_coded_cpu.mdecode_reg_top.reg_src [2] & \mchip.micro_coded_cpu.mdecode_reg_top.reg_src [3]);
	assign _0345_ = _0344_ | _0343_;
	assign _0346_ = _0345_ | \mchip.micro_coded_cpu.mdecode_reg_top.reg_src [4];
	assign _0347_ = \mchip.micro_coded_cpu.mdecode_reg_top.reg_src [3] | ~\mchip.micro_coded_cpu.mdecode_reg_top.reg_src [2];
	assign _0348_ = ~(\mchip.micro_coded_cpu.mdecode_reg_top.reg_src [1] & \mchip.micro_coded_cpu.mdecode_reg_top.reg_src [0]);
	assign _0349_ = _0348_ | _0347_;
	assign _0350_ = _0349_ | \mchip.micro_coded_cpu.mdecode_reg_top.reg_src [4];
	assign _0351_ = \mchip.micro_coded_cpu.reg_file_interface.reg_rd_data_out [0] & ~_0350_;
	assign _0352_ = ~\mchip.micro_coded_cpu.mdecode_reg_top.reg_src [4];
	assign _0353_ = \mchip.micro_coded_cpu.mdecode_reg_top.reg_src [2] | \mchip.micro_coded_cpu.mdecode_reg_top.reg_src [3];
	assign _0354_ = _0353_ | _0343_;
	assign _0355_ = _0352_ & ~_0354_;
	assign _0356_ = (_0355_ ? \mchip.micro_coded_cpu.alu_top.alu_result [0] : _0351_);
	assign _0357_ = \mchip.micro_coded_cpu.mdecode_reg_top.reg_src [1] | ~\mchip.micro_coded_cpu.mdecode_reg_top.reg_src [0];
	assign _0358_ = _0357_ | _0353_;
	assign _0359_ = \mchip.micro_coded_cpu.mdecode_reg_top.reg_src [4] & ~_0358_;
	assign _0360_ = (_0359_ ? \mchip.micro_coded_cpu.mdecode_reg_top.mbranch_target [0] : _0356_);
	assign _0361_ = _0357_ | _0344_;
	assign _0362_ = _0352_ & ~_0361_;
	assign _0363_ = (_0362_ ? \mchip.micro_coded_cpu.m_pc_top.m_pc [0] : _0360_);
	assign _0364_ = \mchip.micro_coded_cpu.mdecode_reg_top.reg_src [2] | ~\mchip.micro_coded_cpu.mdecode_reg_top.reg_src [3];
	assign _0365_ = _0364_ | _0357_;
	assign _0366_ = _0352_ & ~_0365_;
	assign _0367_ = (_0366_ ? \mchip.micro_coded_cpu.mdecode_reg_top.imm [0] : _0363_);
	assign _0368_ = _0348_ | _0344_;
	assign _0369_ = _0352_ & ~_0368_;
	assign _0370_ = (_0369_ ? \mchip.micro_coded_cpu.instr_reg_top.instr_reg [14] : _0367_);
	assign _0371_ = (_0346_ ? _0370_ : \mchip.micro_coded_cpu.instr_reg_top.instr_reg [18]);
	assign _0372_ = \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [41] | \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [42];
	assign _0373_ = \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [43] & ~_0372_;
	assign _0374_ = (_0373_ ? \mchip.micro_coded_cpu.mdecode_reg_top.mbranch_target [0] : _0371_);
	assign _0375_ = (_0245_ ? \mchip.micro_coded_cpu.m_pc_top.m_pc [0] : \mchip.micro_coded_cpu.mdecode_reg_top.mbranch_target [0]);
	assign \mchip.micro_coded_cpu.alu_top.A_bus [0] = (_0108_ ? _0375_ : _0374_);
	assign _0376_ = \mchip.micro_coded_cpu.reg_file_interface.reg_rd_data_out [1] & ~_0350_;
	assign _0377_ = (_0355_ ? \mchip.micro_coded_cpu.alu_top.alu_result [1] : _0376_);
	assign _0378_ = (_0359_ ? \mchip.micro_coded_cpu.mdecode_reg_top.mbranch_target [1] : _0377_);
	assign _0379_ = (_0362_ ? \mchip.micro_coded_cpu.m_pc_top.m_pc [1] : _0378_);
	assign _0380_ = (_0366_ ? \mchip.micro_coded_cpu.mdecode_reg_top.imm [1] : _0379_);
	assign _0381_ = (_0369_ ? \mchip.micro_coded_cpu.instr_reg_top.instr_reg [15] : _0380_);
	assign _0382_ = (_0346_ ? _0381_ : \mchip.micro_coded_cpu.instr_reg_top.instr_reg [19]);
	assign _0383_ = (_0373_ ? \mchip.micro_coded_cpu.mdecode_reg_top.mbranch_target [1] : _0382_);
	assign _0384_ = (_0245_ ? \mchip.micro_coded_cpu.m_pc_top.m_pc [1] : \mchip.micro_coded_cpu.mdecode_reg_top.mbranch_target [1]);
	assign \mchip.micro_coded_cpu.alu_top.A_bus [1] = (_0108_ ? _0384_ : _0383_);
	assign _0385_ = ~\mchip.micro_coded_cpu.mdecode_reg_top.imm [2];
	assign _0386_ = _0350_ | ~\mchip.micro_coded_cpu.reg_file_interface.reg_rd_data_out [2];
	assign _0387_ = (_0355_ ? _0201_ : _0386_);
	assign _0388_ = (_0359_ ? _0251_ : _0387_);
	assign _0389_ = (_0362_ ? _0252_ : _0388_);
	assign _0390_ = (_0366_ ? _0385_ : _0389_);
	assign _0391_ = _0390_ | _0369_;
	assign _0392_ = _0346_ & ~_0391_;
	assign _0393_ = (_0373_ ? \mchip.micro_coded_cpu.mdecode_reg_top.mbranch_target [2] : _0392_);
	assign _0394_ = (_0245_ ? \mchip.micro_coded_cpu.m_pc_top.m_pc [2] : \mchip.micro_coded_cpu.mdecode_reg_top.mbranch_target [2]);
	assign \mchip.micro_coded_cpu.alu_top.A_bus [2] = (_0108_ ? _0394_ : _0393_);
	assign _0395_ = ~\mchip.micro_coded_cpu.mdecode_reg_top.imm [3];
	assign _0396_ = _0350_ | ~\mchip.micro_coded_cpu.reg_file_interface.reg_rd_data_out [3];
	assign _0397_ = (_0355_ ? _0193_ : _0396_);
	assign _0398_ = (_0359_ ? _0256_ : _0397_);
	assign _0399_ = (_0362_ ? _0257_ : _0398_);
	assign _0400_ = (_0366_ ? _0395_ : _0399_);
	assign _0401_ = _0400_ | _0369_;
	assign _0402_ = _0346_ & ~_0401_;
	assign _0403_ = (_0373_ ? \mchip.micro_coded_cpu.mdecode_reg_top.mbranch_target [3] : _0402_);
	assign _0404_ = (_0245_ ? \mchip.micro_coded_cpu.m_pc_top.m_pc [3] : \mchip.micro_coded_cpu.mdecode_reg_top.mbranch_target [3]);
	assign \mchip.micro_coded_cpu.alu_top.A_bus [3] = (_0108_ ? _0404_ : _0403_);
	assign _0405_ = ~\mchip.micro_coded_cpu.mdecode_reg_top.imm [4];
	assign _0406_ = _0350_ | ~\mchip.micro_coded_cpu.reg_file_interface.reg_rd_data_out [4];
	assign _0407_ = (_0355_ ? _0236_ : _0406_);
	assign _0408_ = (_0359_ ? _0261_ : _0407_);
	assign _0409_ = (_0362_ ? _0262_ : _0408_);
	assign _0410_ = (_0366_ ? _0405_ : _0409_);
	assign _0411_ = _0410_ | _0369_;
	assign _0412_ = _0346_ & ~_0411_;
	assign _0413_ = (_0373_ ? \mchip.micro_coded_cpu.mdecode_reg_top.mbranch_target [4] : _0412_);
	assign _0414_ = (_0245_ ? \mchip.micro_coded_cpu.m_pc_top.m_pc [4] : \mchip.micro_coded_cpu.mdecode_reg_top.mbranch_target [4]);
	assign \mchip.micro_coded_cpu.alu_top.A_bus [4] = (_0108_ ? _0414_ : _0413_);
	assign _0415_ = ~\mchip.micro_coded_cpu.mdecode_reg_top.imm [5];
	assign _0416_ = _0350_ | ~\mchip.micro_coded_cpu.reg_file_interface.reg_rd_data_out [5];
	assign _0417_ = (_0355_ ? _0228_ : _0416_);
	assign _0418_ = (_0359_ ? _0267_ : _0417_);
	assign _0419_ = (_0362_ ? _0268_ : _0418_);
	assign _0420_ = (_0366_ ? _0415_ : _0419_);
	assign _0421_ = _0420_ | _0369_;
	assign _0422_ = _0346_ & ~_0421_;
	assign _0423_ = (_0373_ ? \mchip.micro_coded_cpu.mdecode_reg_top.mbranch_target [5] : _0422_);
	assign _0424_ = (_0245_ ? \mchip.micro_coded_cpu.m_pc_top.m_pc [5] : \mchip.micro_coded_cpu.mdecode_reg_top.mbranch_target [5]);
	assign \mchip.micro_coded_cpu.alu_top.A_bus [5] = (_0108_ ? _0424_ : _0423_);
	assign _0425_ = ~\mchip.micro_coded_cpu.mdecode_reg_top.imm [6];
	assign _0426_ = _0350_ | ~\mchip.micro_coded_cpu.reg_file_interface.reg_rd_data_out [6];
	assign _0427_ = (_0355_ ? _0219_ : _0426_);
	assign _0428_ = (_0359_ ? _0272_ : _0427_);
	assign _0429_ = (_0362_ ? _0273_ : _0428_);
	assign _0430_ = (_0366_ ? _0425_ : _0429_);
	assign _0431_ = _0430_ | _0369_;
	assign _0432_ = _0346_ & ~_0431_;
	assign _0433_ = (_0373_ ? \mchip.micro_coded_cpu.mdecode_reg_top.mbranch_target [6] : _0432_);
	assign _0434_ = (_0245_ ? \mchip.micro_coded_cpu.m_pc_top.m_pc [6] : \mchip.micro_coded_cpu.mdecode_reg_top.mbranch_target [6]);
	assign \mchip.micro_coded_cpu.alu_top.A_bus [6] = (_0108_ ? _0434_ : _0433_);
	assign _0435_ = ~\mchip.micro_coded_cpu.mdecode_reg_top.imm [7];
	assign _0436_ = _0350_ | ~\mchip.micro_coded_cpu.reg_file_interface.reg_rd_data_out [7];
	assign _0437_ = (_0355_ ? _0211_ : _0436_);
	assign _0438_ = (_0359_ ? _0278_ : _0437_);
	assign _0439_ = (_0362_ ? _0279_ : _0438_);
	assign _0440_ = (_0366_ ? _0435_ : _0439_);
	assign _0441_ = _0440_ | _0369_;
	assign _0442_ = _0346_ & ~_0441_;
	assign _0443_ = (_0373_ ? \mchip.micro_coded_cpu.mdecode_reg_top.mbranch_target [7] : _0442_);
	assign _0444_ = (_0245_ ? \mchip.micro_coded_cpu.m_pc_top.m_pc [7] : \mchip.micro_coded_cpu.mdecode_reg_top.mbranch_target [7]);
	assign \mchip.micro_coded_cpu.alu_top.A_bus [7] = (_0108_ ? _0444_ : _0443_);
	assign _0445_ = (\mchip.micro_coded_cpu.reg_file_interface.reg_sel_in [0] ? \mchip.micro_coded_cpu.reg_file_interface.mreg_file[1] [0] : \mchip.micro_coded_cpu.reg_file_interface.mreg_file[0] [0]);
	assign _0446_ = (\mchip.micro_coded_cpu.reg_file_interface.reg_sel_in [0] ? \mchip.micro_coded_cpu.reg_file_interface.mreg_file[3] [0] : \mchip.micro_coded_cpu.reg_file_interface.mreg_file[2] [0]);
	assign _0001_[0] = (\mchip.micro_coded_cpu.reg_file_interface.reg_sel_in [1] ? _0446_ : _0445_);
	assign _0447_ = (\mchip.micro_coded_cpu.reg_file_interface.reg_sel_in [0] ? \mchip.micro_coded_cpu.reg_file_interface.mreg_file[1] [1] : \mchip.micro_coded_cpu.reg_file_interface.mreg_file[0] [1]);
	assign _0448_ = (\mchip.micro_coded_cpu.reg_file_interface.reg_sel_in [0] ? \mchip.micro_coded_cpu.reg_file_interface.mreg_file[3] [1] : \mchip.micro_coded_cpu.reg_file_interface.mreg_file[2] [1]);
	assign _0001_[1] = (\mchip.micro_coded_cpu.reg_file_interface.reg_sel_in [1] ? _0448_ : _0447_);
	assign _0449_ = (\mchip.micro_coded_cpu.reg_file_interface.reg_sel_in [0] ? \mchip.micro_coded_cpu.reg_file_interface.mreg_file[1] [2] : \mchip.micro_coded_cpu.reg_file_interface.mreg_file[0] [2]);
	assign _0450_ = (\mchip.micro_coded_cpu.reg_file_interface.reg_sel_in [0] ? \mchip.micro_coded_cpu.reg_file_interface.mreg_file[3] [2] : \mchip.micro_coded_cpu.reg_file_interface.mreg_file[2] [2]);
	assign _0001_[2] = (\mchip.micro_coded_cpu.reg_file_interface.reg_sel_in [1] ? _0450_ : _0449_);
	assign _0451_ = (\mchip.micro_coded_cpu.reg_file_interface.reg_sel_in [0] ? \mchip.micro_coded_cpu.reg_file_interface.mreg_file[1] [3] : \mchip.micro_coded_cpu.reg_file_interface.mreg_file[0] [3]);
	assign _0452_ = (\mchip.micro_coded_cpu.reg_file_interface.reg_sel_in [0] ? \mchip.micro_coded_cpu.reg_file_interface.mreg_file[3] [3] : \mchip.micro_coded_cpu.reg_file_interface.mreg_file[2] [3]);
	assign _0001_[3] = (\mchip.micro_coded_cpu.reg_file_interface.reg_sel_in [1] ? _0452_ : _0451_);
	assign _0453_ = (\mchip.micro_coded_cpu.reg_file_interface.reg_sel_in [0] ? \mchip.micro_coded_cpu.reg_file_interface.mreg_file[1] [4] : \mchip.micro_coded_cpu.reg_file_interface.mreg_file[0] [4]);
	assign _0454_ = (\mchip.micro_coded_cpu.reg_file_interface.reg_sel_in [0] ? \mchip.micro_coded_cpu.reg_file_interface.mreg_file[3] [4] : \mchip.micro_coded_cpu.reg_file_interface.mreg_file[2] [4]);
	assign _0001_[4] = (\mchip.micro_coded_cpu.reg_file_interface.reg_sel_in [1] ? _0454_ : _0453_);
	assign _0455_ = (\mchip.micro_coded_cpu.reg_file_interface.reg_sel_in [0] ? \mchip.micro_coded_cpu.reg_file_interface.mreg_file[1] [5] : \mchip.micro_coded_cpu.reg_file_interface.mreg_file[0] [5]);
	assign _0456_ = (\mchip.micro_coded_cpu.reg_file_interface.reg_sel_in [0] ? \mchip.micro_coded_cpu.reg_file_interface.mreg_file[3] [5] : \mchip.micro_coded_cpu.reg_file_interface.mreg_file[2] [5]);
	assign _0001_[5] = (\mchip.micro_coded_cpu.reg_file_interface.reg_sel_in [1] ? _0456_ : _0455_);
	assign _0457_ = (\mchip.micro_coded_cpu.reg_file_interface.reg_sel_in [0] ? \mchip.micro_coded_cpu.reg_file_interface.mreg_file[1] [6] : \mchip.micro_coded_cpu.reg_file_interface.mreg_file[0] [6]);
	assign _0458_ = (\mchip.micro_coded_cpu.reg_file_interface.reg_sel_in [0] ? \mchip.micro_coded_cpu.reg_file_interface.mreg_file[3] [6] : \mchip.micro_coded_cpu.reg_file_interface.mreg_file[2] [6]);
	assign _0001_[6] = (\mchip.micro_coded_cpu.reg_file_interface.reg_sel_in [1] ? _0458_ : _0457_);
	assign _0459_ = (\mchip.micro_coded_cpu.reg_file_interface.reg_sel_in [0] ? \mchip.micro_coded_cpu.reg_file_interface.mreg_file[1] [7] : \mchip.micro_coded_cpu.reg_file_interface.mreg_file[0] [7]);
	assign _0460_ = (\mchip.micro_coded_cpu.reg_file_interface.reg_sel_in [0] ? \mchip.micro_coded_cpu.reg_file_interface.mreg_file[3] [7] : \mchip.micro_coded_cpu.reg_file_interface.mreg_file[2] [7]);
	assign _0001_[7] = (\mchip.micro_coded_cpu.reg_file_interface.reg_sel_in [1] ? _0460_ : _0459_);
	assign _0461_ = ~\mchip.micro_coded_cpu.m_pc_top.m_pc [1];
	assign _0462_ = (\mchip.micro_coded_cpu.m_inst_to_bit.current_bit_index [0] ? _0461_ : _0155_);
	assign _0463_ = (\mchip.micro_coded_cpu.m_inst_to_bit.current_bit_index [0] ? _0257_ : _0252_);
	assign _0464_ = (\mchip.micro_coded_cpu.m_inst_to_bit.current_bit_index [1] ? _0463_ : _0462_);
	assign _0465_ = ~(\mchip.micro_coded_cpu.m_inst_addr_offset [5] ^ \mchip.micro_coded_cpu.m_pc_top.m_pc [5]);
	assign _0466_ = (\mchip.micro_coded_cpu.m_inst_to_bit.current_bit_index [0] ? _0465_ : _0262_);
	assign _0467_ = \mchip.micro_coded_cpu.m_inst_addr_offset [5] & \mchip.micro_coded_cpu.m_pc_top.m_pc [5];
	assign _0468_ = \mchip.micro_coded_cpu.m_inst_addr_offset [6] ^ \mchip.micro_coded_cpu.m_pc_top.m_pc [6];
	assign _0469_ = ~(_0468_ ^ _0467_);
	assign _0470_ = \mchip.micro_coded_cpu.m_inst_addr_offset [6] & \mchip.micro_coded_cpu.m_pc_top.m_pc [6];
	assign _0471_ = _0468_ & _0467_;
	assign _0472_ = ~(_0471_ | _0470_);
	assign _0473_ = ~(\mchip.micro_coded_cpu.m_inst_addr_offset [7] ^ \mchip.micro_coded_cpu.m_pc_top.m_pc [7]);
	assign _0474_ = ~(_0473_ ^ _0472_);
	assign _0475_ = (\mchip.micro_coded_cpu.m_inst_to_bit.current_bit_index [0] ? _0474_ : _0469_);
	assign _0476_ = (\mchip.micro_coded_cpu.m_inst_to_bit.current_bit_index [1] ? _0475_ : _0466_);
	assign _0477_ = (\mchip.micro_coded_cpu.m_inst_to_bit.current_bit_index [2] ? _0476_ : _0464_);
	assign _0478_ = _0473_ | _0472_;
	assign _0479_ = \mchip.micro_coded_cpu.m_inst_addr_offset [7] & \mchip.micro_coded_cpu.m_pc_top.m_pc [7];
	assign _0480_ = _0478_ & ~_0479_;
	assign _0481_ = _0480_ ^ \mchip.micro_coded_cpu.m_inst_addr_offset [8];
	assign _0482_ = _0481_ | \mchip.micro_coded_cpu.m_inst_to_bit.current_bit_index [0];
	assign _0483_ = _0482_ | \mchip.micro_coded_cpu.m_inst_to_bit.current_bit_index [1];
	assign _0484_ = _0483_ | \mchip.micro_coded_cpu.m_inst_to_bit.current_bit_index [2];
	assign _0485_ = (\mchip.micro_coded_cpu.m_inst_to_bit.current_bit_index [3] ? _0484_ : _0477_);
	assign _0486_ = _0485_ | _0081_;
	assign \mchip.micro_coded_cpu.m_inst_addr_stream  = _0049_ & ~_0486_;
	assign _0487_ = ~\mchip.micro_coded_cpu.mdecode_reg_top.alu_op [2];
	assign _0488_ = ~(\mchip.micro_coded_cpu.mdecode_reg_top.alu_op [1] & \mchip.micro_coded_cpu.mdecode_reg_top.alu_op [0]);
	assign _0489_ = _0487_ & ~_0488_;
	assign _0490_ = \mchip.micro_coded_cpu.mdecode_reg_top.alu_op [1] | ~\mchip.micro_coded_cpu.mdecode_reg_top.alu_op [0];
	assign _0491_ = _0487_ & ~_0490_;
	assign _0492_ = \mchip.micro_coded_cpu.mdecode_reg_top.alu_op [0] | ~\mchip.micro_coded_cpu.mdecode_reg_top.alu_op [1];
	assign _0493_ = _0487_ & ~_0492_;
	assign _0494_ = ~(_0493_ | _0491_);
	assign _0495_ = _0489_ | ~_0494_;
	assign _0496_ = \mchip.micro_coded_cpu.mdecode_reg_top.alu_op [2] & ~\mchip.micro_coded_cpu.mdecode_reg_top.alu_op [1];
	assign _0497_ = \mchip.micro_coded_cpu.mdecode_reg_top.alu_op [1] & \mchip.micro_coded_cpu.mdecode_reg_top.alu_op [2];
	assign _0498_ = _0497_ | _0496_;
	assign _0499_ = _0498_ | _0495_;
	assign _0500_ = \mchip.micro_coded_cpu.alu_top.B_reg [0] & \mchip.micro_coded_cpu.alu_top.A_reg [0];
	assign _0501_ = ~(\mchip.micro_coded_cpu.alu_top.B_reg [0] | \mchip.micro_coded_cpu.alu_top.A_reg [0]);
	assign _0502_ = _0501_ | _0500_;
	assign _0503_ = _0502_ | _0494_;
	assign _0504_ = _0489_ & ~_0501_;
	assign _0505_ = _0503_ & ~_0504_;
	assign _0506_ = \mchip.micro_coded_cpu.mdecode_reg_top.alu_op [1] | \mchip.micro_coded_cpu.mdecode_reg_top.alu_op [0];
	assign _0507_ = \mchip.micro_coded_cpu.mdecode_reg_top.alu_op [2] & ~_0506_;
	assign _0508_ = _0507_ & _0500_;
	assign _0509_ = _0490_ | _0487_;
	assign _0510_ = _0160_ & ~_0509_;
	assign _0511_ = _0510_ | _0508_;
	assign _0512_ = \mchip.micro_coded_cpu.mdecode_reg_top.alu_op [2] & ~_0492_;
	assign _0513_ = \mchip.micro_coded_cpu.alu_top.B_reg [6] | \mchip.micro_coded_cpu.alu_top.B_reg [7];
	assign _0514_ = \mchip.micro_coded_cpu.alu_top.B_reg [4] | \mchip.micro_coded_cpu.alu_top.B_reg [5];
	assign _0515_ = _0514_ | _0513_;
	assign _0516_ = _0515_ | _0160_;
	assign _0517_ = _0516_ | \mchip.micro_coded_cpu.alu_top.B_reg [0];
	assign _0518_ = _0517_ | \mchip.micro_coded_cpu.alu_top.B_reg [1];
	assign _0519_ = _0518_ | \mchip.micro_coded_cpu.alu_top.B_reg [2];
	assign _0520_ = _0519_ | \mchip.micro_coded_cpu.alu_top.B_reg [3];
	assign _0521_ = _0512_ & ~_0520_;
	assign _0522_ = ~\mchip.micro_coded_cpu.alu_top.B_reg [3];
	assign _0523_ = ~\mchip.micro_coded_cpu.alu_top.B_reg [2];
	assign _0524_ = _0515_ | _0184_;
	assign _0525_ = (\mchip.micro_coded_cpu.alu_top.B_reg [0] ? _0524_ : _0516_);
	assign _0526_ = _0515_ | _0200_;
	assign _0527_ = _0515_ | _0192_;
	assign _0528_ = (\mchip.micro_coded_cpu.alu_top.B_reg [0] ? _0527_ : _0526_);
	assign _0529_ = (\mchip.micro_coded_cpu.alu_top.B_reg [1] ? _0528_ : _0525_);
	assign _0530_ = _0515_ | _0235_;
	assign _0531_ = _0515_ | _0227_;
	assign _0532_ = (\mchip.micro_coded_cpu.alu_top.B_reg [0] ? _0531_ : _0530_);
	assign _0533_ = _0515_ | _0218_;
	assign _0534_ = _0515_ | _0210_;
	assign _0535_ = (\mchip.micro_coded_cpu.alu_top.B_reg [0] ? _0534_ : _0533_);
	assign _0536_ = (\mchip.micro_coded_cpu.alu_top.B_reg [1] ? _0535_ : _0532_);
	assign _0537_ = (\mchip.micro_coded_cpu.alu_top.B_reg [2] ? _0536_ : _0529_);
	assign _0538_ = _0522_ & ~_0537_;
	assign _0539_ = _0488_ | _0487_;
	assign _0540_ = _0538_ & ~_0539_;
	assign _0541_ = _0540_ | _0521_;
	assign _0542_ = _0541_ | _0511_;
	assign _0543_ = _0505_ & ~_0542_;
	assign \mchip.micro_coded_cpu.alu_top.alu_result_out [0] = _0499_ & ~_0543_;
	assign _0544_ = (\mchip.micro_coded_cpu.alu_top.B_reg [0] ? _0526_ : _0524_);
	assign _0545_ = (\mchip.micro_coded_cpu.alu_top.B_reg [0] ? _0530_ : _0527_);
	assign _0546_ = (\mchip.micro_coded_cpu.alu_top.B_reg [1] ? _0545_ : _0544_);
	assign _0547_ = (\mchip.micro_coded_cpu.alu_top.B_reg [0] ? _0533_ : _0531_);
	assign _0548_ = _0534_ | \mchip.micro_coded_cpu.alu_top.B_reg [0];
	assign _0549_ = (\mchip.micro_coded_cpu.alu_top.B_reg [1] ? _0548_ : _0547_);
	assign _0550_ = (\mchip.micro_coded_cpu.alu_top.B_reg [2] ? _0549_ : _0546_);
	assign _0551_ = _0550_ | \mchip.micro_coded_cpu.alu_top.B_reg [3];
	assign _0552_ = _0551_ | _0539_;
	assign _0553_ = (\mchip.micro_coded_cpu.alu_top.B_reg [0] ? _0516_ : _0524_);
	assign _0554_ = _0553_ | \mchip.micro_coded_cpu.alu_top.B_reg [1];
	assign _0555_ = _0554_ | \mchip.micro_coded_cpu.alu_top.B_reg [2];
	assign _0556_ = _0555_ | \mchip.micro_coded_cpu.alu_top.B_reg [3];
	assign _0557_ = _0512_ & ~_0556_;
	assign _0558_ = _0552_ & ~_0557_;
	assign _0559_ = ~(\mchip.micro_coded_cpu.alu_top.B_reg [1] & \mchip.micro_coded_cpu.alu_top.A_reg [1]);
	assign _0560_ = _0507_ & ~_0559_;
	assign _0561_ = _0184_ & ~_0509_;
	assign _0562_ = _0561_ | _0560_;
	assign _0563_ = _0558_ & ~_0562_;
	assign _0564_ = ~_0494_;
	assign _0565_ = \mchip.micro_coded_cpu.alu_top.A_reg [0] | ~\mchip.micro_coded_cpu.alu_top.B_reg [0];
	assign _0566_ = \mchip.micro_coded_cpu.alu_top.B_reg [1] ^ \mchip.micro_coded_cpu.alu_top.B_reg [0];
	assign _0567_ = (_0493_ ? \mchip.micro_coded_cpu.alu_top.B_reg [1] : _0566_);
	assign _0568_ = _0567_ ^ \mchip.micro_coded_cpu.alu_top.A_reg [1];
	assign _0569_ = _0568_ ^ _0565_;
	assign _0570_ = _0564_ & ~_0569_;
	assign _0571_ = ~(\mchip.micro_coded_cpu.alu_top.B_reg [1] | \mchip.micro_coded_cpu.alu_top.A_reg [1]);
	assign _0572_ = _0489_ & ~_0571_;
	assign _0573_ = _0572_ | _0570_;
	assign _0574_ = _0563_ & ~_0573_;
	assign \mchip.micro_coded_cpu.alu_top.alu_result_out [1] = _0499_ & ~_0574_;
	assign _0575_ = (\mchip.micro_coded_cpu.alu_top.B_reg [1] ? _0532_ : _0528_);
	assign _0576_ = _0535_ | \mchip.micro_coded_cpu.alu_top.B_reg [1];
	assign _0577_ = (\mchip.micro_coded_cpu.alu_top.B_reg [2] ? _0576_ : _0575_);
	assign _0578_ = _0577_ | \mchip.micro_coded_cpu.alu_top.B_reg [3];
	assign _0579_ = _0578_ | _0539_;
	assign _0580_ = (\mchip.micro_coded_cpu.alu_top.B_reg [0] ? _0524_ : _0526_);
	assign _0581_ = (\mchip.micro_coded_cpu.alu_top.B_reg [1] ? _0517_ : _0580_);
	assign _0582_ = _0581_ | \mchip.micro_coded_cpu.alu_top.B_reg [2];
	assign _0583_ = _0582_ | \mchip.micro_coded_cpu.alu_top.B_reg [3];
	assign _0584_ = _0512_ & ~_0583_;
	assign _0585_ = _0579_ & ~_0584_;
	assign _0586_ = ~(\mchip.micro_coded_cpu.alu_top.B_reg [2] & \mchip.micro_coded_cpu.alu_top.A_reg [2]);
	assign _0587_ = _0507_ & ~_0586_;
	assign _0588_ = _0200_ & ~_0509_;
	assign _0589_ = _0588_ | _0587_;
	assign _0590_ = _0585_ & ~_0589_;
	assign _0591_ = _0565_ & ~_0568_;
	assign _0592_ = \mchip.micro_coded_cpu.alu_top.A_reg [1] & ~_0567_;
	assign _0593_ = _0592_ | _0591_;
	assign _0594_ = \mchip.micro_coded_cpu.alu_top.B_reg [1] | \mchip.micro_coded_cpu.alu_top.B_reg [0];
	assign _0595_ = _0594_ ^ \mchip.micro_coded_cpu.alu_top.B_reg [2];
	assign _0596_ = (_0493_ ? \mchip.micro_coded_cpu.alu_top.B_reg [2] : _0595_);
	assign _0597_ = _0596_ ^ \mchip.micro_coded_cpu.alu_top.A_reg [2];
	assign _0598_ = _0597_ ^ _0593_;
	assign _0599_ = _0564_ & ~_0598_;
	assign _0600_ = ~(\mchip.micro_coded_cpu.alu_top.B_reg [2] | \mchip.micro_coded_cpu.alu_top.A_reg [2]);
	assign _0601_ = _0489_ & ~_0600_;
	assign _0602_ = _0601_ | _0599_;
	assign _0603_ = _0590_ & ~_0602_;
	assign \mchip.micro_coded_cpu.alu_top.alu_result_out [2] = _0499_ & ~_0603_;
	assign _0604_ = (\mchip.micro_coded_cpu.alu_top.B_reg [1] ? _0547_ : _0545_);
	assign _0605_ = _0548_ | \mchip.micro_coded_cpu.alu_top.B_reg [1];
	assign _0606_ = (\mchip.micro_coded_cpu.alu_top.B_reg [2] ? _0605_ : _0604_);
	assign _0607_ = _0606_ | \mchip.micro_coded_cpu.alu_top.B_reg [3];
	assign _0608_ = _0607_ | _0539_;
	assign _0609_ = (\mchip.micro_coded_cpu.alu_top.B_reg [0] ? _0526_ : _0527_);
	assign _0610_ = (\mchip.micro_coded_cpu.alu_top.B_reg [1] ? _0553_ : _0609_);
	assign _0611_ = _0610_ | \mchip.micro_coded_cpu.alu_top.B_reg [2];
	assign _0612_ = _0611_ | \mchip.micro_coded_cpu.alu_top.B_reg [3];
	assign _0613_ = _0512_ & ~_0612_;
	assign _0614_ = _0608_ & ~_0613_;
	assign _0615_ = ~(\mchip.micro_coded_cpu.alu_top.B_reg [3] & \mchip.micro_coded_cpu.alu_top.A_reg [3]);
	assign _0616_ = _0507_ & ~_0615_;
	assign _0617_ = _0192_ & ~_0509_;
	assign _0618_ = _0617_ | _0616_;
	assign _0619_ = _0614_ & ~_0618_;
	assign _0620_ = \mchip.micro_coded_cpu.alu_top.A_reg [2] & ~_0596_;
	assign _0621_ = _0593_ & ~_0597_;
	assign _0622_ = _0621_ | _0620_;
	assign _0623_ = _0523_ & ~_0594_;
	assign _0624_ = _0623_ ^ _0522_;
	assign _0625_ = (_0493_ ? \mchip.micro_coded_cpu.alu_top.B_reg [3] : _0624_);
	assign _0626_ = _0625_ ^ \mchip.micro_coded_cpu.alu_top.A_reg [3];
	assign _0627_ = _0626_ ^ _0622_;
	assign _0628_ = _0564_ & ~_0627_;
	assign _0629_ = ~(\mchip.micro_coded_cpu.alu_top.B_reg [3] | \mchip.micro_coded_cpu.alu_top.A_reg [3]);
	assign _0630_ = _0489_ & ~_0629_;
	assign _0631_ = _0630_ | _0628_;
	assign _0632_ = _0619_ & ~_0631_;
	assign \mchip.micro_coded_cpu.alu_top.alu_result_out [3] = _0499_ & ~_0632_;
	assign _0633_ = _0536_ | \mchip.micro_coded_cpu.alu_top.B_reg [2];
	assign _0634_ = _0633_ | \mchip.micro_coded_cpu.alu_top.B_reg [3];
	assign _0635_ = _0634_ | _0539_;
	assign _0636_ = (\mchip.micro_coded_cpu.alu_top.B_reg [0] ? _0527_ : _0530_);
	assign _0637_ = (\mchip.micro_coded_cpu.alu_top.B_reg [1] ? _0580_ : _0636_);
	assign _0638_ = (\mchip.micro_coded_cpu.alu_top.B_reg [2] ? _0518_ : _0637_);
	assign _0639_ = _0638_ | \mchip.micro_coded_cpu.alu_top.B_reg [3];
	assign _0640_ = _0512_ & ~_0639_;
	assign _0641_ = _0635_ & ~_0640_;
	assign _0642_ = ~(\mchip.micro_coded_cpu.alu_top.B_reg [4] & \mchip.micro_coded_cpu.alu_top.A_reg [4]);
	assign _0643_ = _0507_ & ~_0642_;
	assign _0644_ = _0235_ & ~_0509_;
	assign _0645_ = _0644_ | _0643_;
	assign _0646_ = _0641_ & ~_0645_;
	assign _0647_ = \mchip.micro_coded_cpu.alu_top.A_reg [3] & ~_0625_;
	assign _0648_ = _0620_ & ~_0626_;
	assign _0649_ = _0648_ | _0647_;
	assign _0650_ = _0626_ | _0597_;
	assign _0651_ = _0593_ & ~_0650_;
	assign _0652_ = _0651_ | _0649_;
	assign _0653_ = \mchip.micro_coded_cpu.alu_top.B_reg [2] | \mchip.micro_coded_cpu.alu_top.B_reg [3];
	assign _0654_ = _0653_ | _0594_;
	assign _0655_ = _0654_ ^ \mchip.micro_coded_cpu.alu_top.B_reg [4];
	assign _0656_ = (_0493_ ? \mchip.micro_coded_cpu.alu_top.B_reg [4] : _0655_);
	assign _0657_ = _0656_ ^ \mchip.micro_coded_cpu.alu_top.A_reg [4];
	assign _0658_ = _0657_ ^ _0652_;
	assign _0659_ = _0564_ & ~_0658_;
	assign _0660_ = ~(\mchip.micro_coded_cpu.alu_top.B_reg [4] | \mchip.micro_coded_cpu.alu_top.A_reg [4]);
	assign _0661_ = _0489_ & ~_0660_;
	assign _0662_ = _0661_ | _0659_;
	assign _0663_ = _0646_ & ~_0662_;
	assign \mchip.micro_coded_cpu.alu_top.alu_result_out [4] = _0499_ & ~_0663_;
	assign _0664_ = _0549_ | \mchip.micro_coded_cpu.alu_top.B_reg [2];
	assign _0665_ = _0664_ | \mchip.micro_coded_cpu.alu_top.B_reg [3];
	assign _0666_ = _0665_ | _0539_;
	assign _0667_ = (\mchip.micro_coded_cpu.alu_top.B_reg [0] ? _0530_ : _0531_);
	assign _0668_ = (\mchip.micro_coded_cpu.alu_top.B_reg [1] ? _0609_ : _0667_);
	assign _0669_ = (\mchip.micro_coded_cpu.alu_top.B_reg [2] ? _0554_ : _0668_);
	assign _0670_ = _0669_ | \mchip.micro_coded_cpu.alu_top.B_reg [3];
	assign _0671_ = _0512_ & ~_0670_;
	assign _0672_ = _0666_ & ~_0671_;
	assign _0673_ = ~(\mchip.micro_coded_cpu.alu_top.B_reg [5] & \mchip.micro_coded_cpu.alu_top.A_reg [5]);
	assign _0674_ = _0507_ & ~_0673_;
	assign _0675_ = _0227_ & ~_0509_;
	assign _0676_ = _0675_ | _0674_;
	assign _0677_ = _0672_ & ~_0676_;
	assign _0678_ = \mchip.micro_coded_cpu.alu_top.A_reg [4] & ~_0656_;
	assign _0679_ = _0652_ & ~_0657_;
	assign _0680_ = _0679_ | _0678_;
	assign _0681_ = _0654_ | \mchip.micro_coded_cpu.alu_top.B_reg [4];
	assign _0682_ = _0681_ ^ \mchip.micro_coded_cpu.alu_top.B_reg [5];
	assign _0683_ = (_0493_ ? \mchip.micro_coded_cpu.alu_top.B_reg [5] : _0682_);
	assign _0684_ = _0683_ ^ \mchip.micro_coded_cpu.alu_top.A_reg [5];
	assign _0685_ = _0684_ ^ _0680_;
	assign _0686_ = _0564_ & ~_0685_;
	assign _0687_ = ~(\mchip.micro_coded_cpu.alu_top.B_reg [5] | \mchip.micro_coded_cpu.alu_top.A_reg [5]);
	assign _0688_ = _0489_ & ~_0687_;
	assign _0689_ = _0688_ | _0686_;
	assign _0690_ = _0677_ & ~_0689_;
	assign \mchip.micro_coded_cpu.alu_top.alu_result_out [5] = _0499_ & ~_0690_;
	assign _0691_ = _0576_ | \mchip.micro_coded_cpu.alu_top.B_reg [2];
	assign _0692_ = _0691_ | \mchip.micro_coded_cpu.alu_top.B_reg [3];
	assign _0693_ = _0692_ | _0539_;
	assign _0694_ = (\mchip.micro_coded_cpu.alu_top.B_reg [0] ? _0531_ : _0533_);
	assign _0695_ = (\mchip.micro_coded_cpu.alu_top.B_reg [1] ? _0636_ : _0694_);
	assign _0696_ = (\mchip.micro_coded_cpu.alu_top.B_reg [2] ? _0581_ : _0695_);
	assign _0697_ = _0696_ | \mchip.micro_coded_cpu.alu_top.B_reg [3];
	assign _0698_ = _0512_ & ~_0697_;
	assign _0699_ = _0693_ & ~_0698_;
	assign _0700_ = ~(\mchip.micro_coded_cpu.alu_top.B_reg [6] & \mchip.micro_coded_cpu.alu_top.A_reg [6]);
	assign _0701_ = _0507_ & ~_0700_;
	assign _0702_ = _0218_ & ~_0509_;
	assign _0703_ = _0702_ | _0701_;
	assign _0704_ = _0699_ & ~_0703_;
	assign _0705_ = \mchip.micro_coded_cpu.alu_top.A_reg [5] & ~_0683_;
	assign _0706_ = _0678_ & ~_0684_;
	assign _0707_ = _0706_ | _0705_;
	assign _0708_ = _0684_ | _0657_;
	assign _0709_ = _0652_ & ~_0708_;
	assign _0710_ = _0709_ | _0707_;
	assign _0711_ = ~(_0654_ | _0514_);
	assign _0712_ = ~(_0711_ ^ \mchip.micro_coded_cpu.alu_top.B_reg [6]);
	assign _0713_ = (_0493_ ? \mchip.micro_coded_cpu.alu_top.B_reg [6] : _0712_);
	assign _0714_ = _0713_ ^ \mchip.micro_coded_cpu.alu_top.A_reg [6];
	assign _0715_ = _0714_ ^ _0710_;
	assign _0716_ = _0564_ & ~_0715_;
	assign _0717_ = ~(\mchip.micro_coded_cpu.alu_top.B_reg [6] | \mchip.micro_coded_cpu.alu_top.A_reg [6]);
	assign _0718_ = _0489_ & ~_0717_;
	assign _0719_ = _0718_ | _0716_;
	assign _0720_ = _0704_ & ~_0719_;
	assign \mchip.micro_coded_cpu.alu_top.alu_result_out [6] = _0499_ & ~_0720_;
	assign _0721_ = _0605_ | \mchip.micro_coded_cpu.alu_top.B_reg [2];
	assign _0722_ = _0721_ | \mchip.micro_coded_cpu.alu_top.B_reg [3];
	assign _0723_ = _0722_ | _0539_;
	assign _0724_ = (\mchip.micro_coded_cpu.alu_top.B_reg [0] ? _0533_ : _0534_);
	assign _0725_ = (\mchip.micro_coded_cpu.alu_top.B_reg [1] ? _0667_ : _0724_);
	assign _0726_ = (\mchip.micro_coded_cpu.alu_top.B_reg [2] ? _0610_ : _0725_);
	assign _0727_ = _0726_ | \mchip.micro_coded_cpu.alu_top.B_reg [3];
	assign _0728_ = _0512_ & ~_0727_;
	assign _0729_ = _0723_ & ~_0728_;
	assign _0730_ = ~(\mchip.micro_coded_cpu.alu_top.B_reg [7] & \mchip.micro_coded_cpu.alu_top.A_reg [7]);
	assign _0731_ = _0507_ & ~_0730_;
	assign _0732_ = _0210_ & ~_0509_;
	assign _0733_ = _0732_ | _0731_;
	assign _0734_ = _0729_ & ~_0733_;
	assign _0735_ = _0710_ & ~_0714_;
	assign _0736_ = \mchip.micro_coded_cpu.alu_top.A_reg [6] & ~_0713_;
	assign _0737_ = _0736_ | _0735_;
	assign _0738_ = _0711_ & ~\mchip.micro_coded_cpu.alu_top.B_reg [6];
	assign _0739_ = ~(_0738_ ^ \mchip.micro_coded_cpu.alu_top.B_reg [7]);
	assign _0740_ = (_0493_ ? \mchip.micro_coded_cpu.alu_top.B_reg [7] : _0739_);
	assign _0741_ = _0740_ ^ \mchip.micro_coded_cpu.alu_top.A_reg [7];
	assign _0742_ = _0741_ ^ _0737_;
	assign _0743_ = _0564_ & ~_0742_;
	assign _0744_ = ~(\mchip.micro_coded_cpu.alu_top.B_reg [7] | \mchip.micro_coded_cpu.alu_top.A_reg [7]);
	assign _0745_ = _0489_ & ~_0744_;
	assign _0746_ = _0745_ | _0743_;
	assign _0747_ = _0734_ & ~_0746_;
	assign \mchip.micro_coded_cpu.alu_top.alu_result_out [7] = _0499_ & ~_0747_;
	assign _0748_ = ~(_0043_ & \mchip.micro_coded_cpu.mdecode_reg_top.reg_file_rw );
	assign _0032_ = _0748_ | _0047_;
	assign _0033_ = _0032_ | _0045_;
	assign _0034_ = _0049_ & ~_0033_;
	assign _0035_ = ~(\mchip.micro_coded_cpu.reg_file_interface.reg_sel_in [1] & \mchip.micro_coded_cpu.reg_file_interface.reg_sel_in [0]);
	assign _0029_ = _0034_ & ~_0035_;
	assign \mchip.micro_coded_cpu.load_m_pc_en  = _0246_ | _0071_;
	assign _0036_ = \mchip.micro_coded_cpu.reg_file_interface.reg_sel_in [0] | ~\mchip.micro_coded_cpu.reg_file_interface.reg_sel_in [1];
	assign _0028_ = _0034_ & ~_0036_;
	assign _0037_ = \mchip.micro_coded_cpu.reg_file_interface.reg_sel_in [1] | ~\mchip.micro_coded_cpu.reg_file_interface.reg_sel_in [0];
	assign _0027_ = _0034_ & ~_0037_;
	assign _0038_ = \mchip.micro_coded_cpu.reg_file_interface.reg_sel_in [1] | \mchip.micro_coded_cpu.reg_file_interface.reg_sel_in [0];
	assign _0026_ = _0034_ & ~_0038_;
	assign _0749_[1] = ~(\mchip.micro_coded_cpu.m_inst_to_bit.current_bit_index [1] ^ \mchip.micro_coded_cpu.m_inst_to_bit.current_bit_index [0]);
	assign _0039_ = ~(\mchip.micro_coded_cpu.m_inst_to_bit.current_bit_index [1] | \mchip.micro_coded_cpu.m_inst_to_bit.current_bit_index [0]);
	assign _0749_[2] = _0039_ ^ \mchip.micro_coded_cpu.m_inst_to_bit.current_bit_index [2];
	assign _0040_ = _0039_ & ~\mchip.micro_coded_cpu.m_inst_to_bit.current_bit_index [2];
	assign _0749_[3] = _0040_ ^ \mchip.micro_coded_cpu.m_inst_to_bit.current_bit_index [3];
	reg \mchip.micro_coded_cpu.m_inst_addr_offset_reg[5] ;
	always @(posedge io_in[12]) \mchip.micro_coded_cpu.m_inst_addr_offset_reg[5]  <= _0000_[0];
	assign \mchip.micro_coded_cpu.m_inst_addr_offset [5] = \mchip.micro_coded_cpu.m_inst_addr_offset_reg[5] ;
	reg \mchip.micro_coded_cpu.m_inst_addr_offset_reg[6] ;
	always @(posedge io_in[12]) \mchip.micro_coded_cpu.m_inst_addr_offset_reg[6]  <= _0000_[1];
	assign \mchip.micro_coded_cpu.m_inst_addr_offset [6] = \mchip.micro_coded_cpu.m_inst_addr_offset_reg[6] ;
	reg \mchip.micro_coded_cpu.m_inst_addr_offset_reg[7] ;
	always @(posedge io_in[12]) \mchip.micro_coded_cpu.m_inst_addr_offset_reg[7]  <= _0000_[2];
	assign \mchip.micro_coded_cpu.m_inst_addr_offset [7] = \mchip.micro_coded_cpu.m_inst_addr_offset_reg[7] ;
	reg \mchip.micro_coded_cpu.m_inst_addr_offset_reg[8] ;
	always @(posedge io_in[12]) \mchip.micro_coded_cpu.m_inst_addr_offset_reg[8]  <= _0000_[3];
	assign \mchip.micro_coded_cpu.m_inst_addr_offset [8] = \mchip.micro_coded_cpu.m_inst_addr_offset_reg[8] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.mdecode_reg_top.alu_en_B  <= 1'h0;
		else
			\mchip.micro_coded_cpu.mdecode_reg_top.alu_en_B  <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [8];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [0] <= 1'h0;
		else if (_0030_)
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [0] <= io_in[0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [1] <= 1'h0;
		else if (_0030_)
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [1] <= \mchip.micro_coded_cpu.instr_reg_top.instr_reg [0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [2] <= 1'h0;
		else if (_0030_)
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [2] <= \mchip.micro_coded_cpu.instr_reg_top.instr_reg [1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [3] <= 1'h0;
		else if (_0030_)
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [3] <= \mchip.micro_coded_cpu.instr_reg_top.instr_reg [2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [4] <= 1'h0;
		else if (_0030_)
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [4] <= \mchip.micro_coded_cpu.instr_reg_top.instr_reg [3];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [5] <= 1'h0;
		else if (_0030_)
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [5] <= \mchip.micro_coded_cpu.instr_reg_top.instr_reg [4];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [6] <= 1'h0;
		else if (_0030_)
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [6] <= \mchip.micro_coded_cpu.instr_reg_top.instr_reg [5];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [7] <= 1'h0;
		else if (_0030_)
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [7] <= \mchip.micro_coded_cpu.instr_reg_top.instr_reg [6];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [8] <= 1'h0;
		else if (_0030_)
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [8] <= \mchip.micro_coded_cpu.instr_reg_top.instr_reg [7];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [9] <= 1'h0;
		else if (_0030_)
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [9] <= \mchip.micro_coded_cpu.instr_reg_top.instr_reg [8];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [10] <= 1'h0;
		else if (_0030_)
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [10] <= \mchip.micro_coded_cpu.instr_reg_top.instr_reg [9];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [11] <= 1'h0;
		else if (_0030_)
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [11] <= \mchip.micro_coded_cpu.instr_reg_top.instr_reg [10];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [12] <= 1'h0;
		else if (_0030_)
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [12] <= \mchip.micro_coded_cpu.instr_reg_top.instr_reg [11];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [13] <= 1'h0;
		else if (_0030_)
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [13] <= \mchip.micro_coded_cpu.instr_reg_top.instr_reg [12];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [14] <= 1'h0;
		else if (_0030_)
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [14] <= \mchip.micro_coded_cpu.instr_reg_top.instr_reg [13];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [15] <= 1'h0;
		else if (_0030_)
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [15] <= \mchip.micro_coded_cpu.instr_reg_top.instr_reg [14];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [16] <= 1'h0;
		else if (_0030_)
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [16] <= \mchip.micro_coded_cpu.instr_reg_top.instr_reg [15];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [17] <= 1'h0;
		else if (_0030_)
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [17] <= \mchip.micro_coded_cpu.instr_reg_top.instr_reg [16];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [18] <= 1'h0;
		else if (_0030_)
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [18] <= \mchip.micro_coded_cpu.instr_reg_top.instr_reg [17];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [19] <= 1'h0;
		else if (_0030_)
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [19] <= \mchip.micro_coded_cpu.instr_reg_top.instr_reg [18];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [20] <= 1'h0;
		else if (_0030_)
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [20] <= \mchip.micro_coded_cpu.instr_reg_top.instr_reg [19];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [21] <= 1'h0;
		else if (_0030_)
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [21] <= \mchip.micro_coded_cpu.instr_reg_top.instr_reg [20];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [22] <= 1'h0;
		else if (_0030_)
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [22] <= \mchip.micro_coded_cpu.instr_reg_top.instr_reg [21];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [23] <= 1'h0;
		else if (_0030_)
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [23] <= \mchip.micro_coded_cpu.instr_reg_top.instr_reg [22];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [24] <= 1'h0;
		else if (_0030_)
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [24] <= \mchip.micro_coded_cpu.instr_reg_top.instr_reg [23];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [25] <= 1'h0;
		else if (_0030_)
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [25] <= \mchip.micro_coded_cpu.instr_reg_top.instr_reg [24];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [26] <= 1'h0;
		else if (_0030_)
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [26] <= \mchip.micro_coded_cpu.instr_reg_top.instr_reg [25];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [27] <= 1'h0;
		else if (_0030_)
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [27] <= \mchip.micro_coded_cpu.instr_reg_top.instr_reg [26];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [28] <= 1'h0;
		else if (_0030_)
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [28] <= \mchip.micro_coded_cpu.instr_reg_top.instr_reg [27];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [29] <= 1'h0;
		else if (_0030_)
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [29] <= \mchip.micro_coded_cpu.instr_reg_top.instr_reg [28];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [30] <= 1'h0;
		else if (_0030_)
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [30] <= \mchip.micro_coded_cpu.instr_reg_top.instr_reg [29];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [31] <= 1'h0;
		else if (_0030_)
			\mchip.micro_coded_cpu.instr_reg_top.instr_reg [31] <= \mchip.micro_coded_cpu.instr_reg_top.instr_reg [30];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.m_pc_top.m_pc [0] <= 1'h0;
		else if (\mchip.micro_coded_cpu.load_m_pc_en )
			\mchip.micro_coded_cpu.m_pc_top.m_pc [0] <= \mchip.micro_coded_cpu.m_pc_top.next_m_pc [0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.m_pc_top.m_pc [1] <= 1'h0;
		else if (\mchip.micro_coded_cpu.load_m_pc_en )
			\mchip.micro_coded_cpu.m_pc_top.m_pc [1] <= \mchip.micro_coded_cpu.m_pc_top.next_m_pc [1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.m_pc_top.m_pc [2] <= 1'h0;
		else if (\mchip.micro_coded_cpu.load_m_pc_en )
			\mchip.micro_coded_cpu.m_pc_top.m_pc [2] <= \mchip.micro_coded_cpu.m_pc_top.next_m_pc [2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.m_pc_top.m_pc [3] <= 1'h0;
		else if (\mchip.micro_coded_cpu.load_m_pc_en )
			\mchip.micro_coded_cpu.m_pc_top.m_pc [3] <= \mchip.micro_coded_cpu.m_pc_top.next_m_pc [3];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.m_pc_top.m_pc [4] <= 1'h0;
		else if (\mchip.micro_coded_cpu.load_m_pc_en )
			\mchip.micro_coded_cpu.m_pc_top.m_pc [4] <= \mchip.micro_coded_cpu.m_pc_top.next_m_pc [4];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.m_pc_top.m_pc [5] <= 1'h0;
		else if (\mchip.micro_coded_cpu.load_m_pc_en )
			\mchip.micro_coded_cpu.m_pc_top.m_pc [5] <= \mchip.micro_coded_cpu.m_pc_top.next_m_pc [5];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.m_pc_top.m_pc [6] <= 1'h0;
		else if (\mchip.micro_coded_cpu.load_m_pc_en )
			\mchip.micro_coded_cpu.m_pc_top.m_pc [6] <= \mchip.micro_coded_cpu.m_pc_top.next_m_pc [6];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.m_pc_top.m_pc [7] <= 1'h0;
		else if (\mchip.micro_coded_cpu.load_m_pc_en )
			\mchip.micro_coded_cpu.m_pc_top.m_pc [7] <= \mchip.micro_coded_cpu.m_pc_top.next_m_pc [7];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [0] <= 1'h0;
		else if (_0031_)
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [0] <= io_in[1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [1] <= 1'h0;
		else if (_0031_)
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [1] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [2] <= 1'h0;
		else if (_0031_)
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [2] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [3] <= 1'h0;
		else if (_0031_)
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [3] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [4] <= 1'h0;
		else if (_0031_)
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [4] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [3];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [5] <= 1'h0;
		else if (_0031_)
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [5] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [4];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [6] <= 1'h0;
		else if (_0031_)
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [6] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [5];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [7] <= 1'h0;
		else if (_0031_)
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [7] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [6];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [8] <= 1'h0;
		else if (_0031_)
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [8] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [7];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [9] <= 1'h0;
		else if (_0031_)
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [9] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [8];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [10] <= 1'h0;
		else if (_0031_)
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [10] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [9];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [11] <= 1'h0;
		else if (_0031_)
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [11] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [10];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [12] <= 1'h0;
		else if (_0031_)
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [12] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [11];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [13] <= 1'h0;
		else if (_0031_)
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [13] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [12];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [14] <= 1'h0;
		else if (_0031_)
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [14] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [13];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [15] <= 1'h0;
		else if (_0031_)
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [15] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [14];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [16] <= 1'h0;
		else if (_0031_)
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [16] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [15];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [17] <= 1'h0;
		else if (_0031_)
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [17] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [16];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [18] <= 1'h0;
		else if (_0031_)
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [18] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [17];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [19] <= 1'h0;
		else if (_0031_)
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [19] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [18];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [20] <= 1'h0;
		else if (_0031_)
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [20] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [19];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [21] <= 1'h0;
		else if (_0031_)
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [21] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [20];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [22] <= 1'h0;
		else if (_0031_)
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [22] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [21];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [23] <= 1'h0;
		else if (_0031_)
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [23] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [22];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [24] <= 1'h0;
		else if (_0031_)
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [24] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [23];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [25] <= 1'h0;
		else if (_0031_)
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [25] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [24];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [26] <= 1'h0;
		else if (_0031_)
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [26] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [25];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [27] <= 1'h0;
		else if (_0031_)
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [27] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [26];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [28] <= 1'h0;
		else if (_0031_)
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [28] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [27];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [29] <= 1'h0;
		else if (_0031_)
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [29] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [28];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [30] <= 1'h0;
		else if (_0031_)
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [30] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [29];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [31] <= 1'h0;
		else if (_0031_)
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [31] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [30];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [32] <= 1'h0;
		else if (_0031_)
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [32] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [31];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [33] <= 1'h0;
		else if (_0031_)
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [33] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [32];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [34] <= 1'h0;
		else if (_0031_)
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [34] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [33];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [35] <= 1'h0;
		else if (_0031_)
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [35] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [34];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [36] <= 1'h0;
		else if (_0031_)
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [36] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [35];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [37] <= 1'h0;
		else if (_0031_)
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [37] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [36];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [38] <= 1'h0;
		else if (_0031_)
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [38] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [37];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [39] <= 1'h0;
		else if (_0031_)
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [39] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [38];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [40] <= 1'h0;
		else if (_0031_)
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [40] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [39];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [41] <= 1'h0;
		else if (_0031_)
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [41] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [40];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [42] <= 1'h0;
		else if (_0031_)
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [42] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [41];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [43] <= 1'h0;
		else if (_0031_)
			\mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [43] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [42];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.cpu_fsm_top.current_minst_1 [0] <= 1'h0;
		else if (_0006_)
			\mchip.micro_coded_cpu.cpu_fsm_top.current_minst_1 [0] <= _0012_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.cpu_fsm_top.current_minst_1 [1] <= 1'h0;
		else if (_0006_)
			\mchip.micro_coded_cpu.cpu_fsm_top.current_minst_1 [1] <= _0013_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.cpu_fsm_top.current_minst_1 [2] <= 1'h0;
		else if (_0006_)
			\mchip.micro_coded_cpu.cpu_fsm_top.current_minst_1 [2] <= _0014_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.cpu_fsm_top.current_minst_1 [3] <= 1'h0;
		else if (_0006_)
			\mchip.micro_coded_cpu.cpu_fsm_top.current_minst_1 [3] <= _0015_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.cpu_fsm_top.current_minst_1 [4] <= 1'h0;
		else if (_0006_)
			\mchip.micro_coded_cpu.cpu_fsm_top.current_minst_1 [4] <= _0016_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.cpu_fsm_top.fsm_assist [0] <= 1'h0;
		else if (_0002_)
			\mchip.micro_coded_cpu.cpu_fsm_top.fsm_assist [0] <= _0017_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.cpu_fsm_top.fsm_assist [1] <= 1'h0;
		else if (_0002_)
			\mchip.micro_coded_cpu.cpu_fsm_top.fsm_assist [1] <= _0018_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.cpu_fsm_top.fsm_assist [2] <= 1'h0;
		else if (_0002_)
			\mchip.micro_coded_cpu.cpu_fsm_top.fsm_assist [2] <= _0019_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.cpu_fsm_top.fsm_assist [3] <= 1'h0;
		else if (_0002_)
			\mchip.micro_coded_cpu.cpu_fsm_top.fsm_assist [3] <= _0020_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.cpu_fsm_top.fsm_assist [4] <= 1'h0;
		else if (_0002_)
			\mchip.micro_coded_cpu.cpu_fsm_top.fsm_assist [4] <= _0021_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.cpu_fsm_top.fsm_assist [5] <= 1'h0;
		else if (_0002_)
			\mchip.micro_coded_cpu.cpu_fsm_top.fsm_assist [5] <= _0022_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.reg_file_interface.reg_wr_data_in [0] <= 1'h0;
		else if (_0004_)
			\mchip.micro_coded_cpu.reg_file_interface.reg_wr_data_in [0] <= \mchip.micro_coded_cpu.alu_top.A_bus [0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.reg_file_interface.reg_wr_data_in [1] <= 1'h0;
		else if (_0004_)
			\mchip.micro_coded_cpu.reg_file_interface.reg_wr_data_in [1] <= \mchip.micro_coded_cpu.alu_top.A_bus [1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.reg_file_interface.reg_wr_data_in [2] <= 1'h0;
		else if (_0004_)
			\mchip.micro_coded_cpu.reg_file_interface.reg_wr_data_in [2] <= \mchip.micro_coded_cpu.alu_top.A_bus [2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.reg_file_interface.reg_wr_data_in [3] <= 1'h0;
		else if (_0004_)
			\mchip.micro_coded_cpu.reg_file_interface.reg_wr_data_in [3] <= \mchip.micro_coded_cpu.alu_top.A_bus [3];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.reg_file_interface.reg_wr_data_in [4] <= 1'h0;
		else if (_0004_)
			\mchip.micro_coded_cpu.reg_file_interface.reg_wr_data_in [4] <= \mchip.micro_coded_cpu.alu_top.A_bus [4];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.reg_file_interface.reg_wr_data_in [5] <= 1'h0;
		else if (_0004_)
			\mchip.micro_coded_cpu.reg_file_interface.reg_wr_data_in [5] <= \mchip.micro_coded_cpu.alu_top.A_bus [5];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.reg_file_interface.reg_wr_data_in [6] <= 1'h0;
		else if (_0004_)
			\mchip.micro_coded_cpu.reg_file_interface.reg_wr_data_in [6] <= \mchip.micro_coded_cpu.alu_top.A_bus [6];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.reg_file_interface.reg_wr_data_in [7] <= 1'h0;
		else if (_0004_)
			\mchip.micro_coded_cpu.reg_file_interface.reg_wr_data_in [7] <= \mchip.micro_coded_cpu.alu_top.A_bus [7];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.reg_file_interface.reg_sel_in [0] <= 1'h0;
		else if (_0005_)
			\mchip.micro_coded_cpu.reg_file_interface.reg_sel_in [0] <= \mchip.micro_coded_cpu.alu_top.A_bus [0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.reg_file_interface.reg_sel_in [1] <= 1'h0;
		else if (_0005_)
			\mchip.micro_coded_cpu.reg_file_interface.reg_sel_in [1] <= \mchip.micro_coded_cpu.alu_top.A_bus [1];
	always @(posedge io_in[12])
		if (_0029_)
			\mchip.micro_coded_cpu.reg_file_interface.mreg_file[3] [0] <= \mchip.micro_coded_cpu.reg_file_interface.reg_wr_data_in [0];
	always @(posedge io_in[12])
		if (_0029_)
			\mchip.micro_coded_cpu.reg_file_interface.mreg_file[3] [1] <= \mchip.micro_coded_cpu.reg_file_interface.reg_wr_data_in [1];
	always @(posedge io_in[12])
		if (_0029_)
			\mchip.micro_coded_cpu.reg_file_interface.mreg_file[3] [2] <= \mchip.micro_coded_cpu.reg_file_interface.reg_wr_data_in [2];
	always @(posedge io_in[12])
		if (_0029_)
			\mchip.micro_coded_cpu.reg_file_interface.mreg_file[3] [3] <= \mchip.micro_coded_cpu.reg_file_interface.reg_wr_data_in [3];
	always @(posedge io_in[12])
		if (_0029_)
			\mchip.micro_coded_cpu.reg_file_interface.mreg_file[3] [4] <= \mchip.micro_coded_cpu.reg_file_interface.reg_wr_data_in [4];
	always @(posedge io_in[12])
		if (_0029_)
			\mchip.micro_coded_cpu.reg_file_interface.mreg_file[3] [5] <= \mchip.micro_coded_cpu.reg_file_interface.reg_wr_data_in [5];
	always @(posedge io_in[12])
		if (_0029_)
			\mchip.micro_coded_cpu.reg_file_interface.mreg_file[3] [6] <= \mchip.micro_coded_cpu.reg_file_interface.reg_wr_data_in [6];
	always @(posedge io_in[12])
		if (_0029_)
			\mchip.micro_coded_cpu.reg_file_interface.mreg_file[3] [7] <= \mchip.micro_coded_cpu.reg_file_interface.reg_wr_data_in [7];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.alu_top.B_reg [0] <= 1'h0;
		else if (_0010_)
			\mchip.micro_coded_cpu.alu_top.B_reg [0] <= \mchip.micro_coded_cpu.alu_top.A_bus [0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.alu_top.B_reg [1] <= 1'h0;
		else if (_0010_)
			\mchip.micro_coded_cpu.alu_top.B_reg [1] <= \mchip.micro_coded_cpu.alu_top.A_bus [1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.alu_top.B_reg [2] <= 1'h0;
		else if (_0010_)
			\mchip.micro_coded_cpu.alu_top.B_reg [2] <= \mchip.micro_coded_cpu.alu_top.A_bus [2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.alu_top.B_reg [3] <= 1'h0;
		else if (_0010_)
			\mchip.micro_coded_cpu.alu_top.B_reg [3] <= \mchip.micro_coded_cpu.alu_top.A_bus [3];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.alu_top.B_reg [4] <= 1'h0;
		else if (_0010_)
			\mchip.micro_coded_cpu.alu_top.B_reg [4] <= \mchip.micro_coded_cpu.alu_top.A_bus [4];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.alu_top.B_reg [5] <= 1'h0;
		else if (_0010_)
			\mchip.micro_coded_cpu.alu_top.B_reg [5] <= \mchip.micro_coded_cpu.alu_top.A_bus [5];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.alu_top.B_reg [6] <= 1'h0;
		else if (_0010_)
			\mchip.micro_coded_cpu.alu_top.B_reg [6] <= \mchip.micro_coded_cpu.alu_top.A_bus [6];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.alu_top.B_reg [7] <= 1'h0;
		else if (_0010_)
			\mchip.micro_coded_cpu.alu_top.B_reg [7] <= \mchip.micro_coded_cpu.alu_top.A_bus [7];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.alu_top.A_reg [0] <= 1'h0;
		else if (_0009_)
			\mchip.micro_coded_cpu.alu_top.A_reg [0] <= \mchip.micro_coded_cpu.alu_top.A_bus [0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.alu_top.A_reg [1] <= 1'h0;
		else if (_0009_)
			\mchip.micro_coded_cpu.alu_top.A_reg [1] <= \mchip.micro_coded_cpu.alu_top.A_bus [1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.alu_top.A_reg [2] <= 1'h0;
		else if (_0009_)
			\mchip.micro_coded_cpu.alu_top.A_reg [2] <= \mchip.micro_coded_cpu.alu_top.A_bus [2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.alu_top.A_reg [3] <= 1'h0;
		else if (_0009_)
			\mchip.micro_coded_cpu.alu_top.A_reg [3] <= \mchip.micro_coded_cpu.alu_top.A_bus [3];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.alu_top.A_reg [4] <= 1'h0;
		else if (_0009_)
			\mchip.micro_coded_cpu.alu_top.A_reg [4] <= \mchip.micro_coded_cpu.alu_top.A_bus [4];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.alu_top.A_reg [5] <= 1'h0;
		else if (_0009_)
			\mchip.micro_coded_cpu.alu_top.A_reg [5] <= \mchip.micro_coded_cpu.alu_top.A_bus [5];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.alu_top.A_reg [6] <= 1'h0;
		else if (_0009_)
			\mchip.micro_coded_cpu.alu_top.A_reg [6] <= \mchip.micro_coded_cpu.alu_top.A_bus [6];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.alu_top.A_reg [7] <= 1'h0;
		else if (_0009_)
			\mchip.micro_coded_cpu.alu_top.A_reg [7] <= \mchip.micro_coded_cpu.alu_top.A_bus [7];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.alu_top.alu_result [0] <= 1'h0;
		else if (_0011_)
			\mchip.micro_coded_cpu.alu_top.alu_result [0] <= \mchip.micro_coded_cpu.alu_top.alu_result_out [0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.alu_top.alu_result [1] <= 1'h0;
		else if (_0011_)
			\mchip.micro_coded_cpu.alu_top.alu_result [1] <= \mchip.micro_coded_cpu.alu_top.alu_result_out [1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.alu_top.alu_result [2] <= 1'h0;
		else if (_0011_)
			\mchip.micro_coded_cpu.alu_top.alu_result [2] <= \mchip.micro_coded_cpu.alu_top.alu_result_out [2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.alu_top.alu_result [3] <= 1'h0;
		else if (_0011_)
			\mchip.micro_coded_cpu.alu_top.alu_result [3] <= \mchip.micro_coded_cpu.alu_top.alu_result_out [3];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.alu_top.alu_result [4] <= 1'h0;
		else if (_0011_)
			\mchip.micro_coded_cpu.alu_top.alu_result [4] <= \mchip.micro_coded_cpu.alu_top.alu_result_out [4];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.alu_top.alu_result [5] <= 1'h0;
		else if (_0011_)
			\mchip.micro_coded_cpu.alu_top.alu_result [5] <= \mchip.micro_coded_cpu.alu_top.alu_result_out [5];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.alu_top.alu_result [6] <= 1'h0;
		else if (_0011_)
			\mchip.micro_coded_cpu.alu_top.alu_result [6] <= \mchip.micro_coded_cpu.alu_top.alu_result_out [6];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.alu_top.alu_result [7] <= 1'h0;
		else if (_0011_)
			\mchip.micro_coded_cpu.alu_top.alu_result [7] <= \mchip.micro_coded_cpu.alu_top.alu_result_out [7];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.reg_file_interface.reg_rd_data_out [0] <= 1'h0;
		else if (_0003_)
			\mchip.micro_coded_cpu.reg_file_interface.reg_rd_data_out [0] <= _0001_[0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.reg_file_interface.reg_rd_data_out [1] <= 1'h0;
		else if (_0003_)
			\mchip.micro_coded_cpu.reg_file_interface.reg_rd_data_out [1] <= _0001_[1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.reg_file_interface.reg_rd_data_out [2] <= 1'h0;
		else if (_0003_)
			\mchip.micro_coded_cpu.reg_file_interface.reg_rd_data_out [2] <= _0001_[2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.reg_file_interface.reg_rd_data_out [3] <= 1'h0;
		else if (_0003_)
			\mchip.micro_coded_cpu.reg_file_interface.reg_rd_data_out [3] <= _0001_[3];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.reg_file_interface.reg_rd_data_out [4] <= 1'h0;
		else if (_0003_)
			\mchip.micro_coded_cpu.reg_file_interface.reg_rd_data_out [4] <= _0001_[4];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.reg_file_interface.reg_rd_data_out [5] <= 1'h0;
		else if (_0003_)
			\mchip.micro_coded_cpu.reg_file_interface.reg_rd_data_out [5] <= _0001_[5];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.reg_file_interface.reg_rd_data_out [6] <= 1'h0;
		else if (_0003_)
			\mchip.micro_coded_cpu.reg_file_interface.reg_rd_data_out [6] <= _0001_[6];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.reg_file_interface.reg_rd_data_out [7] <= 1'h0;
		else if (_0003_)
			\mchip.micro_coded_cpu.reg_file_interface.reg_rd_data_out [7] <= _0001_[7];
	always @(posedge io_in[12])
		if (_0028_)
			\mchip.micro_coded_cpu.reg_file_interface.mreg_file[2] [0] <= \mchip.micro_coded_cpu.reg_file_interface.reg_wr_data_in [0];
	always @(posedge io_in[12])
		if (_0028_)
			\mchip.micro_coded_cpu.reg_file_interface.mreg_file[2] [1] <= \mchip.micro_coded_cpu.reg_file_interface.reg_wr_data_in [1];
	always @(posedge io_in[12])
		if (_0028_)
			\mchip.micro_coded_cpu.reg_file_interface.mreg_file[2] [2] <= \mchip.micro_coded_cpu.reg_file_interface.reg_wr_data_in [2];
	always @(posedge io_in[12])
		if (_0028_)
			\mchip.micro_coded_cpu.reg_file_interface.mreg_file[2] [3] <= \mchip.micro_coded_cpu.reg_file_interface.reg_wr_data_in [3];
	always @(posedge io_in[12])
		if (_0028_)
			\mchip.micro_coded_cpu.reg_file_interface.mreg_file[2] [4] <= \mchip.micro_coded_cpu.reg_file_interface.reg_wr_data_in [4];
	always @(posedge io_in[12])
		if (_0028_)
			\mchip.micro_coded_cpu.reg_file_interface.mreg_file[2] [5] <= \mchip.micro_coded_cpu.reg_file_interface.reg_wr_data_in [5];
	always @(posedge io_in[12])
		if (_0028_)
			\mchip.micro_coded_cpu.reg_file_interface.mreg_file[2] [6] <= \mchip.micro_coded_cpu.reg_file_interface.reg_wr_data_in [6];
	always @(posedge io_in[12])
		if (_0028_)
			\mchip.micro_coded_cpu.reg_file_interface.mreg_file[2] [7] <= \mchip.micro_coded_cpu.reg_file_interface.reg_wr_data_in [7];
	always @(posedge io_in[12])
		if (_0027_)
			\mchip.micro_coded_cpu.reg_file_interface.mreg_file[1] [0] <= \mchip.micro_coded_cpu.reg_file_interface.reg_wr_data_in [0];
	always @(posedge io_in[12])
		if (_0027_)
			\mchip.micro_coded_cpu.reg_file_interface.mreg_file[1] [1] <= \mchip.micro_coded_cpu.reg_file_interface.reg_wr_data_in [1];
	always @(posedge io_in[12])
		if (_0027_)
			\mchip.micro_coded_cpu.reg_file_interface.mreg_file[1] [2] <= \mchip.micro_coded_cpu.reg_file_interface.reg_wr_data_in [2];
	always @(posedge io_in[12])
		if (_0027_)
			\mchip.micro_coded_cpu.reg_file_interface.mreg_file[1] [3] <= \mchip.micro_coded_cpu.reg_file_interface.reg_wr_data_in [3];
	always @(posedge io_in[12])
		if (_0027_)
			\mchip.micro_coded_cpu.reg_file_interface.mreg_file[1] [4] <= \mchip.micro_coded_cpu.reg_file_interface.reg_wr_data_in [4];
	always @(posedge io_in[12])
		if (_0027_)
			\mchip.micro_coded_cpu.reg_file_interface.mreg_file[1] [5] <= \mchip.micro_coded_cpu.reg_file_interface.reg_wr_data_in [5];
	always @(posedge io_in[12])
		if (_0027_)
			\mchip.micro_coded_cpu.reg_file_interface.mreg_file[1] [6] <= \mchip.micro_coded_cpu.reg_file_interface.reg_wr_data_in [6];
	always @(posedge io_in[12])
		if (_0027_)
			\mchip.micro_coded_cpu.reg_file_interface.mreg_file[1] [7] <= \mchip.micro_coded_cpu.reg_file_interface.reg_wr_data_in [7];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.mdecode_reg_top.alu_en_A  <= 1'h0;
		else
			\mchip.micro_coded_cpu.mdecode_reg_top.alu_en_A  <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.mdecode_reg_top.reg_file_rw  <= 1'h0;
		else
			\mchip.micro_coded_cpu.mdecode_reg_top.reg_file_rw  <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [5];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.mdecode_reg_top.reg_file_en  <= 1'h0;
		else
			\mchip.micro_coded_cpu.mdecode_reg_top.reg_file_en  <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [4];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.mdecode_reg_top.alu_op [0] <= 1'h0;
		else
			\mchip.micro_coded_cpu.mdecode_reg_top.alu_op [0] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.mdecode_reg_top.alu_op [1] <= 1'h0;
		else
			\mchip.micro_coded_cpu.mdecode_reg_top.alu_op [1] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.mdecode_reg_top.alu_op [2] <= 1'h0;
		else
			\mchip.micro_coded_cpu.mdecode_reg_top.alu_op [2] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [3];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.mdecode_reg_top.is_imm_active  <= 1'h0;
		else
			\mchip.micro_coded_cpu.mdecode_reg_top.is_imm_active  <= \mchip.micro_coded_cpu.mdecode_reg_top.is_imm_active_md ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.mdecode_reg_top.imm [0] <= 1'h0;
		else
			\mchip.micro_coded_cpu.mdecode_reg_top.imm [0] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [20];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.mdecode_reg_top.imm [1] <= 1'h0;
		else
			\mchip.micro_coded_cpu.mdecode_reg_top.imm [1] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [21];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.mdecode_reg_top.imm [2] <= 1'h0;
		else
			\mchip.micro_coded_cpu.mdecode_reg_top.imm [2] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [22];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.mdecode_reg_top.imm [3] <= 1'h0;
		else
			\mchip.micro_coded_cpu.mdecode_reg_top.imm [3] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [23];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.mdecode_reg_top.imm [4] <= 1'h0;
		else
			\mchip.micro_coded_cpu.mdecode_reg_top.imm [4] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [24];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.mdecode_reg_top.imm [5] <= 1'h0;
		else
			\mchip.micro_coded_cpu.mdecode_reg_top.imm [5] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [25];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.mdecode_reg_top.imm [6] <= 1'h0;
		else
			\mchip.micro_coded_cpu.mdecode_reg_top.imm [6] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [26];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.mdecode_reg_top.imm [7] <= 1'h0;
		else
			\mchip.micro_coded_cpu.mdecode_reg_top.imm [7] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [27];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.mdecode_reg_top.reg_src [0] <= 1'h0;
		else
			\mchip.micro_coded_cpu.mdecode_reg_top.reg_src [0] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [36];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.mdecode_reg_top.reg_src [1] <= 1'h0;
		else
			\mchip.micro_coded_cpu.mdecode_reg_top.reg_src [1] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [37];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.mdecode_reg_top.reg_src [2] <= 1'h0;
		else
			\mchip.micro_coded_cpu.mdecode_reg_top.reg_src [2] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [38];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.mdecode_reg_top.reg_src [3] <= 1'h0;
		else
			\mchip.micro_coded_cpu.mdecode_reg_top.reg_src [3] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [39];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.mdecode_reg_top.reg_src [4] <= 1'h0;
		else
			\mchip.micro_coded_cpu.mdecode_reg_top.reg_src [4] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [40];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.mdecode_reg_top.reg_dst [0] <= 1'h0;
		else
			\mchip.micro_coded_cpu.mdecode_reg_top.reg_dst [0] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [31];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.mdecode_reg_top.reg_dst [1] <= 1'h0;
		else
			\mchip.micro_coded_cpu.mdecode_reg_top.reg_dst [1] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [32];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.mdecode_reg_top.reg_dst [2] <= 1'h0;
		else
			\mchip.micro_coded_cpu.mdecode_reg_top.reg_dst [2] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [33];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.mdecode_reg_top.reg_dst [3] <= 1'h0;
		else
			\mchip.micro_coded_cpu.mdecode_reg_top.reg_dst [3] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [34];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.mdecode_reg_top.reg_dst [4] <= 1'h0;
		else
			\mchip.micro_coded_cpu.mdecode_reg_top.reg_dst [4] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [35];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.mdecode_reg_top.mbranch_target [0] <= 1'h0;
		else
			\mchip.micro_coded_cpu.mdecode_reg_top.mbranch_target [0] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [10];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.mdecode_reg_top.mbranch_target [1] <= 1'h0;
		else
			\mchip.micro_coded_cpu.mdecode_reg_top.mbranch_target [1] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [11];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.mdecode_reg_top.mbranch_target [2] <= 1'h0;
		else
			\mchip.micro_coded_cpu.mdecode_reg_top.mbranch_target [2] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [12];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.mdecode_reg_top.mbranch_target [3] <= 1'h0;
		else
			\mchip.micro_coded_cpu.mdecode_reg_top.mbranch_target [3] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [13];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.mdecode_reg_top.mbranch_target [4] <= 1'h0;
		else
			\mchip.micro_coded_cpu.mdecode_reg_top.mbranch_target [4] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [14];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.mdecode_reg_top.mbranch_target [5] <= 1'h0;
		else
			\mchip.micro_coded_cpu.mdecode_reg_top.mbranch_target [5] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [15];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.mdecode_reg_top.mbranch_target [6] <= 1'h0;
		else
			\mchip.micro_coded_cpu.mdecode_reg_top.mbranch_target [6] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [16];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.mdecode_reg_top.mbranch_target [7] <= 1'h0;
		else
			\mchip.micro_coded_cpu.mdecode_reg_top.mbranch_target [7] <= \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [17];
	always @(posedge io_in[12])
		if (_0008_)
			\mchip.micro_coded_cpu.m_inst_to_bit.current_bit_index [0] <= 1'h0;
		else
			\mchip.micro_coded_cpu.m_inst_to_bit.current_bit_index [0] <= _0749_[0];
	always @(posedge io_in[12])
		if (_0008_)
			\mchip.micro_coded_cpu.m_inst_to_bit.current_bit_index [1] <= 1'h0;
		else
			\mchip.micro_coded_cpu.m_inst_to_bit.current_bit_index [1] <= _0749_[1];
	always @(posedge io_in[12])
		if (_0008_)
			\mchip.micro_coded_cpu.m_inst_to_bit.current_bit_index [2] <= 1'h0;
		else
			\mchip.micro_coded_cpu.m_inst_to_bit.current_bit_index [2] <= _0749_[2];
	always @(posedge io_in[12])
		if (_0008_)
			\mchip.micro_coded_cpu.m_inst_to_bit.current_bit_index [3] <= 1'h1;
		else
			\mchip.micro_coded_cpu.m_inst_to_bit.current_bit_index [3] <= _0749_[3];
	always @(posedge io_in[12])
		if (_0026_)
			\mchip.micro_coded_cpu.reg_file_interface.mreg_file[0] [0] <= \mchip.micro_coded_cpu.reg_file_interface.reg_wr_data_in [0];
	always @(posedge io_in[12])
		if (_0026_)
			\mchip.micro_coded_cpu.reg_file_interface.mreg_file[0] [1] <= \mchip.micro_coded_cpu.reg_file_interface.reg_wr_data_in [1];
	always @(posedge io_in[12])
		if (_0026_)
			\mchip.micro_coded_cpu.reg_file_interface.mreg_file[0] [2] <= \mchip.micro_coded_cpu.reg_file_interface.reg_wr_data_in [2];
	always @(posedge io_in[12])
		if (_0026_)
			\mchip.micro_coded_cpu.reg_file_interface.mreg_file[0] [3] <= \mchip.micro_coded_cpu.reg_file_interface.reg_wr_data_in [3];
	always @(posedge io_in[12])
		if (_0026_)
			\mchip.micro_coded_cpu.reg_file_interface.mreg_file[0] [4] <= \mchip.micro_coded_cpu.reg_file_interface.reg_wr_data_in [4];
	always @(posedge io_in[12])
		if (_0026_)
			\mchip.micro_coded_cpu.reg_file_interface.mreg_file[0] [5] <= \mchip.micro_coded_cpu.reg_file_interface.reg_wr_data_in [5];
	always @(posedge io_in[12])
		if (_0026_)
			\mchip.micro_coded_cpu.reg_file_interface.mreg_file[0] [6] <= \mchip.micro_coded_cpu.reg_file_interface.reg_wr_data_in [6];
	always @(posedge io_in[12])
		if (_0026_)
			\mchip.micro_coded_cpu.reg_file_interface.mreg_file[0] [7] <= \mchip.micro_coded_cpu.reg_file_interface.reg_wr_data_in [7];
	reg \mchip.micro_coded_cpu.cpu_fsm_top.cpu_state_reg[0] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.cpu_fsm_top.cpu_state_reg[0]  <= 1'h0;
		else if (_0007_)
			\mchip.micro_coded_cpu.cpu_fsm_top.cpu_state_reg[0]  <= _0023_;
	assign \mchip.micro_coded_cpu.cpu_fsm_top.cpu_state [0] = \mchip.micro_coded_cpu.cpu_fsm_top.cpu_state_reg[0] ;
	reg \mchip.micro_coded_cpu.cpu_fsm_top.cpu_state_reg[1] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.cpu_fsm_top.cpu_state_reg[1]  <= 1'h0;
		else if (_0007_)
			\mchip.micro_coded_cpu.cpu_fsm_top.cpu_state_reg[1]  <= _0024_;
	assign \mchip.micro_coded_cpu.cpu_fsm_top.cpu_state [1] = \mchip.micro_coded_cpu.cpu_fsm_top.cpu_state_reg[1] ;
	reg \mchip.micro_coded_cpu.cpu_fsm_top.cpu_state_reg[2] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.micro_coded_cpu.cpu_fsm_top.cpu_state_reg[2]  <= 1'h0;
		else if (_0007_)
			\mchip.micro_coded_cpu.cpu_fsm_top.cpu_state_reg[2]  <= _0025_;
	assign \mchip.micro_coded_cpu.cpu_fsm_top.cpu_state [2] = \mchip.micro_coded_cpu.cpu_fsm_top.cpu_state_reg[2] ;
	assign io_out = {9'h000, \mchip.micro_coded_cpu.cpu_fsm_top.cpu_state [2:0], \mchip.micro_coded_cpu.m_inst_addr_stream , 1'h0};
	assign \mchip.clock  = io_in[12];
	assign \mchip.io_in  = io_in[11:0];
	assign \mchip.io_out  = {7'h00, \mchip.micro_coded_cpu.cpu_fsm_top.cpu_state [2:0], \mchip.micro_coded_cpu.m_inst_addr_stream , 1'h0};
	assign \mchip.micro_coded_cpu.A_reg  = \mchip.micro_coded_cpu.alu_top.A_reg ;
	assign \mchip.micro_coded_cpu.B_Reg  = 1'h0;
	assign \mchip.micro_coded_cpu.B_reg  = \mchip.micro_coded_cpu.alu_top.B_reg ;
	assign \mchip.micro_coded_cpu.alu_en_A  = \mchip.micro_coded_cpu.mdecode_reg_top.alu_en_A ;
	assign \mchip.micro_coded_cpu.alu_en_A_md  = \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [0];
	assign \mchip.micro_coded_cpu.alu_en_B  = \mchip.micro_coded_cpu.mdecode_reg_top.alu_en_B ;
	assign \mchip.micro_coded_cpu.alu_en_B_md  = \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [8];
	assign \mchip.micro_coded_cpu.alu_op  = \mchip.micro_coded_cpu.mdecode_reg_top.alu_op ;
	assign \mchip.micro_coded_cpu.alu_op_md  = \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [3:1];
	assign \mchip.micro_coded_cpu.alu_result  = \mchip.micro_coded_cpu.alu_top.alu_result ;
	assign \mchip.micro_coded_cpu.alu_top.B_bus  = \mchip.micro_coded_cpu.alu_top.A_bus ;
	assign \mchip.micro_coded_cpu.alu_top.alu.A  = \mchip.micro_coded_cpu.alu_top.A_reg ;
	assign \mchip.micro_coded_cpu.alu_top.alu.B  = \mchip.micro_coded_cpu.alu_top.B_reg ;
	assign \mchip.micro_coded_cpu.alu_top.alu.a_equal_b  = 1'h0;
	assign \mchip.micro_coded_cpu.alu_top.alu.a_greater_b  = 1'h0;
	assign \mchip.micro_coded_cpu.alu_top.alu.alu_op  = \mchip.micro_coded_cpu.mdecode_reg_top.alu_op ;
	assign \mchip.micro_coded_cpu.alu_top.alu.alu_result  = \mchip.micro_coded_cpu.alu_top.alu_result_out ;
	assign \mchip.micro_coded_cpu.alu_top.alu.alu_result_tmp  = \mchip.micro_coded_cpu.alu_top.alu_result_out ;
	assign \mchip.micro_coded_cpu.alu_top.alu.carry_in  = 1'h0;
	assign \mchip.micro_coded_cpu.alu_top.alu.equal  = 1'h0;
	assign \mchip.micro_coded_cpu.alu_top.alu.greater  = 1'h0;
	assign \mchip.micro_coded_cpu.alu_top.alu.zero  = 8'h00;
	assign \mchip.micro_coded_cpu.alu_top.alu_en_A_reg  = \mchip.micro_coded_cpu.mdecode_reg_top.alu_en_A ;
	assign \mchip.micro_coded_cpu.alu_top.alu_en_B_reg  = \mchip.micro_coded_cpu.mdecode_reg_top.alu_en_B ;
	assign \mchip.micro_coded_cpu.alu_top.alu_op  = \mchip.micro_coded_cpu.mdecode_reg_top.alu_op ;
	assign \mchip.micro_coded_cpu.alu_top.carry_in  = 1'h0;
	assign \mchip.micro_coded_cpu.alu_top.cc_equal  = 1'h0;
	assign \mchip.micro_coded_cpu.alu_top.cc_equal_out  = 1'h0;
	assign \mchip.micro_coded_cpu.alu_top.cc_greater  = 1'h0;
	assign \mchip.micro_coded_cpu.alu_top.cc_greater_out  = 1'h0;
	assign \mchip.micro_coded_cpu.alu_top.cpu_state  = {1'h0, \mchip.micro_coded_cpu.cpu_fsm_top.cpu_state [2:0]};
	assign \mchip.micro_coded_cpu.alu_top.sys_clk  = io_in[12];
	assign \mchip.micro_coded_cpu.alu_top.sys_reset  = io_in[13];
	assign \mchip.micro_coded_cpu.branch_target_id  = \mchip.micro_coded_cpu.instr_reg_top.instr_reg [7:0];
	assign \mchip.micro_coded_cpu.cc_equal  = 1'h0;
	assign \mchip.micro_coded_cpu.cc_greater  = 1'h0;
	assign \mchip.micro_coded_cpu.cpu_fsm_top.cpu_state [3] = 1'h0;
	assign \mchip.micro_coded_cpu.cpu_fsm_top.is_micro_nop  = 1'h0;
	assign \mchip.micro_coded_cpu.cpu_fsm_top.is_nop  = 1'h0;
	assign \mchip.micro_coded_cpu.cpu_fsm_top.sys_clk  = io_in[12];
	assign \mchip.micro_coded_cpu.cpu_fsm_top.sys_reset  = io_in[13];
	assign \mchip.micro_coded_cpu.cpu_state  = {1'h0, \mchip.micro_coded_cpu.cpu_fsm_top.cpu_state [2:0]};
	assign \mchip.micro_coded_cpu.imm  = \mchip.micro_coded_cpu.mdecode_reg_top.imm ;
	assign \mchip.micro_coded_cpu.imm_id  = \mchip.micro_coded_cpu.instr_reg_top.instr_reg [7:0];
	assign \mchip.micro_coded_cpu.imm_md  = \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [27:20];
	assign \mchip.micro_coded_cpu.inst_addr_stream  = 1'h0;
	assign \mchip.micro_coded_cpu.inst_to_bit.cpu_state  = {1'h0, \mchip.micro_coded_cpu.cpu_fsm_top.cpu_state [2:0]};
	assign \mchip.micro_coded_cpu.inst_to_bit.inst_addr  = 8'h00;
	assign \mchip.micro_coded_cpu.inst_to_bit.inst_addr_stream  = 1'h0;
	assign \mchip.micro_coded_cpu.inst_to_bit.sys_clk  = io_in[12];
	assign \mchip.micro_coded_cpu.inst_to_bit.sys_reset  = io_in[13];
	assign \mchip.micro_coded_cpu.inst_type  = \mchip.micro_coded_cpu.instr_reg_top.instr_reg [31:27];
	assign \mchip.micro_coded_cpu.instr_in  = io_in[0];
	assign \mchip.micro_coded_cpu.instr_reg  = \mchip.micro_coded_cpu.instr_reg_top.instr_reg ;
	assign \mchip.micro_coded_cpu.instr_reg_top.instr_in  = io_in[0];
	assign \mchip.micro_coded_cpu.instr_reg_top.sys_clk  = io_in[12];
	assign \mchip.micro_coded_cpu.instr_reg_top.sys_reset  = io_in[13];
	assign \mchip.micro_coded_cpu.ir_decode_top.branch_target_id  = \mchip.micro_coded_cpu.instr_reg_top.instr_reg [7:0];
	assign \mchip.micro_coded_cpu.ir_decode_top.imm_id  = \mchip.micro_coded_cpu.instr_reg_top.instr_reg [7:0];
	assign \mchip.micro_coded_cpu.ir_decode_top.inst_type  = \mchip.micro_coded_cpu.instr_reg_top.instr_reg [31:27];
	assign \mchip.micro_coded_cpu.ir_decode_top.instr_in  = \mchip.micro_coded_cpu.instr_reg_top.instr_reg ;
	assign \mchip.micro_coded_cpu.ir_decode_top.is_imm_active_id  = \mchip.micro_coded_cpu.instr_reg_top.instr_reg [26];
	assign \mchip.micro_coded_cpu.ir_decode_top.reg_dst_id  = \mchip.micro_coded_cpu.instr_reg_top.instr_reg [25:22];
	assign \mchip.micro_coded_cpu.ir_decode_top.reg_src_1_id  = \mchip.micro_coded_cpu.instr_reg_top.instr_reg [21:18];
	assign \mchip.micro_coded_cpu.ir_decode_top.reg_src_2_id  = \mchip.micro_coded_cpu.instr_reg_top.instr_reg [17:14];
	assign \mchip.micro_coded_cpu.is_current_inst_nop  = 1'h0;
	assign \mchip.micro_coded_cpu.is_current_micro_inst_nop  = 1'h0;
	assign \mchip.micro_coded_cpu.is_imm_active  = \mchip.micro_coded_cpu.mdecode_reg_top.is_imm_active ;
	assign \mchip.micro_coded_cpu.is_imm_active_id  = \mchip.micro_coded_cpu.instr_reg_top.instr_reg [26];
	assign \mchip.micro_coded_cpu.is_imm_active_md  = \mchip.micro_coded_cpu.mdecode_reg_top.is_imm_active_md ;
	assign \mchip.micro_coded_cpu.load_pc_en  = 1'h0;
	assign \mchip.micro_coded_cpu.m_inst_addr_offset [4:0] = 5'h00;
	assign \mchip.micro_coded_cpu.m_inst_addr_offset_gen.instr_in  = \mchip.micro_coded_cpu.instr_reg_top.instr_reg ;
	assign \mchip.micro_coded_cpu.m_inst_addr_offset_gen.instr_type  = \mchip.micro_coded_cpu.instr_reg_top.instr_reg [31:27];
	assign \mchip.micro_coded_cpu.m_inst_addr_offset_gen.m_inst_addr_base  = {\mchip.micro_coded_cpu.m_inst_addr_offset [8:5], 5'h00};
	assign \mchip.micro_coded_cpu.m_inst_addr_offset_gen.offset  = {\mchip.micro_coded_cpu.m_inst_addr_offset [8:5], 5'h00};
	assign \mchip.micro_coded_cpu.m_inst_decode_top.alu_en_A_md  = \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [0];
	assign \mchip.micro_coded_cpu.m_inst_decode_top.alu_en_B_md  = \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [8];
	assign \mchip.micro_coded_cpu.m_inst_decode_top.alu_op_md  = \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [3:1];
	assign \mchip.micro_coded_cpu.m_inst_decode_top.imm_md  = \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [27:20];
	assign \mchip.micro_coded_cpu.m_inst_decode_top.is_imm_active_md  = \mchip.micro_coded_cpu.mdecode_reg_top.is_imm_active_md ;
	assign \mchip.micro_coded_cpu.m_inst_decode_top.m_args  = \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [9:0];
	assign \mchip.micro_coded_cpu.m_inst_decode_top.mbranch_target_md  = \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [17:10];
	assign \mchip.micro_coded_cpu.m_inst_decode_top.minstr_in  = \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg ;
	assign \mchip.micro_coded_cpu.m_inst_decode_top.minstr_type  = \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [43:41];
	assign \mchip.micro_coded_cpu.m_inst_decode_top.reg_dst_md  = \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [35:31];
	assign \mchip.micro_coded_cpu.m_inst_decode_top.reg_file_en_md  = \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [4];
	assign \mchip.micro_coded_cpu.m_inst_decode_top.reg_file_rw_md  = \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [5];
	assign \mchip.micro_coded_cpu.m_inst_decode_top.reg_src_md  = \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [40:36];
	assign \mchip.micro_coded_cpu.m_inst_to_bit.cpu_state  = {1'h0, \mchip.micro_coded_cpu.cpu_fsm_top.cpu_state [2:0]};
	assign \mchip.micro_coded_cpu.m_inst_to_bit.m_inst_addr  = {4'h0, \mchip.micro_coded_cpu.m_pc_top.m_pc [4:0]};
	assign \mchip.micro_coded_cpu.m_inst_to_bit.m_inst_addr_stream  = \mchip.micro_coded_cpu.m_inst_addr_stream ;
	assign \mchip.micro_coded_cpu.m_inst_to_bit.sys_clk  = io_in[12];
	assign \mchip.micro_coded_cpu.m_inst_to_bit.sys_reset  = io_in[13];
	assign \mchip.micro_coded_cpu.m_instr_in  = io_in[1];
	assign \mchip.micro_coded_cpu.m_instr_reg  = \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg ;
	assign \mchip.micro_coded_cpu.m_instr_reg_top.minstr_in  = io_in[1];
	assign \mchip.micro_coded_cpu.m_instr_reg_top.sys_clk  = io_in[12];
	assign \mchip.micro_coded_cpu.m_instr_reg_top.sys_reset  = io_in[13];
	assign \mchip.micro_coded_cpu.m_pc  = \mchip.micro_coded_cpu.m_pc_top.m_pc ;
	assign \mchip.micro_coded_cpu.m_pc_top.load_m_pc_en  = \mchip.micro_coded_cpu.load_m_pc_en ;
	assign \mchip.micro_coded_cpu.m_pc_top.sys_clk  = io_in[12];
	assign \mchip.micro_coded_cpu.m_pc_top.sys_reset  = io_in[13];
	assign \mchip.micro_coded_cpu.mbranch_target  = \mchip.micro_coded_cpu.mdecode_reg_top.mbranch_target ;
	assign \mchip.micro_coded_cpu.mbranch_target_md  = \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [17:10];
	assign \mchip.micro_coded_cpu.mdecode_reg_top.alu_en_A_md  = \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [0];
	assign \mchip.micro_coded_cpu.mdecode_reg_top.alu_en_B_md  = \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [8];
	assign \mchip.micro_coded_cpu.mdecode_reg_top.alu_op_md  = \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [3:1];
	assign \mchip.micro_coded_cpu.mdecode_reg_top.imm_md  = \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [27:20];
	assign \mchip.micro_coded_cpu.mdecode_reg_top.mbranch_target_md  = \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [17:10];
	assign \mchip.micro_coded_cpu.mdecode_reg_top.reg_dst_md  = \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [35:31];
	assign \mchip.micro_coded_cpu.mdecode_reg_top.reg_file_en_md  = \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [4];
	assign \mchip.micro_coded_cpu.mdecode_reg_top.reg_file_rw_md  = \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [5];
	assign \mchip.micro_coded_cpu.mdecode_reg_top.reg_src_md  = \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [40:36];
	assign \mchip.micro_coded_cpu.mdecode_reg_top.sys_clk  = io_in[12];
	assign \mchip.micro_coded_cpu.mdecode_reg_top.sys_reset  = io_in[13];
	assign \mchip.micro_coded_cpu.minstr_type  = \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [43:41];
	assign \mchip.micro_coded_cpu.mpc_offset  = {4'h0, \mchip.micro_coded_cpu.m_pc_top.m_pc [4:0]};
	assign \mchip.micro_coded_cpu.next_m_pc  = \mchip.micro_coded_cpu.m_pc_top.next_m_pc ;
	assign \mchip.micro_coded_cpu.pc  = 8'h00;
	assign \mchip.micro_coded_cpu.pc_top.load_pc_en  = 1'h0;
	assign \mchip.micro_coded_cpu.pc_top.pc  = 8'h00;
	assign \mchip.micro_coded_cpu.pc_top.sys_clk  = io_in[12];
	assign \mchip.micro_coded_cpu.pc_top.sys_reset  = io_in[13];
	assign \mchip.micro_coded_cpu.reg_dst  = \mchip.micro_coded_cpu.mdecode_reg_top.reg_dst ;
	assign \mchip.micro_coded_cpu.reg_dst_id  = \mchip.micro_coded_cpu.instr_reg_top.instr_reg [25:22];
	assign \mchip.micro_coded_cpu.reg_dst_md  = \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [35:31];
	assign \mchip.micro_coded_cpu.reg_file_en  = \mchip.micro_coded_cpu.mdecode_reg_top.reg_file_en ;
	assign \mchip.micro_coded_cpu.reg_file_en_md  = \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [4];
	assign \mchip.micro_coded_cpu.reg_file_interface.cpu_state  = {1'h0, \mchip.micro_coded_cpu.cpu_fsm_top.cpu_state [2:0]};
	assign \mchip.micro_coded_cpu.reg_file_interface.reg_dst  = \mchip.micro_coded_cpu.instr_reg_top.instr_reg [25:22];
	assign \mchip.micro_coded_cpu.reg_file_interface.reg_file_en  = \mchip.micro_coded_cpu.mdecode_reg_top.reg_file_en ;
	assign \mchip.micro_coded_cpu.reg_file_interface.reg_file_rw  = \mchip.micro_coded_cpu.mdecode_reg_top.reg_file_rw ;
	assign \mchip.micro_coded_cpu.reg_file_interface.reg_rd_data  = \mchip.micro_coded_cpu.reg_file_interface.reg_rd_data_out ;
	assign \mchip.micro_coded_cpu.reg_file_interface.shared_write_bus  = \mchip.micro_coded_cpu.alu_top.A_bus ;
	assign \mchip.micro_coded_cpu.reg_file_interface.sys_clk  = io_in[12];
	assign \mchip.micro_coded_cpu.reg_file_interface.sys_reset  = io_in[13];
	assign \mchip.micro_coded_cpu.reg_file_rw  = \mchip.micro_coded_cpu.mdecode_reg_top.reg_file_rw ;
	assign \mchip.micro_coded_cpu.reg_file_rw_md  = \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [5];
	assign \mchip.micro_coded_cpu.reg_rd_data  = \mchip.micro_coded_cpu.reg_file_interface.reg_rd_data_out ;
	assign \mchip.micro_coded_cpu.reg_src  = \mchip.micro_coded_cpu.mdecode_reg_top.reg_src ;
	assign \mchip.micro_coded_cpu.reg_src_1_id  = \mchip.micro_coded_cpu.instr_reg_top.instr_reg [21:18];
	assign \mchip.micro_coded_cpu.reg_src_2_id  = \mchip.micro_coded_cpu.instr_reg_top.instr_reg [17:14];
	assign \mchip.micro_coded_cpu.reg_src_dst_cmp_branch.A  = \mchip.micro_coded_cpu.alu_top.A_reg ;
	assign \mchip.micro_coded_cpu.reg_src_dst_cmp_branch.B  = 8'h00;
	assign \mchip.micro_coded_cpu.reg_src_dst_cmp_branch.alu_result  = \mchip.micro_coded_cpu.alu_top.alu_result ;
	assign \mchip.micro_coded_cpu.reg_src_dst_cmp_branch.cc_equal  = 1'h0;
	assign \mchip.micro_coded_cpu.reg_src_dst_cmp_branch.cc_greater  = 1'h0;
	assign \mchip.micro_coded_cpu.reg_src_dst_cmp_branch.imm  = \mchip.micro_coded_cpu.mdecode_reg_top.imm ;
	assign \mchip.micro_coded_cpu.reg_src_dst_cmp_branch.is_imm_active  = \mchip.micro_coded_cpu.mdecode_reg_top.is_imm_active ;
	assign \mchip.micro_coded_cpu.reg_src_dst_cmp_branch.reg_dst  = \mchip.micro_coded_cpu.mdecode_reg_top.reg_dst ;
	assign \mchip.micro_coded_cpu.reg_src_md  = \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [40:36];
	assign \mchip.micro_coded_cpu.shared_mcpu_bus.alu_result  = \mchip.micro_coded_cpu.alu_top.alu_result ;
	assign \mchip.micro_coded_cpu.shared_mcpu_bus.cc_equal  = 1'h0;
	assign \mchip.micro_coded_cpu.shared_mcpu_bus.cc_greater  = 1'h0;
	assign \mchip.micro_coded_cpu.shared_mcpu_bus.imm  = \mchip.micro_coded_cpu.mdecode_reg_top.imm ;
	assign \mchip.micro_coded_cpu.shared_mcpu_bus.m_pc  = \mchip.micro_coded_cpu.m_pc_top.m_pc ;
	assign \mchip.micro_coded_cpu.shared_mcpu_bus.mbranch_target  = \mchip.micro_coded_cpu.mdecode_reg_top.mbranch_target ;
	assign \mchip.micro_coded_cpu.shared_mcpu_bus.minstr_type  = \mchip.micro_coded_cpu.m_instr_reg_top.m_instr_reg [43:41];
	assign \mchip.micro_coded_cpu.shared_mcpu_bus.reg_dst  = \mchip.micro_coded_cpu.mdecode_reg_top.reg_dst ;
	assign \mchip.micro_coded_cpu.shared_mcpu_bus.reg_rd_data  = \mchip.micro_coded_cpu.reg_file_interface.reg_rd_data_out ;
	assign \mchip.micro_coded_cpu.shared_mcpu_bus.reg_src  = \mchip.micro_coded_cpu.mdecode_reg_top.reg_src ;
	assign \mchip.micro_coded_cpu.shared_mcpu_bus.rs1  = \mchip.micro_coded_cpu.instr_reg_top.instr_reg [19:18];
	assign \mchip.micro_coded_cpu.shared_mcpu_bus.rs2  = \mchip.micro_coded_cpu.instr_reg_top.instr_reg [15:14];
	assign \mchip.micro_coded_cpu.shared_mcpu_bus.write_bus_out  = \mchip.micro_coded_cpu.alu_top.A_bus ;
	assign \mchip.micro_coded_cpu.shared_write_bus  = \mchip.micro_coded_cpu.alu_top.A_bus ;
	assign \mchip.micro_coded_cpu.sys_clk  = io_in[12];
	assign \mchip.micro_coded_cpu.sys_reset  = io_in[13];
	assign \mchip.reset  = io_in[13];
endmodule
module d29_bwilhelm_i8008 (
	io_in,
	io_out
);
	reg [2:0] _0000_;
	wire _0001_;
	wire _0002_;
	wire _0003_;
	wire _0004_;
	wire _0005_;
	wire _0006_;
	wire _0007_;
	wire _0008_;
	wire _0009_;
	wire _0010_;
	wire _0011_;
	wire _0012_;
	wire _0013_;
	wire _0014_;
	wire _0015_;
	wire _0016_;
	wire _0017_;
	wire _0018_;
	wire _0019_;
	wire _0020_;
	wire _0021_;
	wire _0022_;
	wire _0023_;
	wire _0024_;
	wire _0025_;
	wire _0026_;
	wire _0027_;
	wire _0028_;
	wire _0029_;
	wire _0030_;
	wire _0031_;
	wire _0032_;
	wire _0033_;
	wire _0034_;
	wire _0035_;
	wire _0036_;
	wire _0037_;
	wire _0038_;
	wire _0039_;
	wire _0040_;
	wire _0041_;
	wire _0042_;
	wire _0043_;
	wire _0044_;
	wire _0045_;
	wire _0046_;
	wire _0047_;
	wire _0048_;
	wire _0049_;
	wire _0050_;
	wire _0051_;
	wire _0052_;
	wire _0053_;
	wire _0054_;
	wire _0055_;
	wire _0056_;
	wire _0057_;
	wire _0058_;
	wire _0059_;
	wire _0060_;
	wire _0061_;
	wire _0062_;
	wire _0063_;
	wire _0064_;
	wire _0065_;
	wire _0066_;
	wire _0067_;
	wire _0068_;
	wire _0069_;
	wire _0070_;
	wire _0071_;
	wire _0072_;
	wire _0073_;
	wire _0074_;
	wire _0075_;
	wire _0076_;
	wire _0077_;
	wire _0078_;
	wire _0079_;
	wire _0080_;
	wire _0081_;
	wire _0082_;
	wire _0083_;
	wire _0084_;
	wire _0085_;
	wire _0086_;
	wire _0087_;
	wire _0088_;
	wire _0089_;
	wire _0090_;
	wire _0091_;
	wire _0092_;
	wire _0093_;
	wire _0094_;
	wire _0095_;
	wire _0096_;
	wire _0097_;
	wire _0098_;
	wire _0099_;
	wire _0100_;
	wire _0101_;
	wire _0102_;
	wire _0103_;
	wire _0104_;
	wire _0105_;
	wire _0106_;
	wire _0107_;
	wire _0108_;
	wire _0109_;
	wire _0110_;
	wire _0111_;
	wire _0112_;
	wire _0113_;
	wire _0114_;
	wire _0115_;
	wire _0116_;
	wire _0117_;
	wire _0118_;
	wire _0119_;
	wire _0120_;
	wire _0121_;
	wire _0122_;
	wire _0123_;
	wire _0124_;
	wire _0125_;
	wire _0126_;
	wire _0127_;
	wire _0128_;
	wire _0129_;
	wire _0130_;
	wire _0131_;
	wire _0132_;
	wire _0133_;
	wire _0134_;
	wire _0135_;
	wire _0136_;
	wire _0137_;
	wire _0138_;
	wire _0139_;
	wire _0140_;
	wire _0141_;
	wire _0142_;
	wire _0143_;
	wire _0144_;
	wire _0145_;
	wire _0146_;
	wire _0147_;
	wire _0148_;
	wire _0149_;
	wire _0150_;
	wire _0151_;
	wire _0152_;
	wire _0153_;
	wire _0154_;
	wire _0155_;
	wire _0156_;
	wire _0157_;
	wire _0158_;
	wire _0159_;
	wire _0160_;
	wire _0161_;
	wire _0162_;
	wire _0163_;
	wire _0164_;
	wire _0165_;
	wire _0166_;
	wire _0167_;
	wire _0168_;
	wire _0169_;
	wire _0170_;
	wire _0171_;
	wire _0172_;
	wire _0173_;
	wire _0174_;
	wire _0175_;
	wire _0176_;
	wire _0177_;
	wire _0178_;
	wire _0179_;
	wire _0180_;
	wire _0181_;
	wire _0182_;
	wire _0183_;
	wire _0184_;
	wire _0185_;
	wire _0186_;
	wire _0187_;
	wire _0188_;
	wire _0189_;
	wire _0190_;
	wire _0191_;
	wire _0192_;
	wire _0193_;
	wire _0194_;
	wire _0195_;
	wire _0196_;
	wire _0197_;
	wire _0198_;
	wire _0199_;
	wire _0200_;
	wire _0201_;
	wire _0202_;
	wire _0203_;
	wire _0204_;
	wire _0205_;
	wire _0206_;
	wire _0207_;
	wire _0208_;
	wire _0209_;
	wire _0210_;
	wire _0211_;
	wire _0212_;
	wire _0213_;
	wire _0214_;
	wire _0215_;
	wire _0216_;
	wire _0217_;
	wire _0218_;
	wire _0219_;
	wire _0220_;
	wire _0221_;
	wire _0222_;
	wire _0223_;
	wire _0224_;
	wire _0225_;
	wire _0226_;
	wire _0227_;
	wire _0228_;
	wire _0229_;
	wire _0230_;
	wire _0231_;
	wire _0232_;
	wire _0233_;
	wire _0234_;
	wire _0235_;
	wire _0236_;
	wire _0237_;
	wire _0238_;
	wire _0239_;
	wire _0240_;
	wire _0241_;
	wire _0242_;
	wire _0243_;
	wire _0244_;
	wire _0245_;
	wire _0246_;
	wire _0247_;
	wire _0248_;
	wire _0249_;
	wire _0250_;
	wire _0251_;
	wire _0252_;
	wire _0253_;
	wire _0254_;
	wire _0255_;
	wire _0256_;
	wire _0257_;
	wire _0258_;
	wire _0259_;
	wire _0260_;
	wire _0261_;
	wire _0262_;
	wire _0263_;
	wire _0264_;
	wire _0265_;
	wire _0266_;
	wire _0267_;
	wire _0268_;
	wire _0269_;
	wire _0270_;
	wire _0271_;
	wire _0272_;
	wire _0273_;
	wire _0274_;
	wire _0275_;
	wire _0276_;
	wire _0277_;
	wire _0278_;
	wire _0279_;
	wire _0280_;
	wire _0281_;
	wire _0282_;
	wire _0283_;
	wire _0284_;
	wire _0285_;
	wire _0286_;
	wire _0287_;
	wire _0288_;
	wire _0289_;
	wire _0290_;
	wire _0291_;
	wire _0292_;
	wire _0293_;
	wire _0294_;
	wire _0295_;
	wire _0296_;
	wire _0297_;
	wire _0298_;
	wire _0299_;
	wire _0300_;
	wire _0301_;
	wire _0302_;
	wire _0303_;
	wire _0304_;
	wire _0305_;
	wire _0306_;
	wire _0307_;
	wire _0308_;
	wire _0309_;
	wire _0310_;
	wire _0311_;
	wire _0312_;
	wire _0313_;
	wire _0314_;
	wire _0315_;
	wire _0316_;
	wire _0317_;
	wire _0318_;
	wire _0319_;
	wire _0320_;
	wire _0321_;
	wire _0322_;
	wire _0323_;
	wire _0324_;
	wire _0325_;
	wire _0326_;
	wire _0327_;
	wire _0328_;
	wire _0329_;
	wire _0330_;
	wire _0331_;
	wire _0332_;
	wire _0333_;
	wire _0334_;
	wire _0335_;
	wire _0336_;
	wire _0337_;
	wire _0338_;
	wire _0339_;
	wire _0340_;
	wire _0341_;
	wire _0342_;
	wire _0343_;
	wire _0344_;
	wire _0345_;
	wire _0346_;
	wire _0347_;
	wire _0348_;
	wire _0349_;
	wire _0350_;
	wire _0351_;
	wire _0352_;
	wire _0353_;
	wire _0354_;
	wire _0355_;
	wire _0356_;
	wire _0357_;
	wire _0358_;
	wire _0359_;
	wire _0360_;
	wire _0361_;
	wire _0362_;
	wire _0363_;
	wire _0364_;
	wire _0365_;
	wire _0366_;
	wire _0367_;
	wire _0368_;
	wire _0369_;
	wire _0370_;
	wire _0371_;
	wire _0372_;
	wire _0373_;
	wire _0374_;
	wire _0375_;
	wire _0376_;
	wire _0377_;
	wire _0378_;
	wire _0379_;
	wire _0380_;
	wire _0381_;
	wire _0382_;
	wire _0383_;
	wire _0384_;
	wire _0385_;
	wire _0386_;
	wire _0387_;
	wire _0388_;
	wire _0389_;
	wire _0390_;
	wire _0391_;
	wire _0392_;
	wire _0393_;
	wire _0394_;
	wire _0395_;
	wire _0396_;
	wire _0397_;
	wire _0398_;
	wire _0399_;
	wire _0400_;
	wire _0401_;
	wire _0402_;
	wire _0403_;
	wire _0404_;
	wire _0405_;
	wire _0406_;
	wire _0407_;
	wire _0408_;
	wire _0409_;
	wire _0410_;
	wire _0411_;
	wire _0412_;
	wire _0413_;
	wire _0414_;
	wire _0415_;
	wire _0416_;
	wire _0417_;
	wire _0418_;
	wire _0419_;
	wire _0420_;
	wire _0421_;
	wire _0422_;
	wire _0423_;
	wire _0424_;
	wire _0425_;
	wire _0426_;
	wire _0427_;
	wire _0428_;
	wire _0429_;
	wire _0430_;
	wire _0431_;
	wire _0432_;
	wire _0433_;
	wire _0434_;
	wire _0435_;
	wire _0436_;
	wire _0437_;
	wire _0438_;
	wire _0439_;
	wire _0440_;
	wire _0441_;
	wire _0442_;
	wire _0443_;
	wire _0444_;
	wire _0445_;
	wire _0446_;
	wire _0447_;
	wire _0448_;
	wire _0449_;
	wire _0450_;
	wire _0451_;
	wire _0452_;
	wire _0453_;
	wire _0454_;
	wire _0455_;
	wire _0456_;
	wire _0457_;
	wire _0458_;
	wire _0459_;
	wire _0460_;
	wire _0461_;
	wire _0462_;
	wire _0463_;
	wire _0464_;
	wire _0465_;
	wire _0466_;
	wire _0467_;
	wire _0468_;
	wire _0469_;
	wire _0470_;
	wire _0471_;
	wire _0472_;
	wire _0473_;
	wire _0474_;
	wire _0475_;
	wire _0476_;
	wire _0477_;
	wire _0478_;
	wire _0479_;
	wire _0480_;
	wire _0481_;
	wire _0482_;
	wire _0483_;
	wire _0484_;
	wire _0485_;
	wire _0486_;
	wire _0487_;
	wire _0488_;
	wire _0489_;
	wire _0490_;
	wire _0491_;
	wire _0492_;
	wire _0493_;
	wire _0494_;
	wire _0495_;
	wire _0496_;
	wire _0497_;
	wire _0498_;
	wire _0499_;
	wire _0500_;
	wire _0501_;
	wire _0502_;
	wire _0503_;
	wire _0504_;
	wire _0505_;
	wire _0506_;
	wire _0507_;
	wire _0508_;
	wire _0509_;
	wire _0510_;
	wire _0511_;
	wire _0512_;
	wire _0513_;
	wire _0514_;
	wire _0515_;
	wire _0516_;
	wire _0517_;
	wire _0518_;
	wire _0519_;
	wire _0520_;
	wire _0521_;
	wire _0522_;
	wire _0523_;
	wire _0524_;
	wire _0525_;
	wire _0526_;
	wire _0527_;
	wire _0528_;
	wire _0529_;
	wire _0530_;
	wire _0531_;
	wire _0532_;
	wire _0533_;
	wire _0534_;
	wire _0535_;
	wire _0536_;
	wire _0537_;
	wire _0538_;
	wire _0539_;
	wire _0540_;
	wire _0541_;
	wire _0542_;
	wire _0543_;
	wire _0544_;
	wire _0545_;
	wire _0546_;
	wire _0547_;
	wire _0548_;
	wire _0549_;
	wire _0550_;
	wire _0551_;
	wire _0552_;
	wire _0553_;
	wire _0554_;
	wire _0555_;
	wire _0556_;
	wire _0557_;
	wire _0558_;
	wire _0559_;
	wire _0560_;
	wire _0561_;
	wire _0562_;
	wire _0563_;
	wire _0564_;
	wire _0565_;
	wire _0566_;
	wire _0567_;
	wire _0568_;
	wire _0569_;
	wire _0570_;
	wire _0571_;
	wire _0572_;
	wire _0573_;
	wire _0574_;
	wire _0575_;
	wire _0576_;
	wire _0577_;
	wire _0578_;
	wire _0579_;
	wire _0580_;
	wire _0581_;
	wire _0582_;
	wire _0583_;
	wire _0584_;
	wire _0585_;
	wire _0586_;
	wire _0587_;
	wire _0588_;
	wire _0589_;
	wire _0590_;
	wire _0591_;
	wire _0592_;
	wire _0593_;
	wire _0594_;
	wire _0595_;
	wire _0596_;
	wire _0597_;
	wire _0598_;
	wire _0599_;
	wire _0600_;
	wire _0601_;
	wire _0602_;
	wire _0603_;
	wire _0604_;
	wire _0605_;
	wire _0606_;
	wire _0607_;
	wire _0608_;
	wire _0609_;
	wire _0610_;
	wire _0611_;
	wire _0612_;
	wire _0613_;
	wire _0614_;
	wire _0615_;
	wire _0616_;
	wire _0617_;
	wire _0618_;
	wire _0619_;
	wire _0620_;
	wire _0621_;
	wire _0622_;
	wire _0623_;
	wire _0624_;
	wire _0625_;
	wire _0626_;
	wire _0627_;
	wire _0628_;
	wire _0629_;
	wire _0630_;
	wire _0631_;
	wire _0632_;
	wire _0633_;
	wire _0634_;
	wire _0635_;
	wire _0636_;
	wire _0637_;
	wire _0638_;
	wire _0639_;
	wire _0640_;
	wire _0641_;
	wire _0642_;
	wire _0643_;
	wire _0644_;
	wire _0645_;
	wire _0646_;
	wire _0647_;
	wire _0648_;
	wire _0649_;
	wire _0650_;
	wire _0651_;
	wire _0652_;
	wire _0653_;
	wire _0654_;
	wire _0655_;
	wire _0656_;
	wire _0657_;
	wire _0658_;
	wire _0659_;
	wire _0660_;
	wire _0661_;
	wire _0662_;
	wire _0663_;
	wire _0664_;
	wire _0665_;
	wire _0666_;
	wire _0667_;
	wire _0668_;
	wire _0669_;
	wire _0670_;
	wire _0671_;
	wire _0672_;
	wire _0673_;
	wire _0674_;
	wire _0675_;
	wire _0676_;
	wire _0677_;
	wire _0678_;
	wire _0679_;
	wire _0680_;
	wire _0681_;
	wire _0682_;
	wire _0683_;
	wire _0684_;
	wire _0685_;
	wire _0686_;
	wire _0687_;
	wire _0688_;
	wire _0689_;
	wire _0690_;
	wire _0691_;
	wire _0692_;
	wire _0693_;
	wire _0694_;
	wire _0695_;
	wire _0696_;
	wire _0697_;
	wire _0698_;
	wire _0699_;
	wire _0700_;
	wire _0701_;
	wire _0702_;
	wire _0703_;
	wire _0704_;
	wire _0705_;
	wire _0706_;
	wire _0707_;
	wire _0708_;
	wire _0709_;
	wire _0710_;
	wire _0711_;
	wire _0712_;
	wire _0713_;
	wire _0714_;
	wire _0715_;
	wire _0716_;
	wire _0717_;
	wire _0718_;
	wire _0719_;
	wire _0720_;
	wire _0721_;
	wire _0722_;
	wire _0723_;
	wire _0724_;
	wire _0725_;
	wire _0726_;
	wire _0727_;
	wire _0728_;
	wire _0729_;
	wire _0730_;
	wire _0731_;
	wire _0732_;
	wire _0733_;
	wire _0734_;
	wire _0735_;
	wire _0736_;
	wire _0737_;
	wire _0738_;
	wire _0739_;
	wire _0740_;
	wire _0741_;
	wire _0742_;
	wire _0743_;
	wire _0744_;
	wire _0745_;
	wire _0746_;
	wire _0747_;
	wire _0748_;
	wire _0749_;
	wire _0750_;
	wire _0751_;
	wire _0752_;
	wire _0753_;
	wire _0754_;
	wire _0755_;
	wire _0756_;
	wire _0757_;
	wire _0758_;
	wire _0759_;
	wire _0760_;
	wire _0761_;
	wire _0762_;
	wire _0763_;
	wire _0764_;
	wire _0765_;
	wire _0766_;
	wire _0767_;
	wire _0768_;
	wire _0769_;
	wire _0770_;
	wire _0771_;
	wire _0772_;
	wire _0773_;
	wire _0774_;
	wire _0775_;
	wire _0776_;
	wire _0777_;
	wire _0778_;
	wire _0779_;
	wire _0780_;
	wire _0781_;
	wire _0782_;
	wire _0783_;
	wire _0784_;
	wire _0785_;
	wire _0786_;
	wire _0787_;
	wire _0788_;
	wire _0789_;
	wire _0790_;
	wire _0791_;
	wire _0792_;
	wire _0793_;
	wire _0794_;
	wire _0795_;
	wire _0796_;
	wire _0797_;
	wire _0798_;
	wire _0799_;
	wire _0800_;
	wire _0801_;
	wire _0802_;
	wire _0803_;
	wire _0804_;
	wire _0805_;
	wire _0806_;
	wire _0807_;
	wire _0808_;
	wire _0809_;
	wire _0810_;
	wire _0811_;
	wire _0812_;
	wire _0813_;
	wire _0814_;
	wire _0815_;
	wire _0816_;
	wire _0817_;
	wire _0818_;
	wire _0819_;
	wire _0820_;
	wire _0821_;
	wire _0822_;
	wire _0823_;
	wire _0824_;
	wire _0825_;
	wire _0826_;
	wire _0827_;
	wire _0828_;
	wire _0829_;
	wire _0830_;
	wire _0831_;
	wire _0832_;
	wire _0833_;
	wire _0834_;
	wire _0835_;
	wire _0836_;
	wire _0837_;
	wire _0838_;
	wire _0839_;
	wire _0840_;
	wire _0841_;
	wire _0842_;
	wire _0843_;
	wire _0844_;
	wire _0845_;
	wire _0846_;
	wire _0847_;
	wire _0848_;
	wire _0849_;
	wire _0850_;
	wire _0851_;
	wire _0852_;
	wire _0853_;
	wire _0854_;
	wire _0855_;
	wire _0856_;
	wire _0857_;
	wire _0858_;
	wire _0859_;
	wire _0860_;
	wire _0861_;
	wire _0862_;
	wire _0863_;
	wire _0864_;
	wire _0865_;
	wire _0866_;
	wire _0867_;
	wire _0868_;
	wire _0869_;
	wire _0870_;
	wire _0871_;
	wire _0872_;
	wire _0873_;
	wire _0874_;
	wire _0875_;
	wire _0876_;
	wire _0877_;
	wire _0878_;
	wire _0879_;
	wire _0880_;
	wire _0881_;
	wire _0882_;
	wire _0883_;
	wire _0884_;
	wire _0885_;
	wire _0886_;
	wire _0887_;
	wire _0888_;
	wire _0889_;
	wire _0890_;
	wire _0891_;
	wire _0892_;
	wire _0893_;
	wire _0894_;
	wire _0895_;
	wire _0896_;
	wire _0897_;
	wire _0898_;
	wire _0899_;
	wire _0900_;
	wire _0901_;
	wire _0902_;
	wire _0903_;
	wire _0904_;
	wire _0905_;
	wire _0906_;
	wire _0907_;
	wire _0908_;
	wire _0909_;
	wire _0910_;
	wire _0911_;
	wire _0912_;
	wire _0913_;
	wire _0914_;
	wire _0915_;
	wire _0916_;
	wire _0917_;
	wire _0918_;
	wire _0919_;
	wire _0920_;
	wire _0921_;
	wire _0922_;
	wire _0923_;
	wire _0924_;
	wire _0925_;
	wire _0926_;
	wire _0927_;
	wire _0928_;
	wire _0929_;
	wire _0930_;
	wire _0931_;
	wire _0932_;
	wire _0933_;
	wire _0934_;
	wire _0935_;
	wire _0936_;
	wire _0937_;
	wire _0938_;
	wire _0939_;
	wire _0940_;
	wire _0941_;
	wire _0942_;
	wire _0943_;
	wire _0944_;
	wire _0945_;
	wire _0946_;
	wire _0947_;
	wire _0948_;
	wire _0949_;
	wire _0950_;
	wire _0951_;
	wire _0952_;
	wire _0953_;
	wire _0954_;
	wire _0955_;
	wire _0956_;
	wire _0957_;
	wire _0958_;
	wire _0959_;
	wire _0960_;
	wire _0961_;
	wire _0962_;
	wire _0963_;
	wire _0964_;
	wire _0965_;
	wire _0966_;
	wire _0967_;
	wire _0968_;
	wire _0969_;
	wire _0970_;
	wire _0971_;
	wire _0972_;
	wire _0973_;
	wire _0974_;
	wire _0975_;
	wire _0976_;
	wire _0977_;
	wire _0978_;
	wire _0979_;
	wire _0980_;
	wire _0981_;
	wire _0982_;
	wire _0983_;
	wire _0984_;
	wire _0985_;
	wire _0986_;
	wire _0987_;
	wire _0988_;
	wire _0989_;
	wire _0990_;
	wire _0991_;
	wire _0992_;
	wire _0993_;
	wire _0994_;
	wire _0995_;
	wire _0996_;
	wire _0997_;
	wire _0998_;
	wire _0999_;
	wire _1000_;
	wire _1001_;
	wire _1002_;
	wire _1003_;
	wire _1004_;
	wire _1005_;
	wire _1006_;
	wire _1007_;
	wire _1008_;
	wire _1009_;
	wire _1010_;
	wire _1011_;
	wire _1012_;
	wire _1013_;
	wire _1014_;
	wire _1015_;
	wire _1016_;
	wire _1017_;
	wire _1018_;
	wire _1019_;
	wire _1020_;
	wire _1021_;
	wire _1022_;
	wire _1023_;
	wire _1024_;
	wire _1025_;
	wire _1026_;
	wire _1027_;
	wire _1028_;
	wire _1029_;
	wire _1030_;
	wire _1031_;
	wire _1032_;
	wire _1033_;
	wire _1034_;
	wire _1035_;
	wire _1036_;
	wire _1037_;
	wire _1038_;
	wire _1039_;
	wire _1040_;
	wire _1041_;
	wire _1042_;
	wire _1043_;
	wire _1044_;
	wire _1045_;
	wire _1046_;
	wire _1047_;
	wire _1048_;
	wire _1049_;
	wire _1050_;
	wire _1051_;
	wire _1052_;
	wire _1053_;
	wire _1054_;
	wire _1055_;
	wire _1056_;
	wire _1057_;
	wire _1058_;
	wire _1059_;
	wire _1060_;
	wire _1061_;
	wire _1062_;
	wire _1063_;
	wire _1064_;
	wire _1065_;
	wire _1066_;
	wire _1067_;
	wire _1068_;
	wire _1069_;
	wire _1070_;
	wire _1071_;
	wire _1072_;
	wire _1073_;
	wire _1074_;
	wire _1075_;
	wire _1076_;
	wire _1077_;
	wire _1078_;
	wire _1079_;
	wire _1080_;
	wire _1081_;
	wire _1082_;
	wire _1083_;
	wire _1084_;
	wire _1085_;
	wire _1086_;
	wire _1087_;
	wire _1088_;
	wire _1089_;
	wire _1090_;
	wire _1091_;
	wire _1092_;
	wire _1093_;
	wire _1094_;
	wire _1095_;
	wire _1096_;
	wire _1097_;
	wire _1098_;
	wire _1099_;
	wire _1100_;
	wire _1101_;
	wire _1102_;
	wire _1103_;
	wire _1104_;
	wire _1105_;
	wire _1106_;
	wire _1107_;
	wire _1108_;
	wire _1109_;
	wire _1110_;
	wire _1111_;
	wire _1112_;
	wire _1113_;
	wire _1114_;
	wire _1115_;
	wire _1116_;
	wire _1117_;
	wire _1118_;
	wire _1119_;
	wire _1120_;
	wire _1121_;
	wire _1122_;
	wire _1123_;
	wire _1124_;
	wire _1125_;
	wire _1126_;
	wire _1127_;
	wire _1128_;
	wire _1129_;
	wire _1130_;
	wire _1131_;
	wire _1132_;
	wire _1133_;
	wire _1134_;
	wire _1135_;
	wire _1136_;
	wire _1137_;
	wire _1138_;
	wire _1139_;
	wire _1140_;
	wire _1141_;
	wire _1142_;
	wire _1143_;
	wire _1144_;
	wire _1145_;
	wire _1146_;
	wire _1147_;
	wire _1148_;
	wire _1149_;
	wire _1150_;
	wire _1151_;
	wire _1152_;
	wire _1153_;
	wire _1154_;
	wire _1155_;
	wire _1156_;
	wire _1157_;
	wire _1158_;
	wire _1159_;
	wire _1160_;
	wire _1161_;
	wire _1162_;
	wire _1163_;
	wire _1164_;
	wire _1165_;
	wire _1166_;
	wire _1167_;
	wire _1168_;
	wire _1169_;
	wire _1170_;
	wire _1171_;
	wire _1172_;
	wire _1173_;
	wire _1174_;
	wire _1175_;
	wire _1176_;
	wire _1177_;
	wire _1178_;
	wire _1179_;
	wire _1180_;
	wire _1181_;
	wire _1182_;
	wire _1183_;
	wire _1184_;
	wire _1185_;
	wire _1186_;
	wire _1187_;
	wire _1188_;
	wire _1189_;
	wire _1190_;
	wire _1191_;
	wire _1192_;
	wire _1193_;
	wire _1194_;
	wire _1195_;
	wire _1196_;
	wire _1197_;
	wire _1198_;
	wire _1199_;
	wire _1200_;
	wire _1201_;
	wire _1202_;
	wire _1203_;
	wire _1204_;
	wire _1205_;
	wire _1206_;
	wire _1207_;
	wire _1208_;
	wire _1209_;
	wire _1210_;
	wire _1211_;
	wire _1212_;
	wire _1213_;
	wire _1214_;
	wire _1215_;
	wire _1216_;
	wire _1217_;
	wire _1218_;
	wire _1219_;
	wire _1220_;
	wire _1221_;
	wire _1222_;
	wire _1223_;
	wire _1224_;
	wire _1225_;
	wire _1226_;
	wire _1227_;
	wire _1228_;
	wire _1229_;
	wire _1230_;
	wire _1231_;
	wire _1232_;
	wire _1233_;
	wire _1234_;
	wire _1235_;
	wire _1236_;
	wire _1237_;
	wire _1238_;
	wire _1239_;
	wire _1240_;
	wire _1241_;
	wire _1242_;
	wire _1243_;
	wire _1244_;
	wire _1245_;
	wire _1246_;
	wire _1247_;
	wire _1248_;
	wire _1249_;
	wire _1250_;
	wire _1251_;
	wire _1252_;
	wire _1253_;
	wire _1254_;
	wire _1255_;
	wire _1256_;
	wire _1257_;
	wire _1258_;
	wire _1259_;
	wire _1260_;
	wire _1261_;
	wire _1262_;
	wire _1263_;
	wire _1264_;
	wire _1265_;
	wire _1266_;
	wire _1267_;
	wire _1268_;
	wire _1269_;
	wire _1270_;
	wire _1271_;
	wire _1272_;
	wire _1273_;
	wire _1274_;
	wire _1275_;
	wire _1276_;
	wire _1277_;
	wire _1278_;
	wire _1279_;
	wire _1280_;
	wire _1281_;
	wire _1282_;
	wire _1283_;
	wire _1284_;
	wire _1285_;
	wire _1286_;
	wire _1287_;
	wire _1288_;
	wire _1289_;
	wire _1290_;
	wire _1291_;
	wire _1292_;
	wire _1293_;
	wire _1294_;
	wire _1295_;
	wire _1296_;
	wire _1297_;
	wire _1298_;
	wire _1299_;
	wire _1300_;
	wire _1301_;
	wire _1302_;
	wire _1303_;
	wire _1304_;
	wire _1305_;
	wire _1306_;
	wire _1307_;
	wire _1308_;
	wire _1309_;
	wire _1310_;
	wire _1311_;
	wire _1312_;
	wire _1313_;
	wire _1314_;
	wire _1315_;
	wire _1316_;
	wire _1317_;
	wire _1318_;
	wire _1319_;
	wire _1320_;
	wire _1321_;
	wire _1322_;
	wire _1323_;
	wire _1324_;
	wire _1325_;
	wire _1326_;
	wire _1327_;
	wire _1328_;
	wire _1329_;
	wire _1330_;
	wire _1331_;
	wire _1332_;
	wire _1333_;
	wire _1334_;
	wire _1335_;
	wire _1336_;
	wire _1337_;
	wire _1338_;
	wire _1339_;
	wire _1340_;
	wire _1341_;
	wire _1342_;
	wire _1343_;
	wire _1344_;
	wire _1345_;
	wire _1346_;
	wire _1347_;
	wire _1348_;
	wire _1349_;
	wire _1350_;
	wire _1351_;
	wire _1352_;
	wire _1353_;
	wire _1354_;
	wire _1355_;
	wire _1356_;
	wire _1357_;
	wire _1358_;
	wire _1359_;
	wire _1360_;
	wire _1361_;
	wire _1362_;
	wire _1363_;
	wire _1364_;
	wire _1365_;
	wire _1366_;
	wire _1367_;
	wire _1368_;
	wire _1369_;
	wire _1370_;
	wire _1371_;
	wire _1372_;
	wire _1373_;
	wire _1374_;
	wire _1375_;
	wire _1376_;
	wire _1377_;
	wire _1378_;
	wire _1379_;
	wire _1380_;
	wire _1381_;
	wire _1382_;
	wire _1383_;
	wire _1384_;
	wire _1385_;
	wire _1386_;
	wire _1387_;
	wire _1388_;
	wire _1389_;
	wire _1390_;
	wire _1391_;
	wire _1392_;
	wire _1393_;
	wire _1394_;
	wire _1395_;
	wire _1396_;
	wire _1397_;
	wire _1398_;
	wire _1399_;
	wire _1400_;
	wire _1401_;
	wire _1402_;
	wire _1403_;
	wire _1404_;
	wire _1405_;
	wire _1406_;
	wire _1407_;
	wire _1408_;
	wire _1409_;
	wire _1410_;
	wire _1411_;
	wire _1412_;
	wire _1413_;
	wire _1414_;
	wire _1415_;
	wire _1416_;
	wire _1417_;
	wire _1418_;
	wire _1419_;
	wire _1420_;
	wire _1421_;
	wire _1422_;
	wire _1423_;
	wire _1424_;
	wire _1425_;
	wire _1426_;
	wire _1427_;
	wire _1428_;
	wire _1429_;
	wire _1430_;
	wire _1431_;
	wire _1432_;
	wire _1433_;
	wire _1434_;
	wire _1435_;
	wire _1436_;
	wire _1437_;
	wire _1438_;
	wire _1439_;
	wire _1440_;
	wire _1441_;
	wire _1442_;
	wire _1443_;
	wire _1444_;
	wire _1445_;
	wire _1446_;
	wire _1447_;
	wire _1448_;
	wire _1449_;
	wire _1450_;
	wire _1451_;
	wire _1452_;
	wire _1453_;
	wire _1454_;
	wire _1455_;
	wire _1456_;
	wire _1457_;
	wire _1458_;
	wire _1459_;
	wire _1460_;
	wire _1461_;
	wire _1462_;
	wire _1463_;
	wire _1464_;
	wire _1465_;
	wire _1466_;
	wire _1467_;
	wire _1468_;
	wire _1469_;
	wire _1470_;
	wire _1471_;
	wire _1472_;
	wire _1473_;
	wire _1474_;
	wire _1475_;
	wire _1476_;
	wire _1477_;
	wire _1478_;
	wire _1479_;
	wire _1480_;
	wire _1481_;
	wire _1482_;
	wire _1483_;
	wire _1484_;
	wire _1485_;
	wire _1486_;
	wire _1487_;
	wire _1488_;
	wire _1489_;
	wire _1490_;
	wire _1491_;
	wire _1492_;
	wire _1493_;
	wire _1494_;
	wire _1495_;
	wire _1496_;
	wire _1497_;
	wire [2:0] _1498_;
	wire [2:0] _1499_;
	input wire [13:0] io_in;
	output wire [13:0] io_out;
	wire \mchip.clock ;
	wire [11:0] \mchip.io_in ;
	wire [11:0] \mchip.io_out ;
	wire [7:0] \mchip.my_core.ACC ;
	wire \mchip.my_core.A_en ;
	wire [7:0] \mchip.my_core.A_in ;
	wire [7:0] \mchip.my_core.A_out ;
	wire \mchip.my_core.A_rst ;
	wire [7:0] \mchip.my_core.B_out ;
	wire \mchip.my_core.B_rst ;
	wire [2:0] \mchip.my_core.Brain.D5_3 ;
	wire [2:0] \mchip.my_core.Brain.DDD ;
	wire \mchip.my_core.Brain.Intr ;
	wire \mchip.my_core.Brain.Ready ;
	wire [2:0] \mchip.my_core.Brain.SSS ;
	wire \mchip.my_core.Brain.clk ;
	wire [39:0] \mchip.my_core.Brain.ctrl_signals ;
	reg [2:0] \mchip.my_core.Brain.cycle ;
	wire [3:0] \mchip.my_core.Brain.flags ;
	wire [7:0] \mchip.my_core.Brain.instr ;
	wire [2:0] \mchip.my_core.Brain.next_state ;
	wire \mchip.my_core.Brain.rst ;
	reg [2:0] \mchip.my_core.Brain.state ;
	wire [7:0] \mchip.my_core.D_in ;
	wire [7:0] \mchip.my_core.D_out ;
	wire \mchip.my_core.INTR ;
	reg [7:0] \mchip.my_core.IR.Q ;
	wire \mchip.my_core.IR.clear ;
	wire \mchip.my_core.IR.clk ;
	wire [7:0] \mchip.my_core.IR.d ;
	wire \mchip.my_core.IR.en ;
	wire \mchip.my_core.IR_en ;
	wire \mchip.my_core.IR_rst ;
	reg \mchip.my_core.Intr ;
	wire \mchip.my_core.READY ;
	reg \mchip.my_core.Ready ;
	reg [2:0] \mchip.my_core.SP_SEL.Q ;
	wire \mchip.my_core.SP_SEL.clear ;
	wire \mchip.my_core.SP_SEL.clk ;
	wire [2:0] \mchip.my_core.SP_SEL.d ;
	wire \mchip.my_core.SP_SEL.load ;
	wire \mchip.my_core.SP_SEL.up ;
	wire \mchip.my_core.SP_rst ;
	reg \mchip.my_core.S_Intr ;
	wire [7:0] \mchip.my_core.Stack.RST_AAA ;
	wire [6:0] \mchip.my_core.Stack.Stack_ctrl ;
	wire [7:0] \mchip.my_core.Stack.bus ;
	wire \mchip.my_core.Stack.clk ;
	reg [13:0] \mchip.my_core.Stack.rf[0] ;
	reg [13:0] \mchip.my_core.Stack.rf[1] ;
	reg [13:0] \mchip.my_core.Stack.rf[2] ;
	reg [13:0] \mchip.my_core.Stack.rf[3] ;
	reg [13:0] \mchip.my_core.Stack.rf[4] ;
	reg [13:0] \mchip.my_core.Stack.rf[5] ;
	reg [13:0] \mchip.my_core.Stack.rf[6] ;
	reg [13:0] \mchip.my_core.Stack.rf[7] ;
	wire \mchip.my_core.Stack.rst ;
	wire [2:0] \mchip.my_core.Stack.sel ;
	wire [7:0] \mchip.my_core.Stack.upper ;
	wire \mchip.my_core.Sync ;
	wire [9:0] \mchip.my_core.Unit.ALU_ctrl ;
	wire \mchip.my_core.Unit.Flag_rst ;
	wire [7:0] \mchip.my_core.Unit.a ;
	wire [7:0] \mchip.my_core.Unit.b ;
	wire \mchip.my_core.Unit.clk ;
	wire [3:0] \mchip.my_core.Unit.flag_in ;
	reg [3:0] \mchip.my_core.Unit.flag_reg.Q ;
	wire \mchip.my_core.Unit.flag_reg.clear ;
	wire \mchip.my_core.Unit.flag_reg.clk ;
	wire [3:0] \mchip.my_core.Unit.flag_reg.d ;
	wire \mchip.my_core.Unit.flag_reg.en ;
	wire [3:0] \mchip.my_core.Unit.flags ;
	wire \mchip.my_core.Unit.rst ;
	wire [7:0] \mchip.my_core.bus ;
	wire \mchip.my_core.clk ;
	wire [39:0] \mchip.my_core.ctrl_signals ;
	wire [3:0] \mchip.my_core.flags ;
	wire [7:0] \mchip.my_core.instr ;
	reg [7:0] \mchip.my_core.regA.Q ;
	wire \mchip.my_core.regA.clear ;
	wire \mchip.my_core.regA.clk ;
	wire [7:0] \mchip.my_core.regA.d ;
	wire \mchip.my_core.regA.en ;
	reg [7:0] \mchip.my_core.regB.Q ;
	wire \mchip.my_core.regB.clear ;
	wire \mchip.my_core.regB.clk ;
	wire [7:0] \mchip.my_core.regB.d ;
	wire \mchip.my_core.regB.en ;
	wire [7:0] \mchip.my_core.rf.ACC ;
	wire [7:0] \mchip.my_core.rf.bus ;
	wire \mchip.my_core.rf.clk ;
	reg [7:0] \mchip.my_core.rf.rf[0] ;
	reg [7:0] \mchip.my_core.rf.rf[1] ;
	reg [7:0] \mchip.my_core.rf.rf[2] ;
	reg [7:0] \mchip.my_core.rf.rf[3] ;
	reg [7:0] \mchip.my_core.rf.rf[4] ;
	reg [7:0] \mchip.my_core.rf.rf[5] ;
	reg [7:0] \mchip.my_core.rf.rf[6] ;
	reg [7:0] \mchip.my_core.rf.rf[7] ;
	wire [4:0] \mchip.my_core.rf.rf_ctrl ;
	wire \mchip.my_core.rf.rst ;
	wire \mchip.my_core.rst ;
	wire [2:0] \mchip.my_core.sel_Stack ;
	wire [2:0] \mchip.my_core.state ;
	reg \mchip.my_core.tempR ;
	wire \mchip.reset ;
	assign _0983_ = \mchip.my_core.IR.Q [5] | ~\mchip.my_core.IR.Q [6];
	assign _0984_ = \mchip.my_core.IR.Q [4] | ~\mchip.my_core.IR.Q [0];
	assign _0985_ = _0984_ | _0983_;
	assign _0986_ = _0921_ & ~_0985_;
	assign _0987_ = _0986_ | _0982_;
	assign _0988_ = _0976_ | _0878_;
	assign _0989_ = _0921_ & ~_0988_;
	assign _0990_ = _0947_ & ~\mchip.my_core.IR.Q [7];
	assign _0991_ = _0990_ | _0989_;
	assign _0992_ = _0991_ | _0987_;
	assign _0993_ = _0992_ | _0980_;
	assign _0994_ = _0993_ | _0974_;
	assign _0995_ = ~(_0994_ & _0933_);
	assign _0996_ = _0995_ | _0892_;
	assign _0997_ = \mchip.my_core.Brain.cycle [0] & ~_0996_;
	assign _0998_ = _0997_ | _0972_;
	assign _0999_ = _0998_ | _0952_;
	assign _0003_ = _0999_ | _0940_;
	assign _1000_ = \mchip.my_core.IR.Q [2] | ~\mchip.my_core.IR.Q [3];
	assign _1001_ = ~(_1000_ | _0878_);
	assign _1002_ = \mchip.my_core.IR.Q [4] | \mchip.my_core.IR.Q [5];
	assign _1003_ = ~(_1002_ | _0914_);
	assign _1004_ = _1003_ & _1001_;
	assign _1005_ = \mchip.my_core.IR.Q [3] | \mchip.my_core.IR.Q [2];
	assign _1006_ = ~(_1005_ | _0878_);
	assign _1007_ = _1006_ & _1003_;
	assign _1008_ = ~(_1007_ | _1004_);
	assign _1009_ = \mchip.my_core.IR.Q [6] | \mchip.my_core.IR.Q [2];
	assign _1010_ = _1009_ | _0883_;
	assign _1011_ = _1010_ | \mchip.my_core.IR.Q [7];
	assign _1012_ = \mchip.my_core.IR.Q [1] | ~\mchip.my_core.IR.Q [0];
	assign _1013_ = _1012_ | _1009_;
	assign _1014_ = _0921_ & ~_1013_;
	assign _1015_ = _1011_ & ~_1014_;
	assign _1016_ = _1015_ & _1008_;
	assign _1017_ = \mchip.my_core.IR.Q [5] | ~\mchip.my_core.IR.Q [4];
	assign _1018_ = _1017_ | _0914_;
	assign _1019_ = _1001_ & ~_1018_;
	assign _1020_ = _1006_ & ~_1018_;
	assign _1021_ = _1020_ | _1019_;
	assign _1022_ = _1016_ & ~_1021_;
	assign _1023_ = _0890_ & ~_0899_;
	assign _1024_ = ~_1023_;
	assign _1025_ = _1024_ | _1022_;
	assign _1026_ = \mchip.my_core.Brain.cycle [0] & ~_1025_;
	assign _1027_ = ~(\mchip.my_core.Brain.cycle [0] | \mchip.my_core.Brain.cycle [2]);
	assign _1028_ = _1026_ & ~_1027_;
	assign _1029_ = _1008_ & ~_1021_;
	assign _1030_ = \mchip.my_core.IR.Q [5] & ~_1029_;
	assign _1031_ = _1015_ & ~_1030_;
	assign _1032_ = _1029_ & _1015_;
	assign _1033_ = _1032_ | _1031_;
	assign _1034_ = _1033_ | _1024_;
	assign _0680_ = \mchip.my_core.Brain.cycle [0] & ~_1034_;
	assign _1035_ = ~\mchip.my_core.IR.Q [4];
	assign _1036_ = _1029_ | _1035_;
	assign _1037_ = _1036_ | _1032_;
	assign _1038_ = _1037_ | _1024_;
	assign _1039_ = \mchip.my_core.Brain.cycle [0] & ~_1038_;
	assign _1040_ = ~\mchip.my_core.IR.Q [3];
	assign _1041_ = _1029_ | _1040_;
	assign _1042_ = _0883_ | \mchip.my_core.IR.Q [2];
	assign _1043_ = _1042_ & ~_1015_;
	assign _1044_ = _1041_ & ~_1043_;
	assign _1045_ = _1044_ | _1032_;
	assign _1046_ = _1045_ | _1024_;
	assign _1047_ = \mchip.my_core.Brain.cycle [0] & ~_1046_;
	assign _1048_ = _0680_ & ~_1039_;
	assign _1049_ = _1048_ | ~_1028_;
	assign _1050_ = ~\mchip.my_core.Brain.cycle [2];
	assign _1051_ = (\mchip.my_core.IR.Q [7] ? _0981_ : _0977_);
	assign _1052_ = _1051_ | _1024_;
	assign _1053_ = _1052_ | _1050_;
	assign _1054_ = \mchip.my_core.IR.Q [7] & ~\mchip.my_core.IR.Q [6];
	assign _1055_ = _1054_ | _1007_;
	assign _1056_ = _1015_ & ~_1055_;
	assign _1057_ = _1020_ | _1004_;
	assign _1058_ = _1057_ | _1019_;
	assign _1059_ = _1056_ & ~_1058_;
	assign _1060_ = _1059_ | _1024_;
	assign _1061_ = \mchip.my_core.Brain.cycle [0] & ~_1060_;
	assign _1062_ = _1053_ & ~_1061_;
	assign _1063_ = ~(_1062_ | _1027_);
	assign _0017_ = _1063_ & _1049_;
	assign _1064_ = ~\mchip.my_core.Brain.cycle [0];
	assign _1065_ = \mchip.my_core.Brain.cycle [2] | \mchip.my_core.Brain.cycle [1];
	assign _1066_ = _1064_ & ~_1065_;
	assign _1067_ = ~_1066_;
	assign _1068_ = _0989_ | _0958_;
	assign _1069_ = ~(_1068_ | _0986_);
	assign _1070_ = _1002_ | ~_0880_;
	assign _1071_ = \mchip.my_core.IR.Q [0] & ~_1070_;
	assign _1072_ = _1071_ | _1040_;
	assign _1073_ = _1072_ | _1069_;
	assign _1074_ = _1073_ | _1024_;
	assign _1075_ = _0982_ | _0958_;
	assign _1076_ = ~(_1075_ | _0564_);
	assign _1077_ = ~(_0896_ & \mchip.my_core.Brain.state [2]);
	assign _1078_ = ~(_1077_ | _1076_);
	assign _1079_ = _1074_ & ~_1078_;
	assign _1080_ = _1079_ | _0897_;
	assign _1081_ = _1080_ | _1050_;
	assign _1082_ = _1077_ | _0919_;
	assign _1083_ = \mchip.my_core.Brain.cycle [1] & ~_1082_;
	assign _1084_ = _1081_ & ~_1083_;
	assign _1085_ = ~(_1023_ | _0900_);
	assign _1086_ = ~_0960_;
	assign _1087_ = ~(_1011_ & _1086_);
	assign _1088_ = ~(_1087_ | _1014_);
	assign _1089_ = _1088_ | _1040_;
	assign _1090_ = _1089_ | _1024_;
	assign _1091_ = ~(_1054_ | _0960_);
	assign _1092_ = _1091_ & _1015_;
	assign _1093_ = _1015_ | _1040_;
	assign _1094_ = \mchip.my_core.IR.Q [7] & \mchip.my_core.IR.Q [0];
	assign _1095_ = _1093_ & ~_1094_;
	assign _1096_ = _1095_ | _1092_;
	assign _1097_ = _0900_ & ~_1096_;
	assign _1098_ = _1090_ & ~_1097_;
	assign _1099_ = _1098_ | _1085_;
	assign _1100_ = \mchip.my_core.Brain.cycle [0] & ~_1099_;
	assign _1101_ = _1084_ & ~_1100_;
	assign _1102_ = _1067_ & ~_1101_;
	assign _1103_ = _0897_ & ~_0919_;
	assign _1104_ = ~(_1103_ & \mchip.my_core.Brain.cycle [1]);
	assign _1105_ = _1071_ | _1035_;
	assign _1106_ = _1105_ | _1069_;
	assign _1107_ = _1106_ | _1024_;
	assign _1108_ = (_0897_ ? _1076_ : _1107_);
	assign _1109_ = \mchip.my_core.Brain.cycle [2] & ~_1108_;
	assign _1110_ = _1104_ & ~_1109_;
	assign _1111_ = _1088_ | _1035_;
	assign _1112_ = _1111_ | _1024_;
	assign _1113_ = _1015_ | _1035_;
	assign _1114_ = \mchip.my_core.IR.Q [7] & \mchip.my_core.IR.Q [1];
	assign _1115_ = _1113_ & ~_1114_;
	assign _1116_ = _1115_ | _1092_;
	assign _1117_ = _0900_ & ~_1116_;
	assign _1118_ = _1112_ & ~_1117_;
	assign _1119_ = _1118_ | _1085_;
	assign _1120_ = \mchip.my_core.Brain.cycle [0] & ~_1119_;
	assign _1121_ = _1110_ & ~_1120_;
	assign _1122_ = _1121_ | ~_1067_;
	assign _1123_ = _1122_ | ~_1102_;
	assign _1124_ = ~\mchip.my_core.Brain.cycle [1];
	assign _1125_ = _1082_ & ~_1103_;
	assign _1126_ = _1125_ | _1124_;
	assign _1127_ = ~\mchip.my_core.IR.Q [5];
	assign _1128_ = _1071_ | _1127_;
	assign _1129_ = _1128_ | _1069_;
	assign _1130_ = _1129_ | _1024_;
	assign _1131_ = _1130_ & ~_1078_;
	assign _1132_ = (_0897_ ? _1076_ : _1131_);
	assign _1133_ = \mchip.my_core.Brain.cycle [2] & ~_1132_;
	assign _1134_ = _1126_ & ~_1133_;
	assign _1135_ = _1088_ | _1127_;
	assign _1136_ = _1135_ | _1024_;
	assign _1137_ = _1015_ | _1127_;
	assign _1138_ = \mchip.my_core.IR.Q [7] & \mchip.my_core.IR.Q [2];
	assign _1139_ = _1137_ & ~_1138_;
	assign _1140_ = _1139_ | _1092_;
	assign _1141_ = _0900_ & ~_1140_;
	assign _1142_ = _1136_ & ~_1141_;
	assign _1143_ = _1142_ | _1085_;
	assign _1144_ = \mchip.my_core.Brain.cycle [0] & ~_1143_;
	assign _1145_ = _1134_ & ~_1144_;
	assign _1146_ = _1145_ | ~_1067_;
	assign _1147_ = ~(_1146_ | _1123_);
	assign _1148_ = _1054_ | _1014_;
	assign _1149_ = _1148_ | _1087_;
	assign _1150_ = _1029_ & ~_1149_;
	assign _1151_ = _1068_ | _0987_;
	assign _1152_ = ~(_1151_ | _0978_);
	assign _1153_ = (\mchip.my_core.Brain.cycle [2] ? _1152_ : _1150_);
	assign _1154_ = _1153_ | _1024_;
	assign _1155_ = _1154_ | _1027_;
	assign _1156_ = _1155_ | _1147_;
	assign _1157_ = ~(_1156_ & _0933_);
	assign _1158_ = _0933_ & ~_1156_;
	assign _1159_ = _1158_ & ~_1102_;
	assign _1160_ = _1158_ & _1146_;
	assign _1161_ = _1158_ & ~_1122_;
	assign _1162_ = ~(_1161_ & _1160_);
	assign _1163_ = _1162_ | _1159_;
	assign _0057_ = _1157_ & ~_1163_;
	assign _0005_ = _0057_ | io_in[13];
	assign _1164_ = ~_1159_;
	assign _1165_ = _1162_ | _1164_;
	assign _0056_ = _1157_ & ~_1165_;
	assign _0006_ = _0056_ | io_in[13];
	assign _1166_ = _1161_ | ~_1160_;
	assign _1167_ = _1166_ | _1159_;
	assign _0055_ = _1157_ & ~_1167_;
	assign _0007_ = _0055_ | io_in[13];
	assign _1168_ = _1166_ | _1164_;
	assign _0054_ = _1157_ & ~_1168_;
	assign _0008_ = _0054_ | io_in[13];
	assign _1169_ = _0890_ | _0889_;
	assign _1170_ = (\mchip.my_core.Brain.state [2] ? _0888_ : _0896_);
	assign _1171_ = _1170_ | _0897_;
	assign _1172_ = _1171_ | _1169_;
	assign _1173_ = ~(_0928_ | _0909_);
	assign _1174_ = _1173_ | _1172_;
	assign _1175_ = _1174_ | _1124_;
	assign _1176_ = _0909_ | _0886_;
	assign _1177_ = _0989_ | _0978_;
	assign _1178_ = _1177_ | _0927_;
	assign _1179_ = _1178_ | _1176_;
	assign _1180_ = _0919_ & ~_1179_;
	assign _1181_ = _1180_ | _1172_;
	assign _1182_ = \mchip.my_core.Brain.cycle [2] & ~_1181_;
	assign _1183_ = _1175_ & ~_1182_;
	assign _1184_ = \mchip.my_core.Brain.cycle [0] & ~_1172_;
	assign _1185_ = _1183_ & ~_1184_;
	assign _1186_ = _1185_ | ~_1067_;
	assign _1187_ = ~_0897_;
	assign _1188_ = _1187_ & ~_1023_;
	assign _1189_ = _1188_ | _1173_;
	assign _1190_ = _1189_ | _1124_;
	assign _1191_ = _1180_ | ~_0897_;
	assign _1192_ = \mchip.my_core.Brain.cycle [2] & ~_1191_;
	assign _1193_ = _1190_ & ~_1192_;
	assign _1194_ = _1012_ | _0976_;
	assign _1195_ = _1194_ | \mchip.my_core.IR.Q [7];
	assign _1196_ = _1195_ | _1024_;
	assign _1197_ = _1196_ & ~_0897_;
	assign _1198_ = \mchip.my_core.Brain.cycle [0] & ~_1197_;
	assign _1199_ = _1193_ & ~_1198_;
	assign _1200_ = _1199_ | ~_1067_;
	assign _1201_ = ~(\mchip.my_core.Brain.cycle [0] | \mchip.my_core.Brain.cycle [1]);
	assign _1202_ = (\mchip.my_core.Brain.cycle [1] ? _1173_ : _1195_);
	assign _1203_ = _1202_ | _1085_;
	assign _1204_ = _1203_ | _1124_;
	assign _1205_ = \mchip.my_core.Brain.cycle [0] & ~_1203_;
	assign _1206_ = _1204_ & ~_1205_;
	assign _1207_ = _1206_ | _1201_;
	assign _1208_ = _1200_ & ~_1207_;
	assign _1209_ = _1208_ | _1186_;
	assign _1210_ = ~(_1207_ | _1200_);
	assign _1211_ = _1210_ | _1209_;
	assign _1212_ = _0933_ & ~_1211_;
	assign _1213_ = _0933_ & ~_1207_;
	assign _1214_ = _1213_ | _1212_;
	assign _1215_ = ~(\mchip.my_core.SP_SEL.Q [2] & \mchip.my_core.SP_SEL.Q [1]);
	assign _1216_ = _1215_ | _1498_[0];
	assign _0053_ = _1214_ & ~_1216_;
	assign _0009_ = _0053_ | io_in[13];
	assign _1217_ = _1215_ | \mchip.my_core.SP_SEL.Q [0];
	assign _0052_ = _1214_ & ~_1217_;
	assign _0010_ = _0052_ | io_in[13];
	assign _1218_ = \mchip.my_core.SP_SEL.Q [1] | ~\mchip.my_core.SP_SEL.Q [2];
	assign _1219_ = _1218_ | _1498_[0];
	assign _0051_ = _1214_ & ~_1219_;
	assign _0011_ = _0051_ | io_in[13];
	assign _1220_ = _1218_ | \mchip.my_core.SP_SEL.Q [0];
	assign _0050_ = _1214_ & ~_1220_;
	assign _0012_ = _0050_ | io_in[13];
	assign _1221_ = \mchip.my_core.SP_SEL.Q [2] | ~\mchip.my_core.SP_SEL.Q [1];
	assign _1222_ = _1221_ | _1498_[0];
	assign _0049_ = _1214_ & ~_1222_;
	assign _0013_ = _0049_ | io_in[13];
	assign _1223_ = _1221_ | \mchip.my_core.SP_SEL.Q [0];
	assign _0048_ = _1214_ & ~_1223_;
	assign _0014_ = _0048_ | io_in[13];
	assign _1224_ = \mchip.my_core.SP_SEL.Q [2] | \mchip.my_core.SP_SEL.Q [1];
	assign _1225_ = _1224_ | _1498_[0];
	assign _0047_ = _1214_ & ~_1225_;
	assign _0015_ = _0047_ | io_in[13];
	assign _1226_ = _1224_ | \mchip.my_core.SP_SEL.Q [0];
	assign _0046_ = _1214_ & ~_1226_;
	assign _0016_ = _0046_ | io_in[13];
	assign _1227_ = _0897_ & ~_0899_;
	assign _0019_ = _1227_ | io_in[13];
	assign _1228_ = ~(_1085_ & _0898_);
	assign _1229_ = ~(_1176_ | _0924_);
	assign _1230_ = _0983_ | \mchip.my_core.IR.Q [7];
	assign _1231_ = _0878_ | \mchip.my_core.IR.Q [2];
	assign _1232_ = _1231_ | _1230_;
	assign _1233_ = _1232_ | ~_0876_;
	assign _1234_ = _0886_ & ~_1233_;
	assign _1235_ = _0942_ | \mchip.my_core.IR.Q [7];
	assign _1236_ = _1235_ | _1231_;
	assign _1237_ = _1236_ | _0876_;
	assign _1238_ = _0909_ & ~_1237_;
	assign _1239_ = _1238_ | _1234_;
	assign _1240_ = ~(_1239_ | _0924_);
	assign _1241_ = _1240_ | _1229_;
	assign _1242_ = _1241_ | _1228_;
	assign _1243_ = _1242_ | _1124_;
	assign _1244_ = _1012_ | ~\mchip.my_core.IR.Q [2];
	assign _1245_ = _1244_ | _0914_;
	assign _1246_ = _1245_ | _1228_;
	assign _1247_ = \mchip.my_core.Brain.cycle [0] & ~_1246_;
	assign _1248_ = _1243_ & ~_1247_;
	assign _1249_ = ~(_1248_ | _1201_);
	assign _1250_ = ~\mchip.my_core.SP_SEL.Q [2];
	assign _1251_ = \mchip.my_core.SP_SEL.Q [1] | \mchip.my_core.SP_SEL.Q [0];
	assign _1252_ = _1250_ & ~_1251_;
	assign _1253_ = _1252_ & ~_1249_;
	assign _1254_ = _0981_ | \mchip.my_core.IR.Q [7];
	assign _1255_ = _0956_ | _0877_;
	assign _1256_ = ~(_1255_ | _0914_);
	assign _1257_ = _1254_ & ~_1256_;
	assign _1258_ = _0956_ | _0904_;
	assign _1259_ = ~(_1258_ | _0914_);
	assign _1260_ = _1257_ & ~_1259_;
	assign _1261_ = _1260_ | ~_0900_;
	assign _1262_ = ~_0900_;
	assign _1263_ = _1023_ | ~_0898_;
	assign _1264_ = _1262_ & ~_1263_;
	assign _1265_ = (_1264_ ? _1245_ : _1261_);
	assign _1266_ = \mchip.my_core.Brain.cycle [0] & ~_1265_;
	assign _1267_ = _1243_ & ~_1266_;
	assign _1268_ = _1267_ | _1201_;
	assign _1269_ = _1268_ | _1253_;
	assign _1270_ = ~(\mchip.my_core.SP_SEL.Q [1] & \mchip.my_core.SP_SEL.Q [0]);
	assign _1271_ = _1270_ | _1250_;
	assign _1272_ = _1249_ & ~_1271_;
	assign _1273_ = _1269_ | _1272_;
	assign _0062_ = (_1249_ ? _1273_ : _1269_);
	assign _1274_ = _1048_ & _1028_;
	assign _0018_ = _1063_ & ~_1274_;
	assign _1275_ = ~(_0948_ & _0933_);
	assign _1276_ = _1275_ | _0892_;
	assign _1277_ = \mchip.my_core.Brain.cycle [2] & ~_1276_;
	assign _1278_ = ~(_0909_ & _0876_);
	assign _1279_ = _1278_ | _0893_;
	assign _1280_ = \mchip.my_core.Brain.cycle [1] & ~_1279_;
	assign _1281_ = _0919_ | io_in[13];
	assign _1282_ = _1281_ | _0892_;
	assign _1283_ = \mchip.my_core.Brain.cycle [1] & ~_1282_;
	assign _1284_ = _1283_ | _1280_;
	assign _1285_ = _1284_ | _1277_;
	assign _1286_ = _0564_ | _0941_;
	assign _1287_ = \mchip.my_core.Brain.cycle [0] & ~_1286_;
	assign _1288_ = _0898_ | io_in[13];
	assign _1289_ = \mchip.my_core.Brain.cycle [0] & ~_1288_;
	assign _1290_ = _1289_ | _1287_;
	assign _1291_ = _1023_ & ~io_in[13];
	assign _1292_ = _0876_ | ~_0886_;
	assign _1293_ = _1292_ | _0893_;
	assign _1294_ = \mchip.my_core.Brain.cycle [1] & ~_1293_;
	assign _1295_ = _1294_ | _1291_;
	assign _1296_ = _1295_ | _1290_;
	assign _1297_ = _0954_ | _0892_;
	assign _1298_ = _1297_ | _0970_;
	assign _1299_ = \mchip.my_core.Brain.cycle [0] & ~_1298_;
	assign _1300_ = _1259_ | _1256_;
	assign _1301_ = ~(_1300_ & _0933_);
	assign _1302_ = _1301_ | _0892_;
	assign _1303_ = \mchip.my_core.Brain.cycle [0] & ~_1302_;
	assign _1304_ = _1303_ | _1299_;
	assign _1305_ = _1300_ | _0969_;
	assign _1306_ = _0994_ | io_in[13];
	assign _1307_ = _1306_ | _1305_;
	assign _1308_ = _1307_ | _0892_;
	assign _1309_ = \mchip.my_core.Brain.cycle [0] & ~_1308_;
	assign _1310_ = _1309_ | io_in[13];
	assign _1311_ = _1310_ | _1304_;
	assign _1312_ = _1311_ | _1296_;
	assign _0001_ = _1312_ | _1285_;
	assign _1313_ = _1161_ | _1160_;
	assign _1314_ = _1313_ | _1164_;
	assign _0058_ = _1157_ & ~_1314_;
	assign _0004_ = _0058_ | io_in[13];
	assign \mchip.my_core.IR.en  = \mchip.my_core.Ready  & \mchip.my_core.Brain.cycle [0];
	assign _0020_ = _0062_ ^ _1498_[0];
	assign _1315_ = _1249_ & ~_1273_;
	assign _1316_ = ~(_1315_ ^ \mchip.my_core.SP_SEL.Q [1]);
	assign _1499_[1] = _1316_ ^ \mchip.my_core.SP_SEL.Q [0];
	assign _0021_ = (_0062_ ? \mchip.my_core.SP_SEL.Q [1] : _1499_[1]);
	assign _1317_ = \mchip.my_core.SP_SEL.Q [1] & ~_1315_;
	assign _1318_ = _1316_ & ~_1498_[0];
	assign _1319_ = _1318_ | _1317_;
	assign _1320_ = _1315_ ^ _1250_;
	assign _1499_[2] = _1320_ ^ _1319_;
	assign _0022_ = (_0062_ ? \mchip.my_core.SP_SEL.Q [2] : _1499_[2]);
	assign _1321_ = (_0000_[0] ? \mchip.my_core.Stack.rf[1] [8] : \mchip.my_core.Stack.rf[0] [8]);
	assign _1322_ = (_0000_[0] ? \mchip.my_core.Stack.rf[3] [8] : \mchip.my_core.Stack.rf[2] [8]);
	assign _1323_ = (_0000_[1] ? _1322_ : _1321_);
	assign _1324_ = (_0000_[0] ? \mchip.my_core.Stack.rf[5] [8] : \mchip.my_core.Stack.rf[4] [8]);
	assign _1325_ = (_0000_[0] ? \mchip.my_core.Stack.rf[7] [8] : \mchip.my_core.Stack.rf[6] [8]);
	assign _1326_ = (_0000_[1] ? _1325_ : _1324_);
	assign _1327_ = (_0000_[2] ? _1326_ : _1323_);
	assign _1328_ = (_0000_[0] ? \mchip.my_core.Stack.rf[1] [0] : \mchip.my_core.Stack.rf[0] [0]);
	assign _1329_ = (_0000_[0] ? \mchip.my_core.Stack.rf[3] [0] : \mchip.my_core.Stack.rf[2] [0]);
	assign _1330_ = (_0000_[1] ? _1329_ : _1328_);
	assign _1331_ = (_0000_[0] ? \mchip.my_core.Stack.rf[5] [0] : \mchip.my_core.Stack.rf[4] [0]);
	assign _1332_ = (_0000_[0] ? \mchip.my_core.Stack.rf[7] [0] : \mchip.my_core.Stack.rf[6] [0]);
	assign _1333_ = (_0000_[1] ? _1332_ : _1331_);
	assign _1334_ = (_0000_[2] ? _1333_ : _1330_);
	assign _1335_ = (_1200_ ? _1327_ : _1334_);
	assign _1336_ = _1170_ | _0890_;
	assign _1337_ = _1336_ | _0889_;
	assign _1338_ = _1337_ | _1173_;
	assign _1339_ = _1338_ | _1124_;
	assign _1340_ = _1180_ | _1077_;
	assign _1341_ = (_0897_ ? _1180_ : _1340_);
	assign _1342_ = \mchip.my_core.Brain.cycle [2] & ~_1341_;
	assign _1343_ = _1339_ & ~_1342_;
	assign _1344_ = \mchip.my_core.Brain.cycle [0] & ~_1337_;
	assign _1345_ = _1343_ & ~_1344_;
	assign _1346_ = _1067_ & ~_1345_;
	assign _1347_ = _1102_ & ~_1147_;
	assign _1348_ = (_1347_ ? \mchip.my_core.rf.rf[7] [0] : \mchip.my_core.rf.rf[6] [0]);
	assign _1349_ = ~(_1147_ | _1122_);
	assign _1350_ = (_1347_ ? \mchip.my_core.rf.rf[5] [0] : \mchip.my_core.rf.rf[4] [0]);
	assign _1351_ = (_1349_ ? _1348_ : _1350_);
	assign _1352_ = _1123_ & ~_1146_;
	assign _1353_ = (_1347_ ? \mchip.my_core.rf.rf[3] [0] : \mchip.my_core.rf.rf[2] [0]);
	assign _1354_ = (_1347_ ? \mchip.my_core.rf.rf[1] [0] : \mchip.my_core.rf.rf[0] [0]);
	assign _1355_ = (_1349_ ? _1353_ : _1354_);
	assign _1356_ = (_1352_ ? _1351_ : _1355_);
	assign _1357_ = _1337_ | _1076_;
	assign _1358_ = \mchip.my_core.Brain.cycle [2] & ~_1357_;
	assign _1359_ = _1126_ & ~_1358_;
	assign _1360_ = _1169_ | ~_0898_;
	assign _1361_ = _1360_ | _1150_;
	assign _1362_ = \mchip.my_core.Brain.cycle [0] & ~_1361_;
	assign _1363_ = _1359_ & ~_1362_;
	assign _1364_ = _1067_ & ~_1363_;
	assign _1365_ = _1039_ & _0680_;
	assign _1366_ = ~_1365_;
	assign _1367_ = _1047_ | ~_1039_;
	assign _1368_ = _1367_ | _0680_;
	assign _1369_ = _1368_ | _0866_;
	assign _1370_ = ~(_1047_ & _1039_);
	assign _1371_ = _1370_ | _0680_;
	assign _1372_ = \mchip.my_core.regA.Q [1] & ~_1371_;
	assign _1373_ = _1369_ & ~_1372_;
	assign _1374_ = _1047_ | _1039_;
	assign _1375_ = _1374_ | _0680_;
	assign _1376_ = \mchip.my_core.regA.Q [7] & ~_1375_;
	assign _1377_ = _1039_ | ~_1047_;
	assign _1378_ = _1377_ | _0680_;
	assign _1379_ = \mchip.my_core.regA.Q [1] & ~_1378_;
	assign _1380_ = _1379_ | _1376_;
	assign _1381_ = _1373_ & ~_1380_;
	assign _1382_ = _1048_ & ~\mchip.my_core.regA.Q [0];
	assign _1383_ = _1381_ & ~_1382_;
	assign _1384_ = _1366_ & ~_1383_;
	assign _1385_ = \mchip.my_core.regA.Q [0] & \mchip.my_core.regB.Q [0];
	assign _1386_ = \mchip.my_core.regA.Q [0] | \mchip.my_core.regB.Q [0];
	assign _1387_ = _1386_ & ~_1385_;
	assign _1388_ = ~_1387_;
	assign _1389_ = _1051_ | _1127_;
	assign _1390_ = _1389_ | _1024_;
	assign _1391_ = _1390_ | _1050_;
	assign _1392_ = _1054_ & ~_1127_;
	assign _1393_ = ~(_1392_ & _1023_);
	assign _1394_ = \mchip.my_core.Brain.cycle [0] & ~_1393_;
	assign _1395_ = _1391_ & ~_1394_;
	assign _1396_ = _1395_ | _1027_;
	assign _1397_ = _1051_ | _1035_;
	assign _1398_ = _1397_ | _1024_;
	assign _1399_ = _1398_ | _1050_;
	assign _1400_ = _1054_ & ~_1035_;
	assign _1401_ = ~(_1400_ & _1023_);
	assign _1402_ = \mchip.my_core.Brain.cycle [0] & ~_1401_;
	assign _1403_ = _1399_ & ~_1402_;
	assign _1404_ = ~(_1403_ | _1027_);
	assign _1405_ = _1051_ | _1040_;
	assign _1406_ = _1405_ | _1024_;
	assign _1407_ = _1406_ | _1050_;
	assign _1408_ = _1054_ & ~_1040_;
	assign _1409_ = ~(_1408_ & _1023_);
	assign _1410_ = \mchip.my_core.Brain.cycle [0] & ~_1409_;
	assign _1411_ = _1407_ & ~_1410_;
	assign _1412_ = ~(_1411_ | _1027_);
	assign _1413_ = _1404_ | ~_1412_;
	assign _1414_ = ~(_1413_ | _1396_);
	assign _1415_ = _1414_ & ~_1388_;
	assign _1416_ = ~(_1412_ & _1404_);
	assign _1417_ = _1416_ | _1396_;
	assign _1418_ = \mchip.my_core.regA.Q [0] & ~_1417_;
	assign _1419_ = ~(_1418_ | _1415_);
	assign _1420_ = _1412_ | _1404_;
	assign _1421_ = ~(_1420_ | _1396_);
	assign _1422_ = _1421_ & _1385_;
	assign _1423_ = _1412_ | ~_1404_;
	assign _1424_ = ~(_1423_ | _1396_);
	assign _1425_ = _1424_ & _1386_;
	assign _1426_ = _1425_ | _1422_;
	assign _1427_ = _1419_ & ~_1426_;
	assign _1428_ = _1396_ & ~_1413_;
	assign _1429_ = _1387_ ^ \mchip.my_core.Unit.flag_reg.Q [0];
	assign _1430_ = _1429_ & _1428_;
	assign _1431_ = _1396_ & ~_1423_;
	assign _1432_ = _1431_ & ~_1388_;
	assign _1433_ = _1396_ & ~_1416_;
	assign _1434_ = _1433_ & _1429_;
	assign _1435_ = _1434_ | _1432_;
	assign _1436_ = _1435_ | _1430_;
	assign _1437_ = _1427_ & ~_1436_;
	assign _1438_ = _1404_ & _1396_;
	assign _1439_ = _1438_ | _1428_;
	assign _1440_ = _1396_ & ~_1439_;
	assign _1441_ = (_1440_ ? _1388_ : _1437_);
	assign _1442_ = ~_1441_;
	assign _1443_ = (_1028_ ? _1384_ : _1442_);
	assign _1444_ = _1228_ | _1173_;
	assign _1445_ = _1444_ | _1124_;
	assign _1446_ = ~(_1151_ | _0980_);
	assign _1447_ = _0906_ | ~_0919_;
	assign _1448_ = _1447_ | _0973_;
	assign _1449_ = _1446_ & ~_1448_;
	assign _1450_ = _1449_ | _1228_;
	assign _1451_ = \mchip.my_core.Brain.cycle [2] & ~_1450_;
	assign _1452_ = _1445_ & ~_1451_;
	assign _1453_ = \mchip.my_core.Brain.cycle [0] & ~_1228_;
	assign _1454_ = _1452_ & ~_1453_;
	assign _1455_ = _1454_ | ~_1067_;
	assign _1456_ = io_in[0] & ~_1455_;
	assign _1457_ = _1173_ | _1024_;
	assign _1458_ = _0901_ & ~_1023_;
	assign _1459_ = (_1458_ ? _0919_ : _1457_);
	assign _1460_ = _1459_ | _1124_;
	assign _1461_ = _1069_ | _1024_;
	assign _1462_ = ~(_1449_ & _0564_);
	assign _1463_ = ~(_1462_ | _0892_);
	assign _1464_ = _1461_ & ~_1463_;
	assign _1465_ = _1171_ | _1023_;
	assign _1466_ = _1465_ | ~_0892_;
	assign _1467_ = ~(_0990_ | _0986_);
	assign _1468_ = (_1466_ ? _1464_ : _1467_);
	assign _1469_ = \mchip.my_core.Brain.cycle [2] & ~_1468_;
	assign _1470_ = _1460_ & ~_1469_;
	assign _1471_ = _1195_ & _1086_;
	assign _1472_ = _1471_ | _1024_;
	assign _1473_ = \mchip.my_core.Brain.cycle [0] & ~_1472_;
	assign _1474_ = _1470_ & ~_1473_;
	assign _1475_ = _1067_ & ~_1474_;
	assign _1476_ = (_1475_ ? \mchip.my_core.regB.Q [0] : _1456_);
	assign _1477_ = _1360_ | _1173_;
	assign _1478_ = _1477_ | _1124_;
	assign _1479_ = _1467_ | _1187_;
	assign _1480_ = \mchip.my_core.Brain.cycle [2] & ~_1479_;
	assign _1481_ = _1478_ & ~_1480_;
	assign _1482_ = _1360_ | _1195_;
	assign _1483_ = \mchip.my_core.Brain.cycle [0] & ~_1482_;
	assign _1484_ = _1481_ & ~_1483_;
	assign _1485_ = _1067_ & ~_1484_;
	assign _1486_ = (_1485_ ? \mchip.my_core.regA.Q [0] : _1476_);
	assign _1487_ = _1360_ | ~_1071_;
	assign _1488_ = \mchip.my_core.Brain.cycle [2] & ~_1487_;
	assign _1489_ = (_1488_ ? \mchip.my_core.Unit.flag_reg.Q [0] : _1486_);
	assign _1490_ = (_1063_ ? _1443_ : _1489_);
	assign _1491_ = (_1364_ ? _1356_ : _1490_);
	assign \mchip.my_core.Stack.bus [0] = (_1346_ ? _1335_ : _1491_);
	assign _1492_ = ~_1334_;
	assign _1493_ = \mchip.my_core.Brain.cycle [0] & ~_1196_;
	assign _1494_ = ~_1493_;
	assign _1495_ = _1494_ & \mchip.my_core.Stack.bus [0];
	assign _1496_ = _1208_ & ~io_in[13];
	assign _1497_ = (_1496_ ? _1334_ : _1495_);
	assign _0023_ = (_1212_ ? _1492_ : _1497_);
	assign _0063_ = (_0000_[0] ? \mchip.my_core.Stack.rf[1] [9] : \mchip.my_core.Stack.rf[0] [9]);
	assign _0064_ = (_0000_[0] ? \mchip.my_core.Stack.rf[3] [9] : \mchip.my_core.Stack.rf[2] [9]);
	assign _0065_ = (_0000_[1] ? _0064_ : _0063_);
	assign _0066_ = (_0000_[0] ? \mchip.my_core.Stack.rf[5] [9] : \mchip.my_core.Stack.rf[4] [9]);
	assign _0067_ = (_0000_[0] ? \mchip.my_core.Stack.rf[7] [9] : \mchip.my_core.Stack.rf[6] [9]);
	assign _0068_ = (_0000_[1] ? _0067_ : _0066_);
	assign _0069_ = (_0000_[2] ? _0068_ : _0065_);
	assign _0070_ = (_0000_[0] ? \mchip.my_core.Stack.rf[1] [1] : \mchip.my_core.Stack.rf[0] [1]);
	assign _0071_ = (_0000_[0] ? \mchip.my_core.Stack.rf[3] [1] : \mchip.my_core.Stack.rf[2] [1]);
	assign _0072_ = (_0000_[1] ? _0071_ : _0070_);
	assign _0073_ = (_0000_[0] ? \mchip.my_core.Stack.rf[5] [1] : \mchip.my_core.Stack.rf[4] [1]);
	assign _0074_ = (_0000_[0] ? \mchip.my_core.Stack.rf[7] [1] : \mchip.my_core.Stack.rf[6] [1]);
	assign _0075_ = (_0000_[1] ? _0074_ : _0073_);
	assign _0076_ = (_0000_[2] ? _0075_ : _0072_);
	assign _0077_ = (_1200_ ? _0069_ : _0076_);
	assign _0078_ = (_1347_ ? \mchip.my_core.rf.rf[7] [1] : \mchip.my_core.rf.rf[6] [1]);
	assign _0079_ = (_1347_ ? \mchip.my_core.rf.rf[5] [1] : \mchip.my_core.rf.rf[4] [1]);
	assign _0080_ = (_1349_ ? _0078_ : _0079_);
	assign _0081_ = (_1347_ ? \mchip.my_core.rf.rf[3] [1] : \mchip.my_core.rf.rf[2] [1]);
	assign _0082_ = (_1347_ ? \mchip.my_core.rf.rf[1] [1] : \mchip.my_core.rf.rf[0] [1]);
	assign _0083_ = (_1349_ ? _0081_ : _0082_);
	assign _0084_ = (_1352_ ? _0080_ : _0083_);
	assign _0085_ = ~\mchip.my_core.regA.Q [2];
	assign _0086_ = _1371_ | _0085_;
	assign _0087_ = \mchip.my_core.regA.Q [0] & ~_1368_;
	assign _0088_ = _0086_ & ~_0087_;
	assign _0089_ = \mchip.my_core.regA.Q [0] & ~_1375_;
	assign _0090_ = \mchip.my_core.regA.Q [2] & ~_1378_;
	assign _0091_ = _0090_ | _0089_;
	assign _0092_ = _0088_ & ~_0091_;
	assign _0093_ = ~\mchip.my_core.regA.Q [1];
	assign _0094_ = _0680_ & ~_1377_;
	assign _0095_ = _0094_ ^ _0093_;
	assign _0096_ = _0095_ ^ \mchip.my_core.regA.Q [0];
	assign _0097_ = _1048_ & ~_0096_;
	assign _0098_ = _0092_ & ~_0097_;
	assign _0099_ = _1366_ & ~_0098_;
	assign _0100_ = \mchip.my_core.regB.Q [1] & \mchip.my_core.regA.Q [1];
	assign _0101_ = ~(\mchip.my_core.regB.Q [1] | \mchip.my_core.regA.Q [1]);
	assign _0102_ = ~(_0101_ | _0100_);
	assign _0103_ = _0102_ ^ _1385_;
	assign _0104_ = _0102_ & _1414_;
	assign _0105_ = \mchip.my_core.regA.Q [1] & ~_1417_;
	assign _0106_ = _0105_ | _0104_;
	assign _0107_ = ~_0100_;
	assign _0108_ = _1421_ & ~_0107_;
	assign _0109_ = _1424_ & ~_0101_;
	assign _0110_ = _0109_ | _0108_;
	assign _0111_ = _0110_ | _0106_;
	assign _0112_ = ~(_1387_ & \mchip.my_core.Unit.flag_reg.Q [0]);
	assign _0113_ = _0103_ ^ _0112_;
	assign _0114_ = _1428_ & ~_0113_;
	assign _0115_ = \mchip.my_core.regB.Q [0] & ~\mchip.my_core.regA.Q [0];
	assign _0116_ = _0115_ ^ _0102_;
	assign _0117_ = ~_0116_;
	assign _0118_ = _1431_ & ~_0117_;
	assign _0119_ = \mchip.my_core.Unit.flag_reg.Q [0] & ~_1387_;
	assign _0120_ = ~(_0119_ ^ _0116_);
	assign _0121_ = _1433_ & ~_0120_;
	assign _0122_ = _0121_ | _0118_;
	assign _0123_ = _0122_ | _0114_;
	assign _0124_ = _0123_ | _0111_;
	assign _0125_ = (_1440_ ? _0103_ : _0124_);
	assign _0126_ = (_1028_ ? _0099_ : _0125_);
	assign _0127_ = io_in[1] & ~_1455_;
	assign _0128_ = (_1475_ ? \mchip.my_core.regB.Q [1] : _0127_);
	assign _0129_ = (_1485_ ? \mchip.my_core.regA.Q [1] : _0128_);
	assign _0130_ = (_1488_ ? \mchip.my_core.Unit.flag_reg.Q [1] : _0129_);
	assign _0131_ = (_1063_ ? _0126_ : _0130_);
	assign _0132_ = (_1364_ ? _0084_ : _0131_);
	assign \mchip.my_core.Stack.bus [1] = (_1346_ ? _0077_ : _0132_);
	assign _0133_ = _0076_ ^ _1334_;
	assign _0134_ = \mchip.my_core.Stack.bus [1] & _1494_;
	assign _0135_ = (_1496_ ? _0076_ : _0134_);
	assign _0028_ = (_1212_ ? _0133_ : _0135_);
	assign _0136_ = (_0000_[0] ? \mchip.my_core.Stack.rf[1] [10] : \mchip.my_core.Stack.rf[0] [10]);
	assign _0137_ = (_0000_[0] ? \mchip.my_core.Stack.rf[3] [10] : \mchip.my_core.Stack.rf[2] [10]);
	assign _0138_ = (_0000_[1] ? _0137_ : _0136_);
	assign _0139_ = (_0000_[0] ? \mchip.my_core.Stack.rf[5] [10] : \mchip.my_core.Stack.rf[4] [10]);
	assign _0140_ = (_0000_[0] ? \mchip.my_core.Stack.rf[7] [10] : \mchip.my_core.Stack.rf[6] [10]);
	assign _0141_ = (_0000_[1] ? _0140_ : _0139_);
	assign _0142_ = (_0000_[2] ? _0141_ : _0138_);
	assign _0143_ = (_0000_[0] ? \mchip.my_core.Stack.rf[1] [2] : \mchip.my_core.Stack.rf[0] [2]);
	assign _0144_ = (_0000_[0] ? \mchip.my_core.Stack.rf[3] [2] : \mchip.my_core.Stack.rf[2] [2]);
	assign _0145_ = (_0000_[1] ? _0144_ : _0143_);
	assign _0146_ = (_0000_[0] ? \mchip.my_core.Stack.rf[5] [2] : \mchip.my_core.Stack.rf[4] [2]);
	assign _0147_ = (_0000_[0] ? \mchip.my_core.Stack.rf[7] [2] : \mchip.my_core.Stack.rf[6] [2]);
	assign _0148_ = (_0000_[1] ? _0147_ : _0146_);
	assign _0149_ = (_0000_[2] ? _0148_ : _0145_);
	assign _0150_ = (_1200_ ? _0142_ : _0149_);
	assign _0151_ = (_1347_ ? \mchip.my_core.rf.rf[7] [2] : \mchip.my_core.rf.rf[6] [2]);
	assign _0152_ = (_1347_ ? \mchip.my_core.rf.rf[5] [2] : \mchip.my_core.rf.rf[4] [2]);
	assign _0153_ = (_1349_ ? _0151_ : _0152_);
	assign _0154_ = (_1347_ ? \mchip.my_core.rf.rf[3] [2] : \mchip.my_core.rf.rf[2] [2]);
	assign _0155_ = (_1347_ ? \mchip.my_core.rf.rf[1] [2] : \mchip.my_core.rf.rf[0] [2]);
	assign _0156_ = (_1349_ ? _0154_ : _0155_);
	assign _0157_ = (_1352_ ? _0153_ : _0156_);
	assign _0158_ = ~\mchip.my_core.regA.Q [3];
	assign _0159_ = _1371_ | _0158_;
	assign _0160_ = \mchip.my_core.regA.Q [1] & ~_1368_;
	assign _0161_ = _0159_ & ~_0160_;
	assign _0162_ = \mchip.my_core.regA.Q [1] & ~_1375_;
	assign _0163_ = \mchip.my_core.regA.Q [3] & ~_1378_;
	assign _0164_ = _0163_ | _0162_;
	assign _0165_ = _0161_ & ~_0164_;
	assign _0166_ = _0094_ & ~_0093_;
	assign _0167_ = \mchip.my_core.regA.Q [0] & ~_0095_;
	assign _0168_ = _0167_ | _0166_;
	assign _0169_ = _0094_ ^ _0085_;
	assign _0170_ = _0169_ ^ _0168_;
	assign _0171_ = _1048_ & ~_0170_;
	assign _0172_ = _0165_ & ~_0171_;
	assign _0173_ = _1366_ & ~_0172_;
	assign _0174_ = _0102_ & _1385_;
	assign _0175_ = _0107_ & ~_0174_;
	assign _0176_ = \mchip.my_core.regB.Q [2] & \mchip.my_core.regA.Q [2];
	assign _0177_ = ~(\mchip.my_core.regB.Q [2] | \mchip.my_core.regA.Q [2]);
	assign _0178_ = ~(_0177_ | _0176_);
	assign _0179_ = ~(_0178_ ^ _0175_);
	assign _0180_ = _0112_ | ~_0103_;
	assign _0181_ = _0179_ ^ _0180_;
	assign _0182_ = _1428_ & ~_0181_;
	assign _0183_ = _0115_ | _0102_;
	assign _0184_ = \mchip.my_core.regA.Q [1] & ~\mchip.my_core.regB.Q [1];
	assign _0185_ = _0183_ & ~_0184_;
	assign _0186_ = _0185_ ^ _0178_;
	assign _0187_ = ~_0186_;
	assign _0188_ = _1431_ & ~_0187_;
	assign _0189_ = _0119_ & ~_0116_;
	assign _0190_ = ~_0189_;
	assign _0191_ = _0190_ ^ _0186_;
	assign _0192_ = _1433_ & ~_0191_;
	assign _0193_ = _0192_ | _0188_;
	assign _0194_ = _0193_ | _0182_;
	assign _0195_ = ~_0176_;
	assign _0196_ = _1421_ & ~_0195_;
	assign _0197_ = _1424_ & ~_0177_;
	assign _0198_ = _0197_ | _0196_;
	assign _0199_ = _0178_ & _1414_;
	assign _0200_ = \mchip.my_core.regA.Q [2] & ~_1417_;
	assign _0201_ = _0200_ | _0199_;
	assign _0202_ = _0201_ | _0198_;
	assign _0203_ = _0202_ | _0194_;
	assign _0204_ = (_1440_ ? _0179_ : _0203_);
	assign _0205_ = (_1028_ ? _0173_ : _0204_);
	assign _0206_ = io_in[2] & ~_1455_;
	assign _0207_ = (_1475_ ? \mchip.my_core.regB.Q [2] : _0206_);
	assign _0208_ = (_1485_ ? \mchip.my_core.regA.Q [2] : _0207_);
	assign _0209_ = (_1488_ ? \mchip.my_core.Unit.flag_reg.Q [2] : _0208_);
	assign _0210_ = (_1063_ ? _0205_ : _0209_);
	assign _0211_ = (_1364_ ? _0157_ : _0210_);
	assign \mchip.my_core.Stack.bus [2] = (_1346_ ? _0150_ : _0211_);
	assign _0212_ = _0076_ & _1334_;
	assign _0213_ = _0212_ ^ _0149_;
	assign _0214_ = \mchip.my_core.Stack.bus [2] & _1494_;
	assign _0215_ = (_1496_ ? _0149_ : _0214_);
	assign _0029_ = (_1212_ ? _0213_ : _0215_);
	assign _0216_ = (_0000_[0] ? \mchip.my_core.Stack.rf[1] [11] : \mchip.my_core.Stack.rf[0] [11]);
	assign _0217_ = (_0000_[0] ? \mchip.my_core.Stack.rf[3] [11] : \mchip.my_core.Stack.rf[2] [11]);
	assign _0218_ = (_0000_[1] ? _0217_ : _0216_);
	assign _0219_ = (_0000_[0] ? \mchip.my_core.Stack.rf[5] [11] : \mchip.my_core.Stack.rf[4] [11]);
	assign _0220_ = (_0000_[0] ? \mchip.my_core.Stack.rf[7] [11] : \mchip.my_core.Stack.rf[6] [11]);
	assign _0221_ = (_0000_[1] ? _0220_ : _0219_);
	assign _0222_ = (_0000_[2] ? _0221_ : _0218_);
	assign _0223_ = (_0000_[0] ? \mchip.my_core.Stack.rf[1] [3] : \mchip.my_core.Stack.rf[0] [3]);
	assign _0224_ = (_0000_[0] ? \mchip.my_core.Stack.rf[3] [3] : \mchip.my_core.Stack.rf[2] [3]);
	assign _0225_ = (_0000_[1] ? _0224_ : _0223_);
	assign _0226_ = (_0000_[0] ? \mchip.my_core.Stack.rf[5] [3] : \mchip.my_core.Stack.rf[4] [3]);
	assign _0227_ = (_0000_[0] ? \mchip.my_core.Stack.rf[7] [3] : \mchip.my_core.Stack.rf[6] [3]);
	assign _0228_ = (_0000_[1] ? _0227_ : _0226_);
	assign _0229_ = (_0000_[2] ? _0228_ : _0225_);
	assign _0230_ = (_1200_ ? _0222_ : _0229_);
	assign _0231_ = (_1347_ ? \mchip.my_core.rf.rf[7] [3] : \mchip.my_core.rf.rf[6] [3]);
	assign _0232_ = (_1347_ ? \mchip.my_core.rf.rf[5] [3] : \mchip.my_core.rf.rf[4] [3]);
	assign _0233_ = (_1349_ ? _0231_ : _0232_);
	assign _0234_ = (_1347_ ? \mchip.my_core.rf.rf[3] [3] : \mchip.my_core.rf.rf[2] [3]);
	assign _0235_ = (_1347_ ? \mchip.my_core.rf.rf[1] [3] : \mchip.my_core.rf.rf[0] [3]);
	assign _0236_ = (_1349_ ? _0234_ : _0235_);
	assign _0237_ = (_1352_ ? _0233_ : _0236_);
	assign _0238_ = ~\mchip.my_core.regA.Q [4];
	assign _0239_ = _1371_ | _0238_;
	assign _0240_ = \mchip.my_core.regA.Q [2] & ~_1368_;
	assign _0241_ = _0239_ & ~_0240_;
	assign _0242_ = \mchip.my_core.regA.Q [2] & ~_1375_;
	assign _0243_ = \mchip.my_core.regA.Q [4] & ~_1378_;
	assign _0244_ = _0243_ | _0242_;
	assign _0245_ = _0241_ & ~_0244_;
	assign _0246_ = _0094_ & ~_0085_;
	assign _0247_ = _0168_ & ~_0169_;
	assign _0248_ = _0247_ | _0246_;
	assign _0249_ = _0094_ ^ _0158_;
	assign _0250_ = _0249_ ^ _0248_;
	assign _0251_ = _1048_ & ~_0250_;
	assign _0252_ = _0245_ & ~_0251_;
	assign _0253_ = _1366_ & ~_0252_;
	assign _0254_ = ~(\mchip.my_core.regB.Q [3] & \mchip.my_core.regA.Q [3]);
	assign _0255_ = ~(\mchip.my_core.regB.Q [3] | \mchip.my_core.regA.Q [3]);
	assign _0256_ = _0254_ & ~_0255_;
	assign _0257_ = ~_0256_;
	assign _0258_ = _0178_ & ~_0175_;
	assign _0259_ = _0195_ & ~_0258_;
	assign _0260_ = _0259_ ^ _0257_;
	assign _0261_ = ~_0260_;
	assign _0262_ = _1414_ & ~_0257_;
	assign _0263_ = \mchip.my_core.regA.Q [3] & ~_1417_;
	assign _0264_ = ~(_0263_ | _0262_);
	assign _0265_ = _1421_ & ~_0254_;
	assign _0266_ = _1424_ & ~_0255_;
	assign _0267_ = _0266_ | _0265_;
	assign _0268_ = _0264_ & ~_0267_;
	assign _0269_ = _0180_ | ~_0179_;
	assign _0270_ = _0260_ ^ _0269_;
	assign _0271_ = _1428_ & ~_0270_;
	assign _0272_ = _0185_ | _0178_;
	assign _0273_ = \mchip.my_core.regA.Q [2] & ~\mchip.my_core.regB.Q [2];
	assign _0274_ = _0272_ & ~_0273_;
	assign _0275_ = _0274_ ^ _0256_;
	assign _0276_ = ~_0275_;
	assign _0277_ = _1431_ & ~_0276_;
	assign _0278_ = _0190_ | _0186_;
	assign _0279_ = _0278_ ^ _0275_;
	assign _0280_ = _1433_ & ~_0279_;
	assign _0281_ = _0280_ | _0277_;
	assign _0282_ = _0281_ | _0271_;
	assign _0283_ = _0268_ & ~_0282_;
	assign _0284_ = (_1440_ ? _0261_ : _0283_);
	assign _0285_ = ~_0284_;
	assign _0286_ = (_1028_ ? _0253_ : _0285_);
	assign _0287_ = io_in[3] & ~_1455_;
	assign _0288_ = (_1475_ ? \mchip.my_core.regB.Q [3] : _0287_);
	assign _0289_ = (_1485_ ? \mchip.my_core.regA.Q [3] : _0288_);
	assign _0290_ = (_1488_ ? \mchip.my_core.Unit.flag_reg.Q [3] : _0289_);
	assign _0291_ = (_1063_ ? _0286_ : _0290_);
	assign _0292_ = (_1364_ ? _0237_ : _0291_);
	assign \mchip.my_core.Stack.bus [3] = (_1346_ ? _0230_ : _0292_);
	assign _0293_ = _0212_ & _0149_;
	assign _0294_ = _0293_ ^ _0229_;
	assign _0295_ = (_1496_ ? _0229_ : \mchip.my_core.Stack.bus [3]);
	assign _0030_ = (_1212_ ? _0294_ : _0295_);
	assign _0296_ = (_0000_[0] ? \mchip.my_core.Stack.rf[1] [12] : \mchip.my_core.Stack.rf[0] [12]);
	assign _0297_ = (_0000_[0] ? \mchip.my_core.Stack.rf[3] [12] : \mchip.my_core.Stack.rf[2] [12]);
	assign _0298_ = (_0000_[1] ? _0297_ : _0296_);
	assign _0299_ = (_0000_[0] ? \mchip.my_core.Stack.rf[5] [12] : \mchip.my_core.Stack.rf[4] [12]);
	assign _0300_ = (_0000_[0] ? \mchip.my_core.Stack.rf[7] [12] : \mchip.my_core.Stack.rf[6] [12]);
	assign _0301_ = (_0000_[1] ? _0300_ : _0299_);
	assign _0302_ = (_0000_[2] ? _0301_ : _0298_);
	assign _0303_ = (_0000_[0] ? \mchip.my_core.Stack.rf[1] [4] : \mchip.my_core.Stack.rf[0] [4]);
	assign _0304_ = (_0000_[0] ? \mchip.my_core.Stack.rf[3] [4] : \mchip.my_core.Stack.rf[2] [4]);
	assign _0305_ = (_0000_[1] ? _0304_ : _0303_);
	assign _0306_ = (_0000_[0] ? \mchip.my_core.Stack.rf[5] [4] : \mchip.my_core.Stack.rf[4] [4]);
	assign _0307_ = (_0000_[0] ? \mchip.my_core.Stack.rf[7] [4] : \mchip.my_core.Stack.rf[6] [4]);
	assign _0308_ = (_0000_[1] ? _0307_ : _0306_);
	assign _0309_ = (_0000_[2] ? _0308_ : _0305_);
	assign _0310_ = (_1200_ ? _0302_ : _0309_);
	assign _0311_ = (_1347_ ? \mchip.my_core.rf.rf[7] [4] : \mchip.my_core.rf.rf[6] [4]);
	assign _0312_ = (_1347_ ? \mchip.my_core.rf.rf[5] [4] : \mchip.my_core.rf.rf[4] [4]);
	assign _0313_ = (_1349_ ? _0311_ : _0312_);
	assign _0314_ = (_1347_ ? \mchip.my_core.rf.rf[3] [4] : \mchip.my_core.rf.rf[2] [4]);
	assign _0315_ = (_1347_ ? \mchip.my_core.rf.rf[1] [4] : \mchip.my_core.rf.rf[0] [4]);
	assign _0316_ = (_1349_ ? _0314_ : _0315_);
	assign _0317_ = (_1352_ ? _0313_ : _0316_);
	assign _0318_ = ~\mchip.my_core.regA.Q [5];
	assign _0319_ = _1371_ | _0318_;
	assign _0320_ = \mchip.my_core.regA.Q [3] & ~_1368_;
	assign _0321_ = _0319_ & ~_0320_;
	assign _0322_ = \mchip.my_core.regA.Q [3] & ~_1375_;
	assign _0323_ = \mchip.my_core.regA.Q [5] & ~_1378_;
	assign _0324_ = _0323_ | _0322_;
	assign _0325_ = _0321_ & ~_0324_;
	assign _0326_ = _0094_ & ~_0158_;
	assign _0327_ = _0246_ & ~_0249_;
	assign _0328_ = _0327_ | _0326_;
	assign _0329_ = _0249_ | _0169_;
	assign _0330_ = _0168_ & ~_0329_;
	assign _0331_ = _0330_ | _0328_;
	assign _0332_ = _0094_ ^ _0238_;
	assign _0333_ = _0332_ ^ _0331_;
	assign _0334_ = _1048_ & ~_0333_;
	assign _0335_ = _0325_ & ~_0334_;
	assign _0336_ = _1366_ & ~_0335_;
	assign _0337_ = \mchip.my_core.regB.Q [4] & \mchip.my_core.regA.Q [4];
	assign _0338_ = ~(\mchip.my_core.regB.Q [4] | \mchip.my_core.regA.Q [4]);
	assign _0339_ = ~(_0338_ | _0337_);
	assign _0340_ = ~_0339_;
	assign _0341_ = _0256_ & ~_0195_;
	assign _0342_ = _0254_ & ~_0341_;
	assign _0343_ = _0256_ & _0178_;
	assign _0344_ = _0343_ & ~_0175_;
	assign _0345_ = _0342_ & ~_0344_;
	assign _0346_ = _0345_ ^ _0340_;
	assign _0347_ = ~_0346_;
	assign _0348_ = _1414_ & ~_0340_;
	assign _0349_ = \mchip.my_core.regA.Q [4] & ~_1417_;
	assign _0350_ = ~(_0349_ | _0348_);
	assign _0351_ = ~_0337_;
	assign _0352_ = _1421_ & ~_0351_;
	assign _0353_ = _1424_ & ~_0338_;
	assign _0354_ = _0353_ | _0352_;
	assign _0355_ = _0350_ & ~_0354_;
	assign _0356_ = ~(_0260_ & _0179_);
	assign _0357_ = _0356_ | _0180_;
	assign _0358_ = ~(_0347_ ^ _0357_);
	assign _0359_ = _1428_ & ~_0358_;
	assign _0360_ = \mchip.my_core.regB.Q [3] | ~\mchip.my_core.regA.Q [3];
	assign _0361_ = _0273_ & ~_0256_;
	assign _0362_ = _0360_ & ~_0361_;
	assign _0363_ = _0256_ | _0178_;
	assign _0364_ = ~(_0363_ | _0185_);
	assign _0365_ = _0362_ & ~_0364_;
	assign _0366_ = _0365_ ^ _0339_;
	assign _0367_ = ~_0366_;
	assign _0368_ = _1431_ & ~_0367_;
	assign _0369_ = _0275_ | _0186_;
	assign _0370_ = _0189_ & ~_0369_;
	assign _0371_ = _0370_ ^ _0367_;
	assign _0372_ = _1433_ & ~_0371_;
	assign _0373_ = _0372_ | _0368_;
	assign _0374_ = _0373_ | _0359_;
	assign _0375_ = _0355_ & ~_0374_;
	assign _0376_ = (_1440_ ? _0347_ : _0375_);
	assign _0377_ = ~_0376_;
	assign _0378_ = (_1028_ ? _0336_ : _0377_);
	assign _0379_ = io_in[4] & ~_1455_;
	assign _0380_ = (_1475_ ? \mchip.my_core.regB.Q [4] : _0379_);
	assign _0381_ = (_1485_ ? \mchip.my_core.regA.Q [4] : _0380_);
	assign _0382_ = _0381_ & ~_1488_;
	assign _0383_ = (_1063_ ? _0378_ : _0382_);
	assign _0384_ = (_1364_ ? _0317_ : _0383_);
	assign \mchip.my_core.Stack.bus [4] = (_1346_ ? _0310_ : _0384_);
	assign _0385_ = ~(_0229_ & _0149_);
	assign _0386_ = _0212_ & ~_0385_;
	assign _0387_ = _0386_ ^ _0309_;
	assign _0388_ = (_1496_ ? _0309_ : \mchip.my_core.Stack.bus [4]);
	assign _0031_ = (_1212_ ? _0387_ : _0388_);
	assign _0389_ = (_0000_[0] ? \mchip.my_core.Stack.rf[1] [13] : \mchip.my_core.Stack.rf[0] [13]);
	assign _0390_ = (_0000_[0] ? \mchip.my_core.Stack.rf[3] [13] : \mchip.my_core.Stack.rf[2] [13]);
	assign _0391_ = (_0000_[1] ? _0390_ : _0389_);
	assign _0392_ = (_0000_[0] ? \mchip.my_core.Stack.rf[5] [13] : \mchip.my_core.Stack.rf[4] [13]);
	assign _0393_ = (_0000_[0] ? \mchip.my_core.Stack.rf[7] [13] : \mchip.my_core.Stack.rf[6] [13]);
	assign _0394_ = (_0000_[1] ? _0393_ : _0392_);
	assign _0395_ = (_0000_[2] ? _0394_ : _0391_);
	assign _0396_ = (_0000_[0] ? \mchip.my_core.Stack.rf[1] [5] : \mchip.my_core.Stack.rf[0] [5]);
	assign _0397_ = (_0000_[0] ? \mchip.my_core.Stack.rf[3] [5] : \mchip.my_core.Stack.rf[2] [5]);
	assign _0398_ = (_0000_[1] ? _0397_ : _0396_);
	assign _0399_ = (_0000_[0] ? \mchip.my_core.Stack.rf[5] [5] : \mchip.my_core.Stack.rf[4] [5]);
	assign _0400_ = (_0000_[0] ? \mchip.my_core.Stack.rf[7] [5] : \mchip.my_core.Stack.rf[6] [5]);
	assign _0401_ = (_0000_[1] ? _0400_ : _0399_);
	assign _0402_ = (_0000_[2] ? _0401_ : _0398_);
	assign _0403_ = (_1200_ ? _0395_ : _0402_);
	assign _0404_ = (_1347_ ? \mchip.my_core.rf.rf[7] [5] : \mchip.my_core.rf.rf[6] [5]);
	assign _0405_ = (_1347_ ? \mchip.my_core.rf.rf[5] [5] : \mchip.my_core.rf.rf[4] [5]);
	assign _0406_ = (_1349_ ? _0404_ : _0405_);
	assign _0407_ = (_1347_ ? \mchip.my_core.rf.rf[3] [5] : \mchip.my_core.rf.rf[2] [5]);
	assign _0408_ = (_1347_ ? \mchip.my_core.rf.rf[1] [5] : \mchip.my_core.rf.rf[0] [5]);
	assign _0409_ = (_1349_ ? _0407_ : _0408_);
	assign _0410_ = (_1352_ ? _0406_ : _0409_);
	assign _0411_ = ~\mchip.my_core.regA.Q [6];
	assign _0412_ = _1371_ | _0411_;
	assign _0413_ = \mchip.my_core.regA.Q [4] & ~_1368_;
	assign _0414_ = _0412_ & ~_0413_;
	assign _0415_ = \mchip.my_core.regA.Q [4] & ~_1375_;
	assign _0416_ = \mchip.my_core.regA.Q [6] & ~_1378_;
	assign _0417_ = _0416_ | _0415_;
	assign _0418_ = _0414_ & ~_0417_;
	assign _0419_ = _0094_ & ~_0238_;
	assign _0420_ = _0331_ & ~_0332_;
	assign _0421_ = _0420_ | _0419_;
	assign _0422_ = _0094_ ^ _0318_;
	assign _0423_ = _0422_ ^ _0421_;
	assign _0424_ = _1048_ & ~_0423_;
	assign _0425_ = _0418_ & ~_0424_;
	assign _0426_ = _1366_ & ~_0425_;
	assign _0427_ = ~(\mchip.my_core.regB.Q [5] & \mchip.my_core.regA.Q [5]);
	assign _0428_ = ~(\mchip.my_core.regB.Q [5] | \mchip.my_core.regA.Q [5]);
	assign _0429_ = _0427_ & ~_0428_;
	assign _0430_ = ~_0429_;
	assign _0431_ = _0339_ & ~_0345_;
	assign _0432_ = _0351_ & ~_0431_;
	assign _0433_ = _0432_ ^ _0430_;
	assign _0434_ = _1414_ & ~_0430_;
	assign _0435_ = \mchip.my_core.regA.Q [5] & ~_1417_;
	assign _0436_ = _0435_ | _0434_;
	assign _0437_ = _1421_ & ~_0427_;
	assign _0438_ = _1424_ & ~_0428_;
	assign _0439_ = _0438_ | _0437_;
	assign _0440_ = _0439_ | _0436_;
	assign _0441_ = _0347_ | _0357_;
	assign _0442_ = _0433_ ^ _0441_;
	assign _0443_ = _1428_ & ~_0442_;
	assign _0444_ = _0365_ | _0339_;
	assign _0445_ = \mchip.my_core.regA.Q [4] & ~\mchip.my_core.regB.Q [4];
	assign _0446_ = _0444_ & ~_0445_;
	assign _0447_ = _0446_ ^ _0429_;
	assign _0448_ = ~_0447_;
	assign _0449_ = _1431_ & ~_0448_;
	assign _0450_ = _0370_ & ~_0366_;
	assign _0451_ = _0450_ ^ _0448_;
	assign _0452_ = _1433_ & ~_0451_;
	assign _0453_ = _0452_ | _0449_;
	assign _0454_ = _0453_ | _0443_;
	assign _0455_ = _0454_ | _0440_;
	assign _0456_ = (_1440_ ? _0433_ : _0455_);
	assign _0457_ = (_1028_ ? _0426_ : _0456_);
	assign _0458_ = io_in[5] & ~_1455_;
	assign _0459_ = (_1475_ ? \mchip.my_core.regB.Q [5] : _0458_);
	assign _0460_ = (_1485_ ? \mchip.my_core.regA.Q [5] : _0459_);
	assign _0461_ = _0460_ & ~_1488_;
	assign _0462_ = (_1063_ ? _0457_ : _0461_);
	assign _0463_ = (_1364_ ? _0410_ : _0462_);
	assign \mchip.my_core.Stack.bus [5] = (_1346_ ? _0403_ : _0463_);
	assign _0464_ = _0386_ & _0309_;
	assign _0465_ = _0464_ ^ _0402_;
	assign _0466_ = (_1496_ ? _0402_ : \mchip.my_core.Stack.bus [5]);
	assign _0032_ = (_1212_ ? _0465_ : _0466_);
	assign _0467_ = _1173_ & _0919_;
	assign _0468_ = _0467_ | _1172_;
	assign _0469_ = _0468_ | _1124_;
	assign _0470_ = _1180_ & _1076_;
	assign _0471_ = _0470_ | _1172_;
	assign _0472_ = \mchip.my_core.Brain.cycle [2] & ~_0471_;
	assign _0473_ = _0469_ & ~_0472_;
	assign _0474_ = _1065_ & ~_0473_;
	assign _0475_ = (_0000_[0] ? \mchip.my_core.Stack.rf[1] [6] : \mchip.my_core.Stack.rf[0] [6]);
	assign _0476_ = (_0000_[0] ? \mchip.my_core.Stack.rf[3] [6] : \mchip.my_core.Stack.rf[2] [6]);
	assign _0477_ = (_0000_[1] ? _0476_ : _0475_);
	assign _0478_ = (_0000_[0] ? \mchip.my_core.Stack.rf[5] [6] : \mchip.my_core.Stack.rf[4] [6]);
	assign _0479_ = (_0000_[0] ? \mchip.my_core.Stack.rf[7] [6] : \mchip.my_core.Stack.rf[6] [6]);
	assign _0480_ = (_0000_[1] ? _0479_ : _0478_);
	assign _0481_ = (_0000_[2] ? _0480_ : _0477_);
	assign _0482_ = (_1200_ ? _0474_ : _0481_);
	assign _0483_ = (_1347_ ? \mchip.my_core.rf.rf[7] [6] : \mchip.my_core.rf.rf[6] [6]);
	assign _0484_ = (_1347_ ? \mchip.my_core.rf.rf[5] [6] : \mchip.my_core.rf.rf[4] [6]);
	assign _0485_ = (_1349_ ? _0483_ : _0484_);
	assign _0486_ = (_1347_ ? \mchip.my_core.rf.rf[3] [6] : \mchip.my_core.rf.rf[2] [6]);
	assign _0487_ = (_1347_ ? \mchip.my_core.rf.rf[1] [6] : \mchip.my_core.rf.rf[0] [6]);
	assign _0488_ = (_1349_ ? _0486_ : _0487_);
	assign _0489_ = (_1352_ ? _0485_ : _0488_);
	assign _0490_ = _0489_ | _0474_;
	assign _0491_ = ~\mchip.my_core.regA.Q [7];
	assign _0492_ = _1371_ | _0491_;
	assign _0493_ = \mchip.my_core.regA.Q [5] & ~_1368_;
	assign _0494_ = _0492_ & ~_0493_;
	assign _0495_ = \mchip.my_core.regA.Q [5] & ~_1375_;
	assign _0496_ = \mchip.my_core.regA.Q [7] & ~_1378_;
	assign _0497_ = _0496_ | _0495_;
	assign _0498_ = _0494_ & ~_0497_;
	assign _0499_ = _0094_ & ~_0318_;
	assign _0500_ = _0419_ & ~_0422_;
	assign _0501_ = _0500_ | _0499_;
	assign _0502_ = _0422_ | _0332_;
	assign _0503_ = _0331_ & ~_0502_;
	assign _0504_ = _0503_ | _0501_;
	assign _0505_ = _0094_ ^ _0411_;
	assign _0506_ = _0505_ ^ _0504_;
	assign _0507_ = _1048_ & ~_0506_;
	assign _0508_ = _0498_ & ~_0507_;
	assign _0509_ = _1366_ & ~_0508_;
	assign _0510_ = _0429_ & ~_0351_;
	assign _0511_ = _0510_ | ~_0427_;
	assign _0512_ = ~(_0429_ & _0339_);
	assign _0513_ = ~(_0512_ | _0345_);
	assign _0514_ = _0513_ | _0511_;
	assign _0515_ = \mchip.my_core.regB.Q [6] & \mchip.my_core.regA.Q [6];
	assign _0516_ = ~(\mchip.my_core.regB.Q [6] | \mchip.my_core.regA.Q [6]);
	assign _0517_ = ~(_0516_ | _0515_);
	assign _0518_ = _0517_ ^ _0514_;
	assign _0519_ = ~(_0433_ & _0346_);
	assign _0520_ = _0519_ | _0357_;
	assign _0521_ = ~_0518_;
	assign _0522_ = ~(_0521_ ^ _0520_);
	assign _0523_ = _1428_ & ~_0522_;
	assign _0524_ = _0445_ & ~_0429_;
	assign _0525_ = \mchip.my_core.regA.Q [5] & ~\mchip.my_core.regB.Q [5];
	assign _0526_ = ~(_0525_ | _0524_);
	assign _0527_ = _0429_ | _0339_;
	assign _0528_ = ~(_0527_ | _0365_);
	assign _0529_ = _0526_ & ~_0528_;
	assign _0530_ = _0529_ ^ _0517_;
	assign _0531_ = ~_0530_;
	assign _0532_ = _1431_ & ~_0531_;
	assign _0533_ = _0447_ | _0366_;
	assign _0534_ = _0370_ & ~_0533_;
	assign _0535_ = _0534_ ^ _0531_;
	assign _0536_ = _1433_ & ~_0535_;
	assign _0537_ = _0536_ | _0532_;
	assign _0538_ = _0537_ | _0523_;
	assign _0539_ = ~_0515_;
	assign _0540_ = _1421_ & ~_0539_;
	assign _0541_ = _1424_ & ~_0516_;
	assign _0542_ = _0541_ | _0540_;
	assign _0543_ = _0517_ & _1414_;
	assign _0544_ = \mchip.my_core.regA.Q [6] & ~_1417_;
	assign _0545_ = _0544_ | _0543_;
	assign _0546_ = _0545_ | _0542_;
	assign _0547_ = _0546_ | _0538_;
	assign _0548_ = (_1440_ ? _0518_ : _0547_);
	assign _0549_ = (_1028_ ? _0509_ : _0548_);
	assign _0550_ = _1455_ | ~io_in[6];
	assign _0551_ = ~(_0474_ | \mchip.my_core.regB.Q [6]);
	assign _0552_ = (_1475_ ? _0551_ : _0550_);
	assign _0553_ = (_1485_ ? _0411_ : _0552_);
	assign _0554_ = ~(_0553_ | _1488_);
	assign _0555_ = (_1063_ ? _0549_ : _0554_);
	assign _0556_ = (_1364_ ? _0490_ : _0555_);
	assign \mchip.my_core.Stack.bus [6] = (_1346_ ? _0482_ : _0556_);
	assign _0557_ = ~(_0402_ & _0309_);
	assign _0558_ = _0386_ & ~_0557_;
	assign _0559_ = _0558_ ^ _0481_;
	assign _0560_ = \mchip.my_core.Stack.bus [6] & _1494_;
	assign _0561_ = (_1496_ ? _0481_ : _0560_);
	assign _0033_ = (_1212_ ? _0559_ : _0561_);
	assign _0562_ = _1172_ | _0919_;
	assign _0563_ = _0562_ | _1124_;
	assign _0565_ = _1467_ & ~_0564_;
	assign _0566_ = ~(_1467_ & _1076_);
	assign _0567_ = _1180_ & ~_0566_;
	assign _0568_ = _0567_ | _0565_;
	assign _0569_ = _0568_ | _1172_;
	assign _0570_ = \mchip.my_core.Brain.cycle [2] & ~_0569_;
	assign _0571_ = _0563_ & ~_0570_;
	assign _0572_ = _1065_ & ~_0571_;
	assign _0573_ = (_0000_[0] ? \mchip.my_core.Stack.rf[1] [7] : \mchip.my_core.Stack.rf[0] [7]);
	assign _0574_ = (_0000_[0] ? \mchip.my_core.Stack.rf[3] [7] : \mchip.my_core.Stack.rf[2] [7]);
	assign _0575_ = (_0000_[1] ? _0574_ : _0573_);
	assign _0576_ = (_0000_[0] ? \mchip.my_core.Stack.rf[5] [7] : \mchip.my_core.Stack.rf[4] [7]);
	assign _0577_ = (_0000_[0] ? \mchip.my_core.Stack.rf[7] [7] : \mchip.my_core.Stack.rf[6] [7]);
	assign _0578_ = (_0000_[1] ? _0577_ : _0576_);
	assign _0579_ = (_0000_[2] ? _0578_ : _0575_);
	assign _0580_ = (_1200_ ? _0572_ : _0579_);
	assign _0581_ = (_1347_ ? \mchip.my_core.rf.rf[7] [7] : \mchip.my_core.rf.rf[6] [7]);
	assign _0582_ = (_1347_ ? \mchip.my_core.rf.rf[5] [7] : \mchip.my_core.rf.rf[4] [7]);
	assign _0583_ = (_1349_ ? _0581_ : _0582_);
	assign _0584_ = (_1347_ ? \mchip.my_core.rf.rf[3] [7] : \mchip.my_core.rf.rf[2] [7]);
	assign _0585_ = (_1347_ ? \mchip.my_core.rf.rf[1] [7] : \mchip.my_core.rf.rf[0] [7]);
	assign _0586_ = (_1349_ ? _0584_ : _0585_);
	assign _0587_ = (_1352_ ? _0583_ : _0586_);
	assign _0588_ = _0587_ | _0572_;
	assign _0589_ = _1371_ | _0866_;
	assign _0590_ = \mchip.my_core.regA.Q [6] & ~_1368_;
	assign _0591_ = _0589_ & ~_0590_;
	assign _0592_ = \mchip.my_core.regA.Q [6] & ~_1375_;
	assign _0593_ = \mchip.my_core.regA.Q [0] & ~_1378_;
	assign _0594_ = _0593_ | _0592_;
	assign _0595_ = _0591_ & ~_0594_;
	assign _0596_ = _0504_ & ~_0505_;
	assign _0597_ = _0094_ & ~_0411_;
	assign _0598_ = _0597_ | _0596_;
	assign _0599_ = _0094_ ^ _0491_;
	assign _0600_ = _0599_ ^ _0598_;
	assign _0601_ = _1048_ & ~_0600_;
	assign _0602_ = _0595_ & ~_0601_;
	assign _0603_ = _1366_ & ~_0602_;
	assign _0604_ = _0517_ & _0514_;
	assign _0605_ = _0539_ & ~_0604_;
	assign _0606_ = ~(\mchip.my_core.regB.Q [7] & \mchip.my_core.regA.Q [7]);
	assign _0607_ = ~(\mchip.my_core.regB.Q [7] | \mchip.my_core.regA.Q [7]);
	assign _0608_ = _0606_ & ~_0607_;
	assign _0609_ = ~_0608_;
	assign _0610_ = _0609_ ^ _0605_;
	assign _0611_ = _0521_ | _0520_;
	assign _0612_ = _0610_ ^ _0611_;
	assign _0613_ = _1428_ & ~_0612_;
	assign _0614_ = _0529_ | _0517_;
	assign _0615_ = \mchip.my_core.regA.Q [6] & ~\mchip.my_core.regB.Q [6];
	assign _0616_ = _0614_ & ~_0615_;
	assign _0617_ = _0616_ ^ _0608_;
	assign _0618_ = _0617_ & _1431_;
	assign _0619_ = ~(_0534_ & _0531_);
	assign _0620_ = _0619_ ^ _0617_;
	assign _0621_ = _1433_ & ~_0620_;
	assign _0622_ = _0621_ | _0618_;
	assign _0623_ = _0622_ | _0613_;
	assign _0624_ = _1421_ & ~_0606_;
	assign _0625_ = _1424_ & ~_0607_;
	assign _0626_ = _0625_ | _0624_;
	assign _0627_ = _1414_ & ~_0609_;
	assign _0628_ = \mchip.my_core.regA.Q [7] & ~_1417_;
	assign _0629_ = _0628_ | _0627_;
	assign _0630_ = _0629_ | _0626_;
	assign _0631_ = _0630_ | _0623_;
	assign _0632_ = (_1440_ ? _0610_ : _0631_);
	assign _0633_ = (_1028_ ? _0603_ : _0632_);
	assign _0634_ = _1455_ | ~io_in[7];
	assign _0635_ = ~(_0572_ | \mchip.my_core.regB.Q [7]);
	assign _0636_ = (_1475_ ? _0635_ : _0634_);
	assign _0637_ = (_1485_ ? _0491_ : _0636_);
	assign _0638_ = ~(_0637_ | _1488_);
	assign _0639_ = (_1063_ ? _0633_ : _0638_);
	assign _0640_ = (_1364_ ? _0588_ : _0639_);
	assign \mchip.my_core.Stack.bus [7] = (_1346_ ? _0580_ : _0640_);
	assign _0641_ = _0558_ & _0481_;
	assign _0642_ = _0641_ ^ _0579_;
	assign _0643_ = \mchip.my_core.Stack.bus [7] & _1494_;
	assign _0644_ = (_1496_ ? _0579_ : _0643_);
	assign _0034_ = (_1212_ ? _0642_ : _0644_);
	assign _0645_ = ~(_0579_ & _0481_);
	assign _0646_ = _0645_ | _0557_;
	assign _0647_ = _0386_ & ~_0646_;
	assign _0648_ = _0647_ ^ _1327_;
	assign _0649_ = _1327_ & ~_1493_;
	assign _0650_ = (_1496_ ? \mchip.my_core.Stack.bus [0] : _0649_);
	assign _0035_ = (_1212_ ? _0648_ : _0650_);
	assign _0651_ = _0647_ & _1327_;
	assign _0652_ = _0651_ ^ _0069_;
	assign _0653_ = _0069_ & ~_1493_;
	assign _0654_ = (_1496_ ? \mchip.my_core.Stack.bus [1] : _0653_);
	assign _0036_ = (_1212_ ? _0652_ : _0654_);
	assign _0655_ = ~(_0069_ & _1327_);
	assign _0656_ = _0647_ & ~_0655_;
	assign _0657_ = _0656_ ^ _0142_;
	assign _0658_ = _0142_ & ~_1493_;
	assign _0659_ = (_1496_ ? \mchip.my_core.Stack.bus [2] : _0658_);
	assign _0024_ = (_1212_ ? _0657_ : _0659_);
	assign _0660_ = _0656_ & _0142_;
	assign _0661_ = _0660_ ^ _0222_;
	assign _0662_ = _0222_ & ~_1493_;
	assign _0663_ = (_1496_ ? \mchip.my_core.Stack.bus [3] : _0662_);
	assign _0025_ = (_1212_ ? _0661_ : _0663_);
	assign _0664_ = ~(_0222_ & _0142_);
	assign _0665_ = _0664_ | _0655_;
	assign _0666_ = _0647_ & ~_0665_;
	assign _0667_ = _0666_ ^ _0302_;
	assign _0668_ = _0302_ & ~_1493_;
	assign _0669_ = (_1496_ ? \mchip.my_core.Stack.bus [4] : _0668_);
	assign _0026_ = (_1212_ ? _0667_ : _0669_);
	assign _0670_ = _0666_ & _0302_;
	assign _0671_ = _0670_ ^ _0395_;
	assign _0672_ = _0395_ & ~_1493_;
	assign _0673_ = (_1496_ ? \mchip.my_core.Stack.bus [5] : _0672_);
	assign _0027_ = (_1212_ ? _0671_ : _0673_);
	assign _0674_ = _0897_ & ~_1064_;
	assign \mchip.my_core.regA.d [0] = (_0674_ ? \mchip.my_core.rf.rf[0] [0] : \mchip.my_core.Stack.bus [0]);
	assign \mchip.my_core.regA.d [1] = (_0674_ ? \mchip.my_core.rf.rf[0] [1] : \mchip.my_core.Stack.bus [1]);
	assign \mchip.my_core.regA.d [2] = (_0674_ ? \mchip.my_core.rf.rf[0] [2] : \mchip.my_core.Stack.bus [2]);
	assign \mchip.my_core.regA.d [3] = (_0674_ ? \mchip.my_core.rf.rf[0] [3] : \mchip.my_core.Stack.bus [3]);
	assign \mchip.my_core.regA.d [4] = (_0674_ ? \mchip.my_core.rf.rf[0] [4] : \mchip.my_core.Stack.bus [4]);
	assign \mchip.my_core.regA.d [5] = (_0674_ ? \mchip.my_core.rf.rf[0] [5] : \mchip.my_core.Stack.bus [5]);
	assign \mchip.my_core.regA.d [6] = (_0674_ ? \mchip.my_core.rf.rf[0] [6] : \mchip.my_core.Stack.bus [6]);
	assign \mchip.my_core.regA.d [7] = (_0674_ ? \mchip.my_core.rf.rf[0] [7] : \mchip.my_core.Stack.bus [7]);
	assign _0675_ = _1368_ & _1375_;
	assign _0676_ = \mchip.my_core.regA.Q [7] & ~_0675_;
	assign _0677_ = _1371_ & _1378_;
	assign _0678_ = \mchip.my_core.regA.Q [0] & ~_0677_;
	assign _0679_ = _0678_ | _0676_;
	assign _0681_ = _0679_ & ~_0680_;
	assign _0682_ = _0608_ & ~_0539_;
	assign _0683_ = _0606_ & ~_0682_;
	assign _0684_ = ~(_0608_ & _0517_);
	assign _0685_ = _0511_ & ~_0684_;
	assign _0686_ = _0683_ & ~_0685_;
	assign _0687_ = _0684_ | _0512_;
	assign _0688_ = ~(_0687_ | _0345_);
	assign _0689_ = _0686_ & ~_0688_;
	assign _0690_ = ~_0689_;
	assign _0691_ = ~(_0610_ & _0518_);
	assign _0692_ = _0691_ | _0519_;
	assign _0693_ = ~(_0692_ | _0357_);
	assign _0694_ = _0689_ ^ _0693_;
	assign _0695_ = _1428_ & ~_0694_;
	assign _0696_ = _0617_ | _0530_;
	assign _0697_ = _0696_ | _0533_;
	assign _0698_ = ~(_0696_ | _0533_);
	assign _0699_ = _0698_ & ~_0370_;
	assign _0700_ = _0699_ | _0697_;
	assign _0701_ = _0608_ | _0517_;
	assign _0702_ = _0701_ | _0527_;
	assign _0703_ = _0702_ | _0365_;
	assign _0704_ = ~(_0701_ | _0526_);
	assign _0705_ = _0615_ & ~_0608_;
	assign _0706_ = \mchip.my_core.regA.Q [7] & ~\mchip.my_core.regB.Q [7];
	assign _0707_ = _0706_ | _0705_;
	assign _0708_ = _0707_ | _0704_;
	assign _0709_ = _0703_ & ~_0708_;
	assign _0710_ = _0709_ ^ _0700_;
	assign _0711_ = _1433_ & ~_0710_;
	assign _0712_ = _0711_ | _0695_;
	assign _0713_ = (_1396_ ? _1423_ : _1416_);
	assign _0714_ = _0709_ & ~_0713_;
	assign _0715_ = _0714_ | _0712_;
	assign _0716_ = _1424_ | _1421_;
	assign _0717_ = _0716_ | _1414_;
	assign _0718_ = _0713_ & ~_0717_;
	assign _0719_ = _1433_ | _1428_;
	assign _0720_ = _0718_ & ~_0719_;
	assign _0721_ = (_0720_ ? _0690_ : _0715_);
	assign \mchip.my_core.Unit.flag_reg.d [0] = (_1028_ ? _0681_ : _0721_);
	assign _0722_ = ~(_0126_ | _1443_);
	assign _0723_ = _0286_ | _0205_;
	assign _0724_ = _0722_ & ~_0723_;
	assign _0725_ = _0633_ | _0549_;
	assign _0726_ = ~_0378_;
	assign _0727_ = _0457_ | ~_0726_;
	assign _0728_ = _0727_ | _0725_;
	assign _0729_ = _0724_ & ~_0728_;
	assign _0730_ = _1417_ | _1388_;
	assign _0731_ = ~(_0730_ | _1028_);
	assign _0732_ = _0117_ | _1417_;
	assign _0733_ = ~(_0732_ | _1028_);
	assign _0734_ = ~(_0733_ | _0731_);
	assign _0735_ = _0276_ | _1417_;
	assign _0736_ = ~(_0735_ | _1028_);
	assign _0737_ = _0187_ | _1417_;
	assign _0738_ = ~(_0737_ | _1028_);
	assign _0739_ = _0738_ | _0736_;
	assign _0740_ = _0734_ & ~_0739_;
	assign _0741_ = _1417_ | ~_0617_;
	assign _0742_ = ~(_0741_ | _1028_);
	assign _0743_ = _0531_ | _1417_;
	assign _0744_ = ~(_0743_ | _1028_);
	assign _0745_ = _0744_ | _0742_;
	assign _0746_ = _0448_ | _1417_;
	assign _0747_ = ~(_0746_ | _1028_);
	assign _0748_ = _0367_ | _1417_;
	assign _0749_ = ~(_0748_ | _1028_);
	assign _0750_ = _0749_ | _0747_;
	assign _0751_ = _0750_ | _0745_;
	assign _0752_ = _0740_ & ~_0751_;
	assign _0753_ = (_1417_ ? _0729_ : _0752_);
	assign \mchip.my_core.Unit.flag_reg.d [1] = (_1028_ ? _0729_ : _0753_);
	assign _0754_ = (_1417_ ? _0633_ : _0742_);
	assign \mchip.my_core.Unit.flag_reg.d [2] = (_1028_ ? _0633_ : _0754_);
	assign _0755_ = ~(_0633_ ^ _0549_);
	assign _0756_ = _0457_ ^ _0726_;
	assign _0757_ = _0756_ ^ _0755_;
	assign _0758_ = ~(_0286_ ^ _0205_);
	assign _0759_ = _0126_ ^ _1443_;
	assign _0760_ = _0759_ ^ _0758_;
	assign _0761_ = _0760_ ^ _0757_;
	assign _0762_ = ~(_0744_ ^ _0742_);
	assign _0763_ = ~(_0749_ ^ _0747_);
	assign _0764_ = _0763_ ^ _0762_;
	assign _0765_ = ~(_0738_ ^ _0736_);
	assign _0766_ = _0733_ ^ _0731_;
	assign _0767_ = _0766_ ^ _0765_;
	assign _0768_ = _0767_ ^ _0764_;
	assign _0769_ = (_1417_ ? _0761_ : _0768_);
	assign \mchip.my_core.Unit.flag_reg.d [3] = (_1028_ ? _0761_ : _0769_);
	assign _0037_ = \mchip.my_core.Stack.bus [0] & _1158_;
	assign _0038_ = \mchip.my_core.Stack.bus [1] & _1158_;
	assign _0039_ = \mchip.my_core.Stack.bus [2] & _1158_;
	assign _0040_ = \mchip.my_core.Stack.bus [3] & _1158_;
	assign _0041_ = \mchip.my_core.Stack.bus [4] & _1158_;
	assign _0042_ = \mchip.my_core.Stack.bus [5] & _1158_;
	assign _0043_ = \mchip.my_core.Stack.bus [6] & _1158_;
	assign _0044_ = \mchip.my_core.Stack.bus [7] & _1158_;
	assign _0770_ = ~(_1071_ & _0900_);
	assign _0771_ = _0770_ & ~_1463_;
	assign _0772_ = (\mchip.my_core.Brain.state [2] ? _0890_ : _0896_);
	assign _0773_ = _0772_ | _0900_;
	assign _0774_ = _0773_ | ~_0892_;
	assign _0775_ = ~_0947_;
	assign _0776_ = (\mchip.my_core.IR.Q [7] ? _0957_ : _0775_);
	assign _0777_ = _0989_ | _0986_;
	assign _0778_ = _0776_ & ~_0777_;
	assign _0779_ = _0927_ | ~_1051_;
	assign _0780_ = _0778_ & ~_0779_;
	assign _0781_ = _0564_ | ~_0919_;
	assign _0782_ = _0781_ | _1176_;
	assign _0783_ = _0780_ & ~_0782_;
	assign _0784_ = (_0774_ ? _0771_ : _0783_);
	assign _0785_ = \mchip.my_core.Brain.cycle [2] & ~_0784_;
	assign _0786_ = _0919_ | _0892_;
	assign _0787_ = _1170_ | _1023_;
	assign _0788_ = _0892_ & ~_0787_;
	assign _0789_ = (_0788_ ? _0929_ : _0786_);
	assign _0790_ = \mchip.my_core.Brain.cycle [1] & ~_0789_;
	assign _0791_ = ~(_0790_ | _0785_);
	assign _0792_ = _0791_ & ~_1344_;
	assign \mchip.my_core.Sync  = _1067_ & ~_0792_;
	assign _0793_ = (_0900_ ? _1091_ : _1263_);
	assign _0794_ = _0793_ | _1064_;
	assign _0795_ = _0794_ & ~_1451_;
	assign \mchip.my_core.regB.en  = ~(_0795_ | _1027_);
	assign _0796_ = _0896_ | _0890_;
	assign _0797_ = _0796_ | _0889_;
	assign _0798_ = (_0900_ ? _1022_ : _0797_);
	assign _0799_ = \mchip.my_core.Brain.cycle [0] & ~_0798_;
	assign _0800_ = _1445_ & ~_0799_;
	assign \mchip.my_core.A_en  = ~(_0800_ | _1201_);
	assign _0801_ = _0896_ & \mchip.my_core.Ready ;
	assign _0802_ = _1176_ | ~_0919_;
	assign _0803_ = (_0876_ ? _0886_ : _0909_);
	assign _0804_ = _0802_ & ~_0803_;
	assign _0805_ = ~(_0804_ | _0892_);
	assign _0806_ = _0805_ | _0801_;
	assign _0807_ = _1262_ & ~_0806_;
	assign _0808_ = _0807_ | _0897_;
	assign _0809_ = _0808_ | _1124_;
	assign _0810_ = _0990_ | _0926_;
	assign _0811_ = _0810_ | _0975_;
	assign _0812_ = _0811_ | _1448_;
	assign _0813_ = _0812_ | _0564_;
	assign _0814_ = ~(_0813_ | _0892_);
	assign _0815_ = _0814_ | _0801_;
	assign _0816_ = ~(_0815_ | _0900_);
	assign _0817_ = _0816_ | _0897_;
	assign _0818_ = \mchip.my_core.Brain.cycle [2] & ~_0817_;
	assign _0819_ = _0809_ & ~_0818_;
	assign _0820_ = _1300_ | _0994_;
	assign _0821_ = _0820_ | _0969_;
	assign _0822_ = _0954_ | \mchip.my_core.Intr ;
	assign _0823_ = _0969_ & ~_0822_;
	assign _0824_ = _0876_ ^ _1127_;
	assign _0825_ = _1300_ & ~_0824_;
	assign _0826_ = _0825_ | _0823_;
	assign _0827_ = _0821_ & ~_0826_;
	assign _0828_ = ~(_0827_ | _0892_);
	assign _0829_ = ~(_0828_ | _0801_);
	assign _0830_ = _0900_ & ~_0564_;
	assign _0831_ = _0829_ & ~_0830_;
	assign _0832_ = _0831_ | _0897_;
	assign _0833_ = \mchip.my_core.Brain.cycle [0] & ~_0832_;
	assign _0834_ = _0819_ & ~_0833_;
	assign \mchip.my_core.Brain.next_state [0] = _1067_ & ~_0834_;
	assign _0835_ = _0564_ & ~_1262_;
	assign _0836_ = _0835_ | _1023_;
	assign _0837_ = _0892_ & ~_0836_;
	assign _0838_ = _0837_ | _0897_;
	assign _0839_ = \mchip.my_core.Brain.cycle [0] & ~_0838_;
	assign _0840_ = _1024_ & _0892_;
	assign _0841_ = _0840_ | _0897_;
	assign _0842_ = \mchip.my_core.Brain.cycle [2] & ~_0841_;
	assign _0843_ = \mchip.my_core.Brain.cycle [1] & ~_0841_;
	assign _0844_ = _0843_ | _0842_;
	assign _0845_ = _0844_ | _0839_;
	assign \mchip.my_core.Brain.next_state [1] = _0845_ | _1066_;
	assign _0846_ = _0805_ | _0900_;
	assign _0847_ = ~(_0846_ | _0897_);
	assign _0848_ = _0847_ | _1124_;
	assign _0849_ = _0814_ | _0900_;
	assign _0850_ = ~(_0849_ | _0897_);
	assign _0851_ = \mchip.my_core.Brain.cycle [2] & ~_0850_;
	assign _0852_ = _0848_ & ~_0851_;
	assign _0853_ = _0954_ | ~\mchip.my_core.Intr ;
	assign _0854_ = _0969_ & ~_0853_;
	assign _0855_ = _0854_ | _0825_;
	assign _0856_ = _0821_ & ~_0855_;
	assign _0857_ = ~(_0856_ | _0892_);
	assign _0858_ = _0857_ | _0830_;
	assign _0859_ = ~(_0858_ | _0897_);
	assign _0860_ = \mchip.my_core.Brain.cycle [0] & ~_0859_;
	assign _0861_ = _0852_ & ~_0860_;
	assign \mchip.my_core.Brain.next_state [2] = _1067_ & ~_0861_;
	assign _0862_ = _1160_ | ~_1161_;
	assign _0863_ = _0862_ | _1159_;
	assign _0061_ = _1157_ & ~_0863_;
	assign _0864_ = _0862_ | _1164_;
	assign _0060_ = _1157_ & ~_0864_;
	assign _0865_ = _1313_ | _1159_;
	assign _0059_ = _1157_ & ~_0865_;
	assign _0045_ = \mchip.my_core.S_Intr  | \mchip.my_core.Intr ;
	assign \mchip.my_core.A_rst  = _1247_ | io_in[13];
	assign _1498_[0] = ~\mchip.my_core.SP_SEL.Q [0];
	assign _0866_ = ~\mchip.my_core.Unit.flag_reg.Q [0];
	assign _0867_ = \mchip.my_core.IR.Q [4] & ~\mchip.my_core.IR.Q [3];
	assign _0868_ = _0867_ & ~\mchip.my_core.Unit.flag_reg.Q [2];
	assign _0869_ = ~(\mchip.my_core.IR.Q [4] & \mchip.my_core.IR.Q [3]);
	assign _0870_ = ~(_0869_ | \mchip.my_core.Unit.flag_reg.Q [3]);
	assign _0871_ = _0870_ | _0868_;
	assign _0872_ = \mchip.my_core.IR.Q [3] & ~\mchip.my_core.IR.Q [4];
	assign _0873_ = _0872_ & ~\mchip.my_core.Unit.flag_reg.Q [1];
	assign _0874_ = _0873_ | _0871_;
	assign _0875_ = ~(\mchip.my_core.IR.Q [4] | \mchip.my_core.IR.Q [3]);
	assign _0876_ = (_0875_ ? _0866_ : _0874_);
	assign _0877_ = \mchip.my_core.IR.Q [5] | \mchip.my_core.IR.Q [2];
	assign _0878_ = \mchip.my_core.IR.Q [0] | ~\mchip.my_core.IR.Q [1];
	assign _0879_ = ~(_0878_ | _0877_);
	assign _0880_ = \mchip.my_core.IR.Q [6] & ~\mchip.my_core.IR.Q [7];
	assign _0881_ = ~_0880_;
	assign _0882_ = _0879_ & ~_0881_;
	assign _0883_ = \mchip.my_core.IR.Q [1] | \mchip.my_core.IR.Q [0];
	assign _0884_ = _0883_ | _0877_;
	assign _0885_ = ~(_0884_ | _0881_);
	assign _0886_ = _0885_ | _0882_;
	assign _0887_ = ~(_0886_ & _0876_);
	assign _0888_ = \mchip.my_core.Brain.state [0] & \mchip.my_core.Brain.state [1];
	assign _0889_ = _0888_ & ~\mchip.my_core.Brain.state [2];
	assign _0890_ = \mchip.my_core.Brain.state [0] & ~\mchip.my_core.Brain.state [1];
	assign _0891_ = _0890_ & ~\mchip.my_core.Brain.state [2];
	assign _0892_ = ~(_0891_ | _0889_);
	assign _0893_ = _0892_ | io_in[13];
	assign _0894_ = _0893_ | _0887_;
	assign _0895_ = \mchip.my_core.Brain.cycle [1] & ~_0894_;
	assign _0896_ = ~(\mchip.my_core.Brain.state [0] | \mchip.my_core.Brain.state [1]);
	assign _0897_ = \mchip.my_core.Brain.state [1] & ~\mchip.my_core.Brain.state [0];
	assign _0898_ = ~(_0897_ | _0896_);
	assign _0899_ = ~\mchip.my_core.Brain.state [2];
	assign _0900_ = _0888_ & ~_0899_;
	assign _0901_ = _0898_ & ~_0900_;
	assign _0902_ = _0901_ | io_in[13];
	assign _0903_ = \mchip.my_core.Brain.cycle [1] & ~_0902_;
	assign _0904_ = \mchip.my_core.IR.Q [2] | ~\mchip.my_core.IR.Q [5];
	assign _0905_ = _0904_ | _0878_;
	assign _0906_ = ~(_0905_ | _0881_);
	assign _0907_ = _0904_ | _0883_;
	assign _0908_ = _0880_ & ~_0907_;
	assign _0909_ = _0908_ | _0906_;
	assign _0910_ = _0876_ | ~_0909_;
	assign _0911_ = _0910_ | _0893_;
	assign _0912_ = \mchip.my_core.Brain.cycle [1] & ~_0911_;
	assign _0913_ = _0912_ | _0903_;
	assign _0914_ = \mchip.my_core.IR.Q [6] | \mchip.my_core.IR.Q [7];
	assign _0915_ = ~(\mchip.my_core.IR.Q [4] & \mchip.my_core.IR.Q [5]);
	assign _0916_ = _0915_ | _0914_;
	assign _0917_ = \mchip.my_core.IR.Q [3] & \mchip.my_core.IR.Q [2];
	assign _0918_ = _0878_ | ~_0917_;
	assign _0919_ = _0918_ | _0916_;
	assign _0920_ = _0919_ & ~_0909_;
	assign _0921_ = ~\mchip.my_core.IR.Q [7];
	assign _0922_ = ~(\mchip.my_core.IR.Q [6] & \mchip.my_core.IR.Q [2]);
	assign _0923_ = _0922_ | _0878_;
	assign _0924_ = _0921_ & ~_0923_;
	assign _0925_ = _0922_ | _0883_;
	assign _0926_ = _0921_ & ~_0925_;
	assign _0927_ = _0926_ | _0924_;
	assign _0928_ = _0927_ | _0886_;
	assign _0929_ = _0920_ & ~_0928_;
	assign _0930_ = _0929_ | _0893_;
	assign _0931_ = \mchip.my_core.Brain.cycle [2] & ~_0930_;
	assign _0932_ = _0892_ | _0886_;
	assign _0933_ = ~io_in[13];
	assign _0934_ = ~(_0919_ & _0933_);
	assign _0935_ = _0934_ | _0932_;
	assign _0936_ = _0935_ | _0909_;
	assign _0937_ = \mchip.my_core.Brain.cycle [1] & ~_0936_;
	assign _0938_ = _0937_ | _0931_;
	assign _0939_ = _0938_ | _0913_;
	assign _0002_ = _0939_ | _0895_;
	assign _0940_ = \mchip.my_core.Brain.cycle [2] & ~_0902_;
	assign _0941_ = ~(_0900_ & _0933_);
	assign _0942_ = ~(\mchip.my_core.IR.Q [6] & \mchip.my_core.IR.Q [5]);
	assign _0943_ = ~(_0942_ | _0869_);
	assign _0564_ = _0943_ & ~_0921_;
	assign _0944_ = _0941_ | ~_0564_;
	assign _0945_ = \mchip.my_core.Brain.cycle [0] & ~_0944_;
	assign _0946_ = _0892_ | ~_0929_;
	assign _0947_ = \mchip.my_core.IR.Q [6] & \mchip.my_core.IR.Q [0];
	assign _0948_ = (\mchip.my_core.IR.Q [7] ? _0943_ : _0947_);
	assign _0949_ = _0948_ | io_in[13];
	assign _0950_ = _0949_ | _0946_;
	assign _0951_ = \mchip.my_core.Brain.cycle [2] & ~_0950_;
	assign _0952_ = _0951_ | _0945_;
	assign _0953_ = \mchip.my_core.IR.Q [5] & ~_0869_;
	assign _0954_ = \mchip.my_core.IR.Q [7] & ~_0953_;
	assign _0955_ = _0892_ | ~_0954_;
	assign _0956_ = ~(\mchip.my_core.IR.Q [1] & \mchip.my_core.IR.Q [0]);
	assign _0957_ = _0956_ | _0922_;
	assign _0958_ = \mchip.my_core.IR.Q [7] & ~_0957_;
	assign _0959_ = _0917_ & ~_0956_;
	assign _0960_ = \mchip.my_core.IR.Q [6] & \mchip.my_core.IR.Q [7];
	assign _0961_ = _0915_ | ~_0960_;
	assign _0962_ = _0959_ & ~_0961_;
	assign _0963_ = \mchip.my_core.IR.Q [2] | \mchip.my_core.IR.Q [1];
	assign _0964_ = _0875_ & ~_0963_;
	assign _0965_ = \mchip.my_core.IR.Q [6] | \mchip.my_core.IR.Q [5];
	assign _0966_ = _0965_ | \mchip.my_core.IR.Q [7];
	assign _0967_ = _0964_ & ~_0966_;
	assign _0968_ = _0967_ | _0962_;
	assign _0969_ = _0968_ | _0958_;
	assign _0970_ = ~(_0969_ & _0933_);
	assign _0971_ = _0970_ | _0955_;
	assign _0972_ = \mchip.my_core.Brain.cycle [0] & ~_0971_;
	assign _0973_ = _0908_ | _0882_;
	assign _0974_ = _0973_ | _0906_;
	assign _0975_ = _0924_ | _0885_;
	assign _0976_ = \mchip.my_core.IR.Q [6] | ~\mchip.my_core.IR.Q [2];
	assign _0977_ = _0976_ | _0883_;
	assign _0978_ = _0921_ & ~_0977_;
	assign _0979_ = _0978_ | _0926_;
	assign _0980_ = _0979_ | _0975_;
	assign _0981_ = _0976_ | _0956_;
	assign _0982_ = \mchip.my_core.IR.Q [7] & ~_0981_;
	always @(posedge io_in[12])
		if (_0013_)
			if (!_0049_)
				\mchip.my_core.Stack.rf[3] [0] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[3] [0] <= _0023_;
	always @(posedge io_in[12])
		if (_0013_)
			if (!_0049_)
				\mchip.my_core.Stack.rf[3] [1] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[3] [1] <= _0028_;
	always @(posedge io_in[12])
		if (_0013_)
			if (!_0049_)
				\mchip.my_core.Stack.rf[3] [2] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[3] [2] <= _0029_;
	always @(posedge io_in[12])
		if (_0013_)
			if (!_0049_)
				\mchip.my_core.Stack.rf[3] [3] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[3] [3] <= _0030_;
	always @(posedge io_in[12])
		if (_0013_)
			if (!_0049_)
				\mchip.my_core.Stack.rf[3] [4] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[3] [4] <= _0031_;
	always @(posedge io_in[12])
		if (_0013_)
			if (!_0049_)
				\mchip.my_core.Stack.rf[3] [5] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[3] [5] <= _0032_;
	always @(posedge io_in[12])
		if (_0013_)
			if (!_0049_)
				\mchip.my_core.Stack.rf[3] [6] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[3] [6] <= _0033_;
	always @(posedge io_in[12])
		if (_0013_)
			if (!_0049_)
				\mchip.my_core.Stack.rf[3] [7] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[3] [7] <= _0034_;
	always @(posedge io_in[12])
		if (_0013_)
			if (!_0049_)
				\mchip.my_core.Stack.rf[3] [8] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[3] [8] <= _0035_;
	always @(posedge io_in[12])
		if (_0013_)
			if (!_0049_)
				\mchip.my_core.Stack.rf[3] [9] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[3] [9] <= _0036_;
	always @(posedge io_in[12])
		if (_0013_)
			if (!_0049_)
				\mchip.my_core.Stack.rf[3] [10] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[3] [10] <= _0024_;
	always @(posedge io_in[12])
		if (_0013_)
			if (!_0049_)
				\mchip.my_core.Stack.rf[3] [11] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[3] [11] <= _0025_;
	always @(posedge io_in[12])
		if (_0013_)
			if (!_0049_)
				\mchip.my_core.Stack.rf[3] [12] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[3] [12] <= _0026_;
	always @(posedge io_in[12])
		if (_0013_)
			if (!_0049_)
				\mchip.my_core.Stack.rf[3] [13] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[3] [13] <= _0027_;
	always @(posedge io_in[12])
		if (_0009_)
			if (!_0053_)
				\mchip.my_core.Stack.rf[7] [0] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[7] [0] <= _0023_;
	always @(posedge io_in[12])
		if (_0009_)
			if (!_0053_)
				\mchip.my_core.Stack.rf[7] [1] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[7] [1] <= _0028_;
	always @(posedge io_in[12])
		if (_0009_)
			if (!_0053_)
				\mchip.my_core.Stack.rf[7] [2] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[7] [2] <= _0029_;
	always @(posedge io_in[12])
		if (_0009_)
			if (!_0053_)
				\mchip.my_core.Stack.rf[7] [3] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[7] [3] <= _0030_;
	always @(posedge io_in[12])
		if (_0009_)
			if (!_0053_)
				\mchip.my_core.Stack.rf[7] [4] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[7] [4] <= _0031_;
	always @(posedge io_in[12])
		if (_0009_)
			if (!_0053_)
				\mchip.my_core.Stack.rf[7] [5] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[7] [5] <= _0032_;
	always @(posedge io_in[12])
		if (_0009_)
			if (!_0053_)
				\mchip.my_core.Stack.rf[7] [6] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[7] [6] <= _0033_;
	always @(posedge io_in[12])
		if (_0009_)
			if (!_0053_)
				\mchip.my_core.Stack.rf[7] [7] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[7] [7] <= _0034_;
	always @(posedge io_in[12])
		if (_0009_)
			if (!_0053_)
				\mchip.my_core.Stack.rf[7] [8] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[7] [8] <= _0035_;
	always @(posedge io_in[12])
		if (_0009_)
			if (!_0053_)
				\mchip.my_core.Stack.rf[7] [9] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[7] [9] <= _0036_;
	always @(posedge io_in[12])
		if (_0009_)
			if (!_0053_)
				\mchip.my_core.Stack.rf[7] [10] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[7] [10] <= _0024_;
	always @(posedge io_in[12])
		if (_0009_)
			if (!_0053_)
				\mchip.my_core.Stack.rf[7] [11] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[7] [11] <= _0025_;
	always @(posedge io_in[12])
		if (_0009_)
			if (!_0053_)
				\mchip.my_core.Stack.rf[7] [12] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[7] [12] <= _0026_;
	always @(posedge io_in[12])
		if (_0009_)
			if (!_0053_)
				\mchip.my_core.Stack.rf[7] [13] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[7] [13] <= _0027_;
	always @(posedge io_in[12])
		if (_0059_)
			\mchip.my_core.rf.rf[5] [0] <= _0037_;
	always @(posedge io_in[12])
		if (_0059_)
			\mchip.my_core.rf.rf[5] [1] <= _0038_;
	always @(posedge io_in[12])
		if (_0059_)
			\mchip.my_core.rf.rf[5] [2] <= _0039_;
	always @(posedge io_in[12])
		if (_0059_)
			\mchip.my_core.rf.rf[5] [3] <= _0040_;
	always @(posedge io_in[12])
		if (_0059_)
			\mchip.my_core.rf.rf[5] [4] <= _0041_;
	always @(posedge io_in[12])
		if (_0059_)
			\mchip.my_core.rf.rf[5] [5] <= _0042_;
	always @(posedge io_in[12])
		if (_0059_)
			\mchip.my_core.rf.rf[5] [6] <= _0043_;
	always @(posedge io_in[12])
		if (_0059_)
			\mchip.my_core.rf.rf[5] [7] <= _0044_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.my_core.rf.rf[6] [0] <= 1'h0;
		else if (_0060_)
			\mchip.my_core.rf.rf[6] [0] <= _0037_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.my_core.rf.rf[6] [1] <= 1'h0;
		else if (_0060_)
			\mchip.my_core.rf.rf[6] [1] <= _0038_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.my_core.rf.rf[6] [2] <= 1'h0;
		else if (_0060_)
			\mchip.my_core.rf.rf[6] [2] <= _0039_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.my_core.rf.rf[6] [3] <= 1'h0;
		else if (_0060_)
			\mchip.my_core.rf.rf[6] [3] <= _0040_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.my_core.rf.rf[6] [4] <= 1'h0;
		else if (_0060_)
			\mchip.my_core.rf.rf[6] [4] <= _0041_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.my_core.rf.rf[6] [5] <= 1'h0;
		else if (_0060_)
			\mchip.my_core.rf.rf[6] [5] <= _0042_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.my_core.rf.rf[6] [6] <= 1'h0;
		else if (_0060_)
			\mchip.my_core.rf.rf[6] [6] <= _0043_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.my_core.rf.rf[6] [7] <= 1'h0;
		else if (_0060_)
			\mchip.my_core.rf.rf[6] [7] <= _0044_;
	always @(posedge io_in[12])
		if (_0004_)
			if (!_0058_)
				\mchip.my_core.rf.rf[4] [0] <= 1'h0;
			else
				\mchip.my_core.rf.rf[4] [0] <= _0037_;
	always @(posedge io_in[12])
		if (_0004_)
			if (!_0058_)
				\mchip.my_core.rf.rf[4] [1] <= 1'h0;
			else
				\mchip.my_core.rf.rf[4] [1] <= _0038_;
	always @(posedge io_in[12])
		if (_0004_)
			if (!_0058_)
				\mchip.my_core.rf.rf[4] [2] <= 1'h0;
			else
				\mchip.my_core.rf.rf[4] [2] <= _0039_;
	always @(posedge io_in[12])
		if (_0004_)
			if (!_0058_)
				\mchip.my_core.rf.rf[4] [3] <= 1'h0;
			else
				\mchip.my_core.rf.rf[4] [3] <= _0040_;
	always @(posedge io_in[12])
		if (_0004_)
			if (!_0058_)
				\mchip.my_core.rf.rf[4] [4] <= 1'h0;
			else
				\mchip.my_core.rf.rf[4] [4] <= _0041_;
	always @(posedge io_in[12])
		if (_0004_)
			if (!_0058_)
				\mchip.my_core.rf.rf[4] [5] <= 1'h0;
			else
				\mchip.my_core.rf.rf[4] [5] <= _0042_;
	always @(posedge io_in[12])
		if (_0004_)
			if (!_0058_)
				\mchip.my_core.rf.rf[4] [6] <= 1'h0;
			else
				\mchip.my_core.rf.rf[4] [6] <= _0043_;
	always @(posedge io_in[12])
		if (_0004_)
			if (!_0058_)
				\mchip.my_core.rf.rf[4] [7] <= 1'h0;
			else
				\mchip.my_core.rf.rf[4] [7] <= _0044_;
	always @(posedge io_in[12])
		if (_0005_)
			if (!_0057_)
				\mchip.my_core.rf.rf[3] [0] <= 1'h0;
			else
				\mchip.my_core.rf.rf[3] [0] <= _0037_;
	always @(posedge io_in[12])
		if (_0005_)
			if (!_0057_)
				\mchip.my_core.rf.rf[3] [1] <= 1'h0;
			else
				\mchip.my_core.rf.rf[3] [1] <= _0038_;
	always @(posedge io_in[12])
		if (_0005_)
			if (!_0057_)
				\mchip.my_core.rf.rf[3] [2] <= 1'h0;
			else
				\mchip.my_core.rf.rf[3] [2] <= _0039_;
	always @(posedge io_in[12])
		if (_0005_)
			if (!_0057_)
				\mchip.my_core.rf.rf[3] [3] <= 1'h0;
			else
				\mchip.my_core.rf.rf[3] [3] <= _0040_;
	always @(posedge io_in[12])
		if (_0005_)
			if (!_0057_)
				\mchip.my_core.rf.rf[3] [4] <= 1'h0;
			else
				\mchip.my_core.rf.rf[3] [4] <= _0041_;
	always @(posedge io_in[12])
		if (_0005_)
			if (!_0057_)
				\mchip.my_core.rf.rf[3] [5] <= 1'h0;
			else
				\mchip.my_core.rf.rf[3] [5] <= _0042_;
	always @(posedge io_in[12])
		if (_0005_)
			if (!_0057_)
				\mchip.my_core.rf.rf[3] [6] <= 1'h0;
			else
				\mchip.my_core.rf.rf[3] [6] <= _0043_;
	always @(posedge io_in[12])
		if (_0005_)
			if (!_0057_)
				\mchip.my_core.rf.rf[3] [7] <= 1'h0;
			else
				\mchip.my_core.rf.rf[3] [7] <= _0044_;
	always @(posedge io_in[12])
		if (_0006_)
			if (!_0056_)
				\mchip.my_core.rf.rf[2] [0] <= 1'h0;
			else
				\mchip.my_core.rf.rf[2] [0] <= _0037_;
	always @(posedge io_in[12])
		if (_0006_)
			if (!_0056_)
				\mchip.my_core.rf.rf[2] [1] <= 1'h0;
			else
				\mchip.my_core.rf.rf[2] [1] <= _0038_;
	always @(posedge io_in[12])
		if (_0006_)
			if (!_0056_)
				\mchip.my_core.rf.rf[2] [2] <= 1'h0;
			else
				\mchip.my_core.rf.rf[2] [2] <= _0039_;
	always @(posedge io_in[12])
		if (_0006_)
			if (!_0056_)
				\mchip.my_core.rf.rf[2] [3] <= 1'h0;
			else
				\mchip.my_core.rf.rf[2] [3] <= _0040_;
	always @(posedge io_in[12])
		if (_0006_)
			if (!_0056_)
				\mchip.my_core.rf.rf[2] [4] <= 1'h0;
			else
				\mchip.my_core.rf.rf[2] [4] <= _0041_;
	always @(posedge io_in[12])
		if (_0006_)
			if (!_0056_)
				\mchip.my_core.rf.rf[2] [5] <= 1'h0;
			else
				\mchip.my_core.rf.rf[2] [5] <= _0042_;
	always @(posedge io_in[12])
		if (_0006_)
			if (!_0056_)
				\mchip.my_core.rf.rf[2] [6] <= 1'h0;
			else
				\mchip.my_core.rf.rf[2] [6] <= _0043_;
	always @(posedge io_in[12])
		if (_0006_)
			if (!_0056_)
				\mchip.my_core.rf.rf[2] [7] <= 1'h0;
			else
				\mchip.my_core.rf.rf[2] [7] <= _0044_;
	always @(posedge io_in[12])
		if (_0007_)
			if (!_0055_)
				\mchip.my_core.rf.rf[1] [0] <= 1'h0;
			else
				\mchip.my_core.rf.rf[1] [0] <= _0037_;
	always @(posedge io_in[12])
		if (_0007_)
			if (!_0055_)
				\mchip.my_core.rf.rf[1] [1] <= 1'h0;
			else
				\mchip.my_core.rf.rf[1] [1] <= _0038_;
	always @(posedge io_in[12])
		if (_0007_)
			if (!_0055_)
				\mchip.my_core.rf.rf[1] [2] <= 1'h0;
			else
				\mchip.my_core.rf.rf[1] [2] <= _0039_;
	always @(posedge io_in[12])
		if (_0007_)
			if (!_0055_)
				\mchip.my_core.rf.rf[1] [3] <= 1'h0;
			else
				\mchip.my_core.rf.rf[1] [3] <= _0040_;
	always @(posedge io_in[12])
		if (_0007_)
			if (!_0055_)
				\mchip.my_core.rf.rf[1] [4] <= 1'h0;
			else
				\mchip.my_core.rf.rf[1] [4] <= _0041_;
	always @(posedge io_in[12])
		if (_0007_)
			if (!_0055_)
				\mchip.my_core.rf.rf[1] [5] <= 1'h0;
			else
				\mchip.my_core.rf.rf[1] [5] <= _0042_;
	always @(posedge io_in[12])
		if (_0007_)
			if (!_0055_)
				\mchip.my_core.rf.rf[1] [6] <= 1'h0;
			else
				\mchip.my_core.rf.rf[1] [6] <= _0043_;
	always @(posedge io_in[12])
		if (_0007_)
			if (!_0055_)
				\mchip.my_core.rf.rf[1] [7] <= 1'h0;
			else
				\mchip.my_core.rf.rf[1] [7] <= _0044_;
	always @(posedge io_in[12])
		if (_0008_)
			if (!_0054_)
				\mchip.my_core.rf.rf[0] [0] <= 1'h0;
			else
				\mchip.my_core.rf.rf[0] [0] <= _0037_;
	always @(posedge io_in[12])
		if (_0008_)
			if (!_0054_)
				\mchip.my_core.rf.rf[0] [1] <= 1'h0;
			else
				\mchip.my_core.rf.rf[0] [1] <= _0038_;
	always @(posedge io_in[12])
		if (_0008_)
			if (!_0054_)
				\mchip.my_core.rf.rf[0] [2] <= 1'h0;
			else
				\mchip.my_core.rf.rf[0] [2] <= _0039_;
	always @(posedge io_in[12])
		if (_0008_)
			if (!_0054_)
				\mchip.my_core.rf.rf[0] [3] <= 1'h0;
			else
				\mchip.my_core.rf.rf[0] [3] <= _0040_;
	always @(posedge io_in[12])
		if (_0008_)
			if (!_0054_)
				\mchip.my_core.rf.rf[0] [4] <= 1'h0;
			else
				\mchip.my_core.rf.rf[0] [4] <= _0041_;
	always @(posedge io_in[12])
		if (_0008_)
			if (!_0054_)
				\mchip.my_core.rf.rf[0] [5] <= 1'h0;
			else
				\mchip.my_core.rf.rf[0] [5] <= _0042_;
	always @(posedge io_in[12])
		if (_0008_)
			if (!_0054_)
				\mchip.my_core.rf.rf[0] [6] <= 1'h0;
			else
				\mchip.my_core.rf.rf[0] [6] <= _0043_;
	always @(posedge io_in[12])
		if (_0008_)
			if (!_0054_)
				\mchip.my_core.rf.rf[0] [7] <= 1'h0;
			else
				\mchip.my_core.rf.rf[0] [7] <= _0044_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0000_[0] <= 1'h0;
		else
			_0000_[0] <= _0020_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0000_[1] <= 1'h0;
		else
			_0000_[1] <= _0021_;
	always @(posedge io_in[12])
		if (io_in[13])
			_0000_[2] <= 1'h0;
		else
			_0000_[2] <= _0022_;
	always @(posedge io_in[12])
		if (_0010_)
			if (!_0052_)
				\mchip.my_core.Stack.rf[6] [0] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[6] [0] <= _0023_;
	always @(posedge io_in[12])
		if (_0010_)
			if (!_0052_)
				\mchip.my_core.Stack.rf[6] [1] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[6] [1] <= _0028_;
	always @(posedge io_in[12])
		if (_0010_)
			if (!_0052_)
				\mchip.my_core.Stack.rf[6] [2] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[6] [2] <= _0029_;
	always @(posedge io_in[12])
		if (_0010_)
			if (!_0052_)
				\mchip.my_core.Stack.rf[6] [3] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[6] [3] <= _0030_;
	always @(posedge io_in[12])
		if (_0010_)
			if (!_0052_)
				\mchip.my_core.Stack.rf[6] [4] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[6] [4] <= _0031_;
	always @(posedge io_in[12])
		if (_0010_)
			if (!_0052_)
				\mchip.my_core.Stack.rf[6] [5] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[6] [5] <= _0032_;
	always @(posedge io_in[12])
		if (_0010_)
			if (!_0052_)
				\mchip.my_core.Stack.rf[6] [6] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[6] [6] <= _0033_;
	always @(posedge io_in[12])
		if (_0010_)
			if (!_0052_)
				\mchip.my_core.Stack.rf[6] [7] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[6] [7] <= _0034_;
	always @(posedge io_in[12])
		if (_0010_)
			if (!_0052_)
				\mchip.my_core.Stack.rf[6] [8] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[6] [8] <= _0035_;
	always @(posedge io_in[12])
		if (_0010_)
			if (!_0052_)
				\mchip.my_core.Stack.rf[6] [9] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[6] [9] <= _0036_;
	always @(posedge io_in[12])
		if (_0010_)
			if (!_0052_)
				\mchip.my_core.Stack.rf[6] [10] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[6] [10] <= _0024_;
	always @(posedge io_in[12])
		if (_0010_)
			if (!_0052_)
				\mchip.my_core.Stack.rf[6] [11] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[6] [11] <= _0025_;
	always @(posedge io_in[12])
		if (_0010_)
			if (!_0052_)
				\mchip.my_core.Stack.rf[6] [12] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[6] [12] <= _0026_;
	always @(posedge io_in[12])
		if (_0010_)
			if (!_0052_)
				\mchip.my_core.Stack.rf[6] [13] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[6] [13] <= _0027_;
	always @(posedge io_in[12])
		if (_0011_)
			if (!_0051_)
				\mchip.my_core.Stack.rf[5] [0] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[5] [0] <= _0023_;
	always @(posedge io_in[12])
		if (_0011_)
			if (!_0051_)
				\mchip.my_core.Stack.rf[5] [1] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[5] [1] <= _0028_;
	always @(posedge io_in[12])
		if (_0011_)
			if (!_0051_)
				\mchip.my_core.Stack.rf[5] [2] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[5] [2] <= _0029_;
	always @(posedge io_in[12])
		if (_0011_)
			if (!_0051_)
				\mchip.my_core.Stack.rf[5] [3] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[5] [3] <= _0030_;
	always @(posedge io_in[12])
		if (_0011_)
			if (!_0051_)
				\mchip.my_core.Stack.rf[5] [4] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[5] [4] <= _0031_;
	always @(posedge io_in[12])
		if (_0011_)
			if (!_0051_)
				\mchip.my_core.Stack.rf[5] [5] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[5] [5] <= _0032_;
	always @(posedge io_in[12])
		if (_0011_)
			if (!_0051_)
				\mchip.my_core.Stack.rf[5] [6] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[5] [6] <= _0033_;
	always @(posedge io_in[12])
		if (_0011_)
			if (!_0051_)
				\mchip.my_core.Stack.rf[5] [7] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[5] [7] <= _0034_;
	always @(posedge io_in[12])
		if (_0011_)
			if (!_0051_)
				\mchip.my_core.Stack.rf[5] [8] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[5] [8] <= _0035_;
	always @(posedge io_in[12])
		if (_0011_)
			if (!_0051_)
				\mchip.my_core.Stack.rf[5] [9] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[5] [9] <= _0036_;
	always @(posedge io_in[12])
		if (_0011_)
			if (!_0051_)
				\mchip.my_core.Stack.rf[5] [10] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[5] [10] <= _0024_;
	always @(posedge io_in[12])
		if (_0011_)
			if (!_0051_)
				\mchip.my_core.Stack.rf[5] [11] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[5] [11] <= _0025_;
	always @(posedge io_in[12])
		if (_0011_)
			if (!_0051_)
				\mchip.my_core.Stack.rf[5] [12] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[5] [12] <= _0026_;
	always @(posedge io_in[12])
		if (_0011_)
			if (!_0051_)
				\mchip.my_core.Stack.rf[5] [13] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[5] [13] <= _0027_;
	always @(posedge io_in[12])
		if (_0012_)
			if (!_0050_)
				\mchip.my_core.Stack.rf[4] [0] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[4] [0] <= _0023_;
	always @(posedge io_in[12])
		if (_0012_)
			if (!_0050_)
				\mchip.my_core.Stack.rf[4] [1] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[4] [1] <= _0028_;
	always @(posedge io_in[12])
		if (_0012_)
			if (!_0050_)
				\mchip.my_core.Stack.rf[4] [2] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[4] [2] <= _0029_;
	always @(posedge io_in[12])
		if (_0012_)
			if (!_0050_)
				\mchip.my_core.Stack.rf[4] [3] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[4] [3] <= _0030_;
	always @(posedge io_in[12])
		if (_0012_)
			if (!_0050_)
				\mchip.my_core.Stack.rf[4] [4] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[4] [4] <= _0031_;
	always @(posedge io_in[12])
		if (_0012_)
			if (!_0050_)
				\mchip.my_core.Stack.rf[4] [5] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[4] [5] <= _0032_;
	always @(posedge io_in[12])
		if (_0012_)
			if (!_0050_)
				\mchip.my_core.Stack.rf[4] [6] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[4] [6] <= _0033_;
	always @(posedge io_in[12])
		if (_0012_)
			if (!_0050_)
				\mchip.my_core.Stack.rf[4] [7] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[4] [7] <= _0034_;
	always @(posedge io_in[12])
		if (_0012_)
			if (!_0050_)
				\mchip.my_core.Stack.rf[4] [8] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[4] [8] <= _0035_;
	always @(posedge io_in[12])
		if (_0012_)
			if (!_0050_)
				\mchip.my_core.Stack.rf[4] [9] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[4] [9] <= _0036_;
	always @(posedge io_in[12])
		if (_0012_)
			if (!_0050_)
				\mchip.my_core.Stack.rf[4] [10] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[4] [10] <= _0024_;
	always @(posedge io_in[12])
		if (_0012_)
			if (!_0050_)
				\mchip.my_core.Stack.rf[4] [11] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[4] [11] <= _0025_;
	always @(posedge io_in[12])
		if (_0012_)
			if (!_0050_)
				\mchip.my_core.Stack.rf[4] [12] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[4] [12] <= _0026_;
	always @(posedge io_in[12])
		if (_0012_)
			if (!_0050_)
				\mchip.my_core.Stack.rf[4] [13] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[4] [13] <= _0027_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.my_core.Unit.flag_reg.Q [0] <= 1'h0;
		else if (_0018_)
			\mchip.my_core.Unit.flag_reg.Q [0] <= \mchip.my_core.Unit.flag_reg.d [0];
	always @(posedge io_in[12])
		if (_0019_)
			\mchip.my_core.Intr  <= 1'h0;
		else
			\mchip.my_core.Intr  <= _0045_;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.my_core.tempR  <= 1'h0;
		else
			\mchip.my_core.tempR  <= io_in[9];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.my_core.Ready  <= 1'h0;
		else
			\mchip.my_core.Ready  <= \mchip.my_core.tempR ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.my_core.IR.Q [0] <= 1'h0;
		else if (\mchip.my_core.IR.en )
			\mchip.my_core.IR.Q [0] <= io_in[0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.my_core.IR.Q [1] <= 1'h0;
		else if (\mchip.my_core.IR.en )
			\mchip.my_core.IR.Q [1] <= io_in[1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.my_core.IR.Q [2] <= 1'h0;
		else if (\mchip.my_core.IR.en )
			\mchip.my_core.IR.Q [2] <= io_in[2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.my_core.IR.Q [3] <= 1'h0;
		else if (\mchip.my_core.IR.en )
			\mchip.my_core.IR.Q [3] <= io_in[3];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.my_core.IR.Q [4] <= 1'h0;
		else if (\mchip.my_core.IR.en )
			\mchip.my_core.IR.Q [4] <= io_in[4];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.my_core.IR.Q [5] <= 1'h0;
		else if (\mchip.my_core.IR.en )
			\mchip.my_core.IR.Q [5] <= io_in[5];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.my_core.IR.Q [6] <= 1'h0;
		else if (\mchip.my_core.IR.en )
			\mchip.my_core.IR.Q [6] <= io_in[6];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.my_core.IR.Q [7] <= 1'h0;
		else if (\mchip.my_core.IR.en )
			\mchip.my_core.IR.Q [7] <= io_in[7];
	always @(posedge io_in[12])
		if (\mchip.my_core.A_rst )
			\mchip.my_core.regA.Q [0] <= 1'h0;
		else if (\mchip.my_core.A_en )
			\mchip.my_core.regA.Q [0] <= \mchip.my_core.regA.d [0];
	always @(posedge io_in[12])
		if (\mchip.my_core.A_rst )
			\mchip.my_core.regA.Q [1] <= 1'h0;
		else if (\mchip.my_core.A_en )
			\mchip.my_core.regA.Q [1] <= \mchip.my_core.regA.d [1];
	always @(posedge io_in[12])
		if (\mchip.my_core.A_rst )
			\mchip.my_core.regA.Q [2] <= 1'h0;
		else if (\mchip.my_core.A_en )
			\mchip.my_core.regA.Q [2] <= \mchip.my_core.regA.d [2];
	always @(posedge io_in[12])
		if (\mchip.my_core.A_rst )
			\mchip.my_core.regA.Q [3] <= 1'h0;
		else if (\mchip.my_core.A_en )
			\mchip.my_core.regA.Q [3] <= \mchip.my_core.regA.d [3];
	always @(posedge io_in[12])
		if (\mchip.my_core.A_rst )
			\mchip.my_core.regA.Q [4] <= 1'h0;
		else if (\mchip.my_core.A_en )
			\mchip.my_core.regA.Q [4] <= \mchip.my_core.regA.d [4];
	always @(posedge io_in[12])
		if (\mchip.my_core.A_rst )
			\mchip.my_core.regA.Q [5] <= 1'h0;
		else if (\mchip.my_core.A_en )
			\mchip.my_core.regA.Q [5] <= \mchip.my_core.regA.d [5];
	always @(posedge io_in[12])
		if (\mchip.my_core.A_rst )
			\mchip.my_core.regA.Q [6] <= 1'h0;
		else if (\mchip.my_core.A_en )
			\mchip.my_core.regA.Q [6] <= \mchip.my_core.regA.d [6];
	always @(posedge io_in[12])
		if (\mchip.my_core.A_rst )
			\mchip.my_core.regA.Q [7] <= 1'h0;
		else if (\mchip.my_core.A_en )
			\mchip.my_core.regA.Q [7] <= \mchip.my_core.regA.d [7];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.my_core.regB.Q [0] <= 1'h0;
		else if (\mchip.my_core.regB.en )
			\mchip.my_core.regB.Q [0] <= \mchip.my_core.Stack.bus [0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.my_core.regB.Q [1] <= 1'h0;
		else if (\mchip.my_core.regB.en )
			\mchip.my_core.regB.Q [1] <= \mchip.my_core.Stack.bus [1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.my_core.regB.Q [2] <= 1'h0;
		else if (\mchip.my_core.regB.en )
			\mchip.my_core.regB.Q [2] <= \mchip.my_core.Stack.bus [2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.my_core.regB.Q [3] <= 1'h0;
		else if (\mchip.my_core.regB.en )
			\mchip.my_core.regB.Q [3] <= \mchip.my_core.Stack.bus [3];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.my_core.regB.Q [4] <= 1'h0;
		else if (\mchip.my_core.regB.en )
			\mchip.my_core.regB.Q [4] <= \mchip.my_core.Stack.bus [4];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.my_core.regB.Q [5] <= 1'h0;
		else if (\mchip.my_core.regB.en )
			\mchip.my_core.regB.Q [5] <= \mchip.my_core.Stack.bus [5];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.my_core.regB.Q [6] <= 1'h0;
		else if (\mchip.my_core.regB.en )
			\mchip.my_core.regB.Q [6] <= \mchip.my_core.Stack.bus [6];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.my_core.regB.Q [7] <= 1'h0;
		else if (\mchip.my_core.regB.en )
			\mchip.my_core.regB.Q [7] <= \mchip.my_core.Stack.bus [7];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.my_core.Unit.flag_reg.Q [1] <= 1'h0;
		else if (_0017_)
			\mchip.my_core.Unit.flag_reg.Q [1] <= \mchip.my_core.Unit.flag_reg.d [1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.my_core.Unit.flag_reg.Q [2] <= 1'h0;
		else if (_0017_)
			\mchip.my_core.Unit.flag_reg.Q [2] <= \mchip.my_core.Unit.flag_reg.d [2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.my_core.Unit.flag_reg.Q [3] <= 1'h0;
		else if (_0017_)
			\mchip.my_core.Unit.flag_reg.Q [3] <= \mchip.my_core.Unit.flag_reg.d [3];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.my_core.SP_SEL.Q [0] <= 1'h0;
		else if (!_0062_)
			\mchip.my_core.SP_SEL.Q [0] <= _1498_[0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.my_core.SP_SEL.Q [1] <= 1'h0;
		else if (!_0062_)
			\mchip.my_core.SP_SEL.Q [1] <= _1499_[1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.my_core.SP_SEL.Q [2] <= 1'h0;
		else if (!_0062_)
			\mchip.my_core.SP_SEL.Q [2] <= _1499_[2];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.my_core.Brain.state [0] <= 1'h0;
		else
			\mchip.my_core.Brain.state [0] <= \mchip.my_core.Brain.next_state [0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.my_core.Brain.state [1] <= 1'h1;
		else
			\mchip.my_core.Brain.state [1] <= \mchip.my_core.Brain.next_state [1];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.my_core.Brain.state [2] <= 1'h0;
		else
			\mchip.my_core.Brain.state [2] <= \mchip.my_core.Brain.next_state [2];
	always @(posedge io_in[12])
		if (_0019_)
			\mchip.my_core.S_Intr  <= 1'h0;
		else
			\mchip.my_core.S_Intr  <= io_in[8];
	always @(posedge io_in[12])
		if (_0015_)
			if (!_0047_)
				\mchip.my_core.Stack.rf[1] [0] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[1] [0] <= _0023_;
	always @(posedge io_in[12])
		if (_0015_)
			if (!_0047_)
				\mchip.my_core.Stack.rf[1] [1] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[1] [1] <= _0028_;
	always @(posedge io_in[12])
		if (_0015_)
			if (!_0047_)
				\mchip.my_core.Stack.rf[1] [2] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[1] [2] <= _0029_;
	always @(posedge io_in[12])
		if (_0015_)
			if (!_0047_)
				\mchip.my_core.Stack.rf[1] [3] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[1] [3] <= _0030_;
	always @(posedge io_in[12])
		if (_0015_)
			if (!_0047_)
				\mchip.my_core.Stack.rf[1] [4] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[1] [4] <= _0031_;
	always @(posedge io_in[12])
		if (_0015_)
			if (!_0047_)
				\mchip.my_core.Stack.rf[1] [5] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[1] [5] <= _0032_;
	always @(posedge io_in[12])
		if (_0015_)
			if (!_0047_)
				\mchip.my_core.Stack.rf[1] [6] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[1] [6] <= _0033_;
	always @(posedge io_in[12])
		if (_0015_)
			if (!_0047_)
				\mchip.my_core.Stack.rf[1] [7] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[1] [7] <= _0034_;
	always @(posedge io_in[12])
		if (_0015_)
			if (!_0047_)
				\mchip.my_core.Stack.rf[1] [8] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[1] [8] <= _0035_;
	always @(posedge io_in[12])
		if (_0015_)
			if (!_0047_)
				\mchip.my_core.Stack.rf[1] [9] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[1] [9] <= _0036_;
	always @(posedge io_in[12])
		if (_0015_)
			if (!_0047_)
				\mchip.my_core.Stack.rf[1] [10] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[1] [10] <= _0024_;
	always @(posedge io_in[12])
		if (_0015_)
			if (!_0047_)
				\mchip.my_core.Stack.rf[1] [11] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[1] [11] <= _0025_;
	always @(posedge io_in[12])
		if (_0015_)
			if (!_0047_)
				\mchip.my_core.Stack.rf[1] [12] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[1] [12] <= _0026_;
	always @(posedge io_in[12])
		if (_0015_)
			if (!_0047_)
				\mchip.my_core.Stack.rf[1] [13] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[1] [13] <= _0027_;
	always @(posedge io_in[12]) \mchip.my_core.Brain.cycle [0] <= _0001_;
	always @(posedge io_in[12]) \mchip.my_core.Brain.cycle [1] <= _0002_;
	always @(posedge io_in[12]) \mchip.my_core.Brain.cycle [2] <= _0003_;
	always @(posedge io_in[12])
		if (_0016_)
			if (!_0046_)
				\mchip.my_core.Stack.rf[0] [0] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[0] [0] <= _0023_;
	always @(posedge io_in[12])
		if (_0016_)
			if (!_0046_)
				\mchip.my_core.Stack.rf[0] [1] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[0] [1] <= _0028_;
	always @(posedge io_in[12])
		if (_0016_)
			if (!_0046_)
				\mchip.my_core.Stack.rf[0] [2] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[0] [2] <= _0029_;
	always @(posedge io_in[12])
		if (_0016_)
			if (!_0046_)
				\mchip.my_core.Stack.rf[0] [3] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[0] [3] <= _0030_;
	always @(posedge io_in[12])
		if (_0016_)
			if (!_0046_)
				\mchip.my_core.Stack.rf[0] [4] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[0] [4] <= _0031_;
	always @(posedge io_in[12])
		if (_0016_)
			if (!_0046_)
				\mchip.my_core.Stack.rf[0] [5] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[0] [5] <= _0032_;
	always @(posedge io_in[12])
		if (_0016_)
			if (!_0046_)
				\mchip.my_core.Stack.rf[0] [6] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[0] [6] <= _0033_;
	always @(posedge io_in[12])
		if (_0016_)
			if (!_0046_)
				\mchip.my_core.Stack.rf[0] [7] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[0] [7] <= _0034_;
	always @(posedge io_in[12])
		if (_0016_)
			if (!_0046_)
				\mchip.my_core.Stack.rf[0] [8] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[0] [8] <= _0035_;
	always @(posedge io_in[12])
		if (_0016_)
			if (!_0046_)
				\mchip.my_core.Stack.rf[0] [9] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[0] [9] <= _0036_;
	always @(posedge io_in[12])
		if (_0016_)
			if (!_0046_)
				\mchip.my_core.Stack.rf[0] [10] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[0] [10] <= _0024_;
	always @(posedge io_in[12])
		if (_0016_)
			if (!_0046_)
				\mchip.my_core.Stack.rf[0] [11] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[0] [11] <= _0025_;
	always @(posedge io_in[12])
		if (_0016_)
			if (!_0046_)
				\mchip.my_core.Stack.rf[0] [12] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[0] [12] <= _0026_;
	always @(posedge io_in[12])
		if (_0016_)
			if (!_0046_)
				\mchip.my_core.Stack.rf[0] [13] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[0] [13] <= _0027_;
	always @(posedge io_in[12])
		if (_0014_)
			if (!_0048_)
				\mchip.my_core.Stack.rf[2] [0] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[2] [0] <= _0023_;
	always @(posedge io_in[12])
		if (_0014_)
			if (!_0048_)
				\mchip.my_core.Stack.rf[2] [1] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[2] [1] <= _0028_;
	always @(posedge io_in[12])
		if (_0014_)
			if (!_0048_)
				\mchip.my_core.Stack.rf[2] [2] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[2] [2] <= _0029_;
	always @(posedge io_in[12])
		if (_0014_)
			if (!_0048_)
				\mchip.my_core.Stack.rf[2] [3] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[2] [3] <= _0030_;
	always @(posedge io_in[12])
		if (_0014_)
			if (!_0048_)
				\mchip.my_core.Stack.rf[2] [4] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[2] [4] <= _0031_;
	always @(posedge io_in[12])
		if (_0014_)
			if (!_0048_)
				\mchip.my_core.Stack.rf[2] [5] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[2] [5] <= _0032_;
	always @(posedge io_in[12])
		if (_0014_)
			if (!_0048_)
				\mchip.my_core.Stack.rf[2] [6] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[2] [6] <= _0033_;
	always @(posedge io_in[12])
		if (_0014_)
			if (!_0048_)
				\mchip.my_core.Stack.rf[2] [7] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[2] [7] <= _0034_;
	always @(posedge io_in[12])
		if (_0014_)
			if (!_0048_)
				\mchip.my_core.Stack.rf[2] [8] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[2] [8] <= _0035_;
	always @(posedge io_in[12])
		if (_0014_)
			if (!_0048_)
				\mchip.my_core.Stack.rf[2] [9] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[2] [9] <= _0036_;
	always @(posedge io_in[12])
		if (_0014_)
			if (!_0048_)
				\mchip.my_core.Stack.rf[2] [10] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[2] [10] <= _0024_;
	always @(posedge io_in[12])
		if (_0014_)
			if (!_0048_)
				\mchip.my_core.Stack.rf[2] [11] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[2] [11] <= _0025_;
	always @(posedge io_in[12])
		if (_0014_)
			if (!_0048_)
				\mchip.my_core.Stack.rf[2] [12] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[2] [12] <= _0026_;
	always @(posedge io_in[12])
		if (_0014_)
			if (!_0048_)
				\mchip.my_core.Stack.rf[2] [13] <= 1'h0;
			else
				\mchip.my_core.Stack.rf[2] [13] <= _0027_;
	always @(posedge io_in[12])
		if (_0061_)
			\mchip.my_core.rf.rf[7] [0] <= _0037_;
	always @(posedge io_in[12])
		if (_0061_)
			\mchip.my_core.rf.rf[7] [1] <= _0038_;
	always @(posedge io_in[12])
		if (_0061_)
			\mchip.my_core.rf.rf[7] [2] <= _0039_;
	always @(posedge io_in[12])
		if (_0061_)
			\mchip.my_core.rf.rf[7] [3] <= _0040_;
	always @(posedge io_in[12])
		if (_0061_)
			\mchip.my_core.rf.rf[7] [4] <= _0041_;
	always @(posedge io_in[12])
		if (_0061_)
			\mchip.my_core.rf.rf[7] [5] <= _0042_;
	always @(posedge io_in[12])
		if (_0061_)
			\mchip.my_core.rf.rf[7] [6] <= _0043_;
	always @(posedge io_in[12])
		if (_0061_)
			\mchip.my_core.rf.rf[7] [7] <= _0044_;
	assign _1498_[2:1] = 2'h0;
	assign _1499_[0] = _1498_[0];
	assign io_out = {2'h0, \mchip.my_core.Sync , \mchip.my_core.Brain.state , \mchip.my_core.Stack.bus };
	assign \mchip.clock  = io_in[12];
	assign \mchip.io_in  = io_in[11:0];
	assign \mchip.io_out  = {\mchip.my_core.Sync , \mchip.my_core.Brain.state , \mchip.my_core.Stack.bus };
	assign \mchip.my_core.ACC  = \mchip.my_core.rf.rf[0] ;
	assign \mchip.my_core.A_in  = \mchip.my_core.regA.d ;
	assign \mchip.my_core.A_out  = \mchip.my_core.regA.Q ;
	assign \mchip.my_core.B_out  = \mchip.my_core.regB.Q ;
	assign \mchip.my_core.B_rst  = io_in[13];
	assign \mchip.my_core.Brain.D5_3  = \mchip.my_core.IR.Q [5:3];
	assign \mchip.my_core.Brain.DDD  = \mchip.my_core.IR.Q [5:3];
	assign \mchip.my_core.Brain.Intr  = \mchip.my_core.Intr ;
	assign \mchip.my_core.Brain.Ready  = \mchip.my_core.Ready ;
	assign \mchip.my_core.Brain.SSS  = \mchip.my_core.IR.Q [2:0];
	assign \mchip.my_core.Brain.clk  = io_in[12];
	assign \mchip.my_core.Brain.ctrl_signals  = {1'h0, \mchip.my_core.Sync , 5'h00, \mchip.my_core.A_en , 2'h0, \mchip.my_core.regB.en , 29'h00000000};
	assign \mchip.my_core.Brain.flags  = \mchip.my_core.Unit.flag_reg.Q ;
	assign \mchip.my_core.Brain.instr  = \mchip.my_core.IR.Q ;
	assign \mchip.my_core.Brain.rst  = io_in[13];
	assign \mchip.my_core.D_in  = io_in[7:0];
	assign \mchip.my_core.D_out  = \mchip.my_core.Stack.bus ;
	assign \mchip.my_core.INTR  = io_in[8];
	assign \mchip.my_core.IR.clear  = io_in[13];
	assign \mchip.my_core.IR.clk  = io_in[12];
	assign \mchip.my_core.IR.d  = io_in[7:0];
	assign \mchip.my_core.IR_en  = \mchip.my_core.IR.en ;
	assign \mchip.my_core.IR_rst  = io_in[13];
	assign \mchip.my_core.READY  = io_in[9];
	assign \mchip.my_core.SP_SEL.clear  = io_in[13];
	assign \mchip.my_core.SP_SEL.clk  = io_in[12];
	assign \mchip.my_core.SP_SEL.d  = 3'h0;
	assign \mchip.my_core.SP_SEL.load  = 1'h0;
	assign \mchip.my_core.SP_SEL.up  = 1'h0;
	assign \mchip.my_core.SP_rst  = io_in[13];
	assign \mchip.my_core.Stack.RST_AAA  = {2'h0, \mchip.my_core.Stack.bus [5:3], 3'h0};
	assign \mchip.my_core.Stack.Stack_ctrl  = 7'h00;
	assign \mchip.my_core.Stack.clk  = io_in[12];
	assign \mchip.my_core.Stack.rst  = io_in[13];
	assign \mchip.my_core.Stack.sel  = \mchip.my_core.SP_SEL.Q ;
	assign \mchip.my_core.Stack.upper  = 8'h00;
	assign \mchip.my_core.Unit.ALU_ctrl  = 10'h000;
	assign \mchip.my_core.Unit.Flag_rst  = io_in[13];
	assign \mchip.my_core.Unit.a  = \mchip.my_core.regA.Q ;
	assign \mchip.my_core.Unit.b  = \mchip.my_core.regB.Q ;
	assign \mchip.my_core.Unit.clk  = io_in[12];
	assign \mchip.my_core.Unit.flag_in  = \mchip.my_core.Unit.flag_reg.d ;
	assign \mchip.my_core.Unit.flag_reg.clear  = io_in[13];
	assign \mchip.my_core.Unit.flag_reg.clk  = io_in[12];
	assign \mchip.my_core.Unit.flag_reg.en  = 1'h0;
	assign \mchip.my_core.Unit.flags  = \mchip.my_core.Unit.flag_reg.Q ;
	assign \mchip.my_core.Unit.rst  = io_in[13];
	assign \mchip.my_core.bus  = \mchip.my_core.Stack.bus ;
	assign \mchip.my_core.clk  = io_in[12];
	assign \mchip.my_core.ctrl_signals  = {1'h0, \mchip.my_core.Sync , 5'h00, \mchip.my_core.A_en , 2'h0, \mchip.my_core.regB.en , 29'h00000000};
	assign \mchip.my_core.flags  = \mchip.my_core.Unit.flag_reg.Q ;
	assign \mchip.my_core.instr  = \mchip.my_core.IR.Q ;
	assign \mchip.my_core.regA.clear  = \mchip.my_core.A_rst ;
	assign \mchip.my_core.regA.clk  = io_in[12];
	assign \mchip.my_core.regA.en  = \mchip.my_core.A_en ;
	assign \mchip.my_core.regB.clear  = io_in[13];
	assign \mchip.my_core.regB.clk  = io_in[12];
	assign \mchip.my_core.regB.d  = \mchip.my_core.Stack.bus ;
	assign \mchip.my_core.rf.ACC  = \mchip.my_core.rf.rf[0] ;
	assign \mchip.my_core.rf.bus  = \mchip.my_core.Stack.bus ;
	assign \mchip.my_core.rf.clk  = io_in[12];
	assign \mchip.my_core.rf.rf_ctrl  = 5'h00;
	assign \mchip.my_core.rf.rst  = io_in[13];
	assign \mchip.my_core.rst  = io_in[13];
	assign \mchip.my_core.sel_Stack  = \mchip.my_core.SP_SEL.Q ;
	assign \mchip.my_core.state  = \mchip.my_core.Brain.state ;
	assign \mchip.reset  = io_in[13];
endmodule
module d30_yuchingw_fpga (
	io_in,
	io_out
);
	wire _00_;
	wire _01_;
	wire _02_;
	wire _03_;
	wire _04_;
	wire _05_;
	wire _06_;
	wire _07_;
	wire _08_;
	wire _09_;
	wire _10_;
	wire _11_;
	wire _12_;
	wire _13_;
	wire _14_;
	wire _15_;
	wire _16_;
	wire _17_;
	wire _18_;
	wire _19_;
	wire _20_;
	wire _21_;
	input wire [13:0] io_in;
	output wire [13:0] io_out;
	wire \mchip.clock ;
	wire [11:0] \mchip.io_in ;
	wire [11:0] \mchip.io_out ;
	wire \mchip.reset ;
	wire [4:0] \mchip.setData ;
	wire [15:0] \mchip.top.CLBOut ;
	wire [3:0] \mchip.top.addr0.LUTConfig ;
	wire \mchip.top.addr0.clock ;
	wire [3:0] \mchip.top.addr0.data.D ;
	wire \mchip.top.addr0.data.clock ;
	wire \mchip.top.addr0.data.reset ;
	wire \mchip.top.addr0.dataSel.D ;
	wire \mchip.top.addr0.dataSel.clock ;
	wire \mchip.top.addr0.dataSel.reset ;
	wire \mchip.top.addr0.letVal.clock ;
	wire \mchip.top.addr0.letVal.en ;
	wire \mchip.top.addr0.letVal.reset ;
	wire \mchip.top.addr0.memSel_in ;
	wire \mchip.top.addr0.out ;
	wire \mchip.top.addr0.reset ;
	wire [3:0] \mchip.top.addr1.LUTConfig ;
	wire \mchip.top.addr1.clock ;
	wire [3:0] \mchip.top.addr1.data.D ;
	wire \mchip.top.addr1.data.clock ;
	wire \mchip.top.addr1.data.reset ;
	wire \mchip.top.addr1.dataSel.D ;
	wire \mchip.top.addr1.dataSel.clock ;
	wire \mchip.top.addr1.dataSel.reset ;
	wire \mchip.top.addr1.letVal.clock ;
	wire \mchip.top.addr1.letVal.en ;
	wire \mchip.top.addr1.letVal.reset ;
	wire \mchip.top.addr1.memSel_in ;
	wire \mchip.top.addr1.out ;
	wire \mchip.top.addr1.reset ;
	wire [3:0] \mchip.top.addr10.LUTConfig ;
	wire \mchip.top.addr10.clock ;
	wire [3:0] \mchip.top.addr10.data.D ;
	wire \mchip.top.addr10.data.clock ;
	wire \mchip.top.addr10.data.reset ;
	wire \mchip.top.addr10.dataSel.D ;
	wire \mchip.top.addr10.dataSel.clock ;
	wire \mchip.top.addr10.dataSel.reset ;
	wire \mchip.top.addr10.letVal.clock ;
	wire \mchip.top.addr10.letVal.en ;
	wire \mchip.top.addr10.letVal.reset ;
	wire \mchip.top.addr10.memSel_in ;
	wire \mchip.top.addr10.out ;
	wire \mchip.top.addr10.reset ;
	wire [1:0] \mchip.top.addr10.sel ;
	wire [3:0] \mchip.top.addr11.LUTConfig ;
	wire \mchip.top.addr11.clock ;
	wire [3:0] \mchip.top.addr11.data.D ;
	wire \mchip.top.addr11.data.clock ;
	wire \mchip.top.addr11.data.reset ;
	wire \mchip.top.addr11.dataSel.D ;
	wire \mchip.top.addr11.dataSel.clock ;
	wire \mchip.top.addr11.dataSel.reset ;
	wire \mchip.top.addr11.letVal.clock ;
	wire \mchip.top.addr11.letVal.en ;
	wire \mchip.top.addr11.letVal.reset ;
	wire \mchip.top.addr11.memSel_in ;
	wire \mchip.top.addr11.out ;
	wire \mchip.top.addr11.reset ;
	wire [1:0] \mchip.top.addr11.sel ;
	wire [3:0] \mchip.top.addr12.LUTConfig ;
	wire [3:0] \mchip.top.addr12.LUTData ;
	wire \mchip.top.addr12.clock ;
	wire [3:0] \mchip.top.addr12.data.D ;
	wire [3:0] \mchip.top.addr12.data.Q ;
	wire \mchip.top.addr12.data.clock ;
	wire \mchip.top.addr12.data.reset ;
	wire \mchip.top.addr12.dataSel.D ;
	reg \mchip.top.addr12.dataSel.Q ;
	wire \mchip.top.addr12.dataSel.clock ;
	wire \mchip.top.addr12.dataSel.reset ;
	wire \mchip.top.addr12.letVal.D ;
	reg \mchip.top.addr12.letVal.Q ;
	wire \mchip.top.addr12.letVal.clock ;
	wire \mchip.top.addr12.letVal.en ;
	wire \mchip.top.addr12.letVal.reset ;
	wire \mchip.top.addr12.memSel_in ;
	wire \mchip.top.addr12.memSel_mem ;
	wire \mchip.top.addr12.out ;
	wire \mchip.top.addr12.regData ;
	wire \mchip.top.addr12.reset ;
	wire [1:0] \mchip.top.addr12.sel ;
	wire [3:0] \mchip.top.addr13.LUTConfig ;
	wire [3:0] \mchip.top.addr13.LUTData ;
	wire \mchip.top.addr13.clock ;
	wire [3:0] \mchip.top.addr13.data.D ;
	wire [3:0] \mchip.top.addr13.data.Q ;
	wire \mchip.top.addr13.data.clock ;
	wire \mchip.top.addr13.data.reset ;
	wire \mchip.top.addr13.dataSel.D ;
	reg \mchip.top.addr13.dataSel.Q ;
	wire \mchip.top.addr13.dataSel.clock ;
	wire \mchip.top.addr13.dataSel.reset ;
	wire \mchip.top.addr13.letVal.D ;
	reg \mchip.top.addr13.letVal.Q ;
	wire \mchip.top.addr13.letVal.clock ;
	wire \mchip.top.addr13.letVal.en ;
	wire \mchip.top.addr13.letVal.reset ;
	wire \mchip.top.addr13.memSel_in ;
	wire \mchip.top.addr13.memSel_mem ;
	wire \mchip.top.addr13.out ;
	wire \mchip.top.addr13.regData ;
	wire \mchip.top.addr13.reset ;
	wire [1:0] \mchip.top.addr13.sel ;
	wire [3:0] \mchip.top.addr14.LUTConfig ;
	wire [3:0] \mchip.top.addr14.LUTData ;
	wire \mchip.top.addr14.clock ;
	wire [3:0] \mchip.top.addr14.data.D ;
	wire [3:0] \mchip.top.addr14.data.Q ;
	wire \mchip.top.addr14.data.clock ;
	wire \mchip.top.addr14.data.reset ;
	wire \mchip.top.addr14.dataSel.D ;
	reg \mchip.top.addr14.dataSel.Q ;
	wire \mchip.top.addr14.dataSel.clock ;
	wire \mchip.top.addr14.dataSel.reset ;
	wire \mchip.top.addr14.letVal.D ;
	reg \mchip.top.addr14.letVal.Q ;
	wire \mchip.top.addr14.letVal.clock ;
	wire \mchip.top.addr14.letVal.en ;
	wire \mchip.top.addr14.letVal.reset ;
	wire \mchip.top.addr14.memSel_in ;
	wire \mchip.top.addr14.memSel_mem ;
	wire \mchip.top.addr14.out ;
	wire \mchip.top.addr14.regData ;
	wire \mchip.top.addr14.reset ;
	wire [1:0] \mchip.top.addr14.sel ;
	wire [3:0] \mchip.top.addr15.LUTConfig ;
	wire [3:0] \mchip.top.addr15.LUTData ;
	wire \mchip.top.addr15.clock ;
	wire [3:0] \mchip.top.addr15.data.D ;
	wire [3:0] \mchip.top.addr15.data.Q ;
	wire \mchip.top.addr15.data.clock ;
	wire \mchip.top.addr15.data.reset ;
	wire \mchip.top.addr15.dataSel.D ;
	reg \mchip.top.addr15.dataSel.Q ;
	wire \mchip.top.addr15.dataSel.clock ;
	wire \mchip.top.addr15.dataSel.reset ;
	wire \mchip.top.addr15.letVal.D ;
	reg \mchip.top.addr15.letVal.Q ;
	wire \mchip.top.addr15.letVal.clock ;
	wire \mchip.top.addr15.letVal.en ;
	wire \mchip.top.addr15.letVal.reset ;
	wire \mchip.top.addr15.memSel_in ;
	wire \mchip.top.addr15.memSel_mem ;
	wire \mchip.top.addr15.out ;
	wire \mchip.top.addr15.regData ;
	wire \mchip.top.addr15.reset ;
	wire [1:0] \mchip.top.addr15.sel ;
	wire [3:0] \mchip.top.addr2.LUTConfig ;
	wire \mchip.top.addr2.clock ;
	wire [3:0] \mchip.top.addr2.data.D ;
	wire \mchip.top.addr2.data.clock ;
	wire \mchip.top.addr2.data.reset ;
	wire \mchip.top.addr2.dataSel.D ;
	wire \mchip.top.addr2.dataSel.clock ;
	wire \mchip.top.addr2.dataSel.reset ;
	wire \mchip.top.addr2.letVal.clock ;
	wire \mchip.top.addr2.letVal.en ;
	wire \mchip.top.addr2.letVal.reset ;
	wire \mchip.top.addr2.memSel_in ;
	wire \mchip.top.addr2.out ;
	wire \mchip.top.addr2.reset ;
	wire [3:0] \mchip.top.addr3.LUTConfig ;
	wire \mchip.top.addr3.clock ;
	wire [3:0] \mchip.top.addr3.data.D ;
	wire \mchip.top.addr3.data.clock ;
	wire \mchip.top.addr3.data.reset ;
	wire \mchip.top.addr3.dataSel.D ;
	wire \mchip.top.addr3.dataSel.clock ;
	wire \mchip.top.addr3.dataSel.reset ;
	wire \mchip.top.addr3.letVal.clock ;
	wire \mchip.top.addr3.letVal.en ;
	wire \mchip.top.addr3.letVal.reset ;
	wire \mchip.top.addr3.memSel_in ;
	wire \mchip.top.addr3.out ;
	wire \mchip.top.addr3.reset ;
	wire [3:0] \mchip.top.addr4.LUTConfig ;
	wire \mchip.top.addr4.clock ;
	wire [3:0] \mchip.top.addr4.data.D ;
	wire \mchip.top.addr4.data.clock ;
	wire \mchip.top.addr4.data.reset ;
	wire \mchip.top.addr4.dataSel.D ;
	wire \mchip.top.addr4.dataSel.clock ;
	wire \mchip.top.addr4.dataSel.reset ;
	wire \mchip.top.addr4.letVal.clock ;
	wire \mchip.top.addr4.letVal.en ;
	wire \mchip.top.addr4.letVal.reset ;
	wire \mchip.top.addr4.memSel_in ;
	wire \mchip.top.addr4.out ;
	wire \mchip.top.addr4.reset ;
	wire [1:0] \mchip.top.addr4.sel ;
	wire [3:0] \mchip.top.addr5.LUTConfig ;
	wire \mchip.top.addr5.clock ;
	wire [3:0] \mchip.top.addr5.data.D ;
	wire \mchip.top.addr5.data.clock ;
	wire \mchip.top.addr5.data.reset ;
	wire \mchip.top.addr5.dataSel.D ;
	wire \mchip.top.addr5.dataSel.clock ;
	wire \mchip.top.addr5.dataSel.reset ;
	wire \mchip.top.addr5.letVal.clock ;
	wire \mchip.top.addr5.letVal.en ;
	wire \mchip.top.addr5.letVal.reset ;
	wire \mchip.top.addr5.memSel_in ;
	wire \mchip.top.addr5.out ;
	wire \mchip.top.addr5.reset ;
	wire [1:0] \mchip.top.addr5.sel ;
	wire [3:0] \mchip.top.addr6.LUTConfig ;
	wire \mchip.top.addr6.clock ;
	wire [3:0] \mchip.top.addr6.data.D ;
	wire \mchip.top.addr6.data.clock ;
	wire \mchip.top.addr6.data.reset ;
	wire \mchip.top.addr6.dataSel.D ;
	wire \mchip.top.addr6.dataSel.clock ;
	wire \mchip.top.addr6.dataSel.reset ;
	wire \mchip.top.addr6.letVal.clock ;
	wire \mchip.top.addr6.letVal.en ;
	wire \mchip.top.addr6.letVal.reset ;
	wire \mchip.top.addr6.memSel_in ;
	wire \mchip.top.addr6.out ;
	wire \mchip.top.addr6.reset ;
	wire [1:0] \mchip.top.addr6.sel ;
	wire [3:0] \mchip.top.addr7.LUTConfig ;
	wire \mchip.top.addr7.clock ;
	wire [3:0] \mchip.top.addr7.data.D ;
	wire \mchip.top.addr7.data.clock ;
	wire \mchip.top.addr7.data.reset ;
	wire \mchip.top.addr7.dataSel.D ;
	wire \mchip.top.addr7.dataSel.clock ;
	wire \mchip.top.addr7.dataSel.reset ;
	wire \mchip.top.addr7.letVal.clock ;
	wire \mchip.top.addr7.letVal.en ;
	wire \mchip.top.addr7.letVal.reset ;
	wire \mchip.top.addr7.memSel_in ;
	wire \mchip.top.addr7.out ;
	wire \mchip.top.addr7.reset ;
	wire [1:0] \mchip.top.addr7.sel ;
	wire [3:0] \mchip.top.addr8.LUTConfig ;
	wire \mchip.top.addr8.clock ;
	wire [3:0] \mchip.top.addr8.data.D ;
	wire \mchip.top.addr8.data.clock ;
	wire \mchip.top.addr8.data.reset ;
	wire \mchip.top.addr8.dataSel.D ;
	wire \mchip.top.addr8.dataSel.clock ;
	wire \mchip.top.addr8.dataSel.reset ;
	wire \mchip.top.addr8.letVal.clock ;
	wire \mchip.top.addr8.letVal.en ;
	wire \mchip.top.addr8.letVal.reset ;
	wire \mchip.top.addr8.memSel_in ;
	wire \mchip.top.addr8.out ;
	wire \mchip.top.addr8.reset ;
	wire [1:0] \mchip.top.addr8.sel ;
	wire [3:0] \mchip.top.addr9.LUTConfig ;
	wire \mchip.top.addr9.clock ;
	wire [3:0] \mchip.top.addr9.data.D ;
	wire \mchip.top.addr9.data.clock ;
	wire \mchip.top.addr9.data.reset ;
	wire \mchip.top.addr9.dataSel.D ;
	wire \mchip.top.addr9.dataSel.clock ;
	wire \mchip.top.addr9.dataSel.reset ;
	wire \mchip.top.addr9.letVal.clock ;
	wire \mchip.top.addr9.letVal.en ;
	wire \mchip.top.addr9.letVal.reset ;
	wire \mchip.top.addr9.memSel_in ;
	wire \mchip.top.addr9.out ;
	wire \mchip.top.addr9.reset ;
	wire [1:0] \mchip.top.addr9.sel ;
	wire \mchip.top.clock ;
	wire \mchip.top.inputSel0.clock ;
	wire [1:0] \mchip.top.inputSel0.regInput.D ;
	wire \mchip.top.inputSel0.regInput.clock ;
	wire \mchip.top.inputSel0.regInput.reset ;
	wire \mchip.top.inputSel0.reset ;
	wire [1:0] \mchip.top.inputSel0.selConfig ;
	wire \mchip.top.inputSel1.clock ;
	wire [1:0] \mchip.top.inputSel1.regInput.D ;
	wire \mchip.top.inputSel1.regInput.clock ;
	wire \mchip.top.inputSel1.regInput.reset ;
	wire \mchip.top.inputSel1.reset ;
	wire [1:0] \mchip.top.inputSel1.selConfig ;
	wire \mchip.top.inputSel2.clock ;
	wire [1:0] \mchip.top.inputSel2.regInput.D ;
	wire \mchip.top.inputSel2.regInput.clock ;
	wire \mchip.top.inputSel2.regInput.reset ;
	wire \mchip.top.inputSel2.reset ;
	wire [1:0] \mchip.top.inputSel2.selConfig ;
	wire \mchip.top.inputSel3.clock ;
	wire [1:0] \mchip.top.inputSel3.regInput.D ;
	wire \mchip.top.inputSel3.regInput.clock ;
	wire \mchip.top.inputSel3.regInput.reset ;
	wire \mchip.top.inputSel3.reset ;
	wire [1:0] \mchip.top.inputSel3.selConfig ;
	wire \mchip.top.inputSel4.clock ;
	wire [1:0] \mchip.top.inputSel4.regInput.D ;
	wire \mchip.top.inputSel4.regInput.clock ;
	wire \mchip.top.inputSel4.regInput.reset ;
	wire \mchip.top.inputSel4.reset ;
	wire [1:0] \mchip.top.inputSel4.selConfig ;
	wire \mchip.top.inputSel5.clock ;
	wire [1:0] \mchip.top.inputSel5.regInput.D ;
	wire \mchip.top.inputSel5.regInput.clock ;
	wire \mchip.top.inputSel5.regInput.reset ;
	wire \mchip.top.inputSel5.reset ;
	wire [1:0] \mchip.top.inputSel5.selConfig ;
	wire \mchip.top.inputSel6.clock ;
	wire [1:0] \mchip.top.inputSel6.regInput.D ;
	wire \mchip.top.inputSel6.regInput.clock ;
	wire \mchip.top.inputSel6.regInput.reset ;
	wire \mchip.top.inputSel6.reset ;
	wire [1:0] \mchip.top.inputSel6.selConfig ;
	wire \mchip.top.inputSel7.clock ;
	wire [1:0] \mchip.top.inputSel7.regInput.D ;
	wire \mchip.top.inputSel7.regInput.clock ;
	wire \mchip.top.inputSel7.regInput.reset ;
	wire \mchip.top.inputSel7.reset ;
	wire [1:0] \mchip.top.inputSel7.selConfig ;
	wire [3:0] \mchip.top.out ;
	wire \mchip.top.reset ;
	wire [4:0] \mchip.top.setData ;
	wire \mchip.top.switch16.clock ;
	wire [3:0] \mchip.top.switch16.data.D ;
	wire \mchip.top.switch16.data.clock ;
	wire \mchip.top.switch16.data.reset ;
	wire [11:0] \mchip.top.switch16.inputs ;
	wire \mchip.top.switch16.out ;
	wire \mchip.top.switch16.reset ;
	wire [3:0] \mchip.top.switch16.selectConfig ;
	wire \mchip.top.switch17.clock ;
	wire [3:0] \mchip.top.switch17.data.D ;
	wire \mchip.top.switch17.data.clock ;
	wire \mchip.top.switch17.data.reset ;
	wire [11:0] \mchip.top.switch17.inputs ;
	wire \mchip.top.switch17.out ;
	wire \mchip.top.switch17.reset ;
	wire [3:0] \mchip.top.switch17.selectConfig ;
	wire \mchip.top.switch18.clock ;
	wire [3:0] \mchip.top.switch18.data.D ;
	wire \mchip.top.switch18.data.clock ;
	wire \mchip.top.switch18.data.reset ;
	wire [11:0] \mchip.top.switch18.inputs ;
	wire \mchip.top.switch18.out ;
	wire \mchip.top.switch18.reset ;
	wire [3:0] \mchip.top.switch18.selectConfig ;
	wire \mchip.top.switch19.clock ;
	wire [3:0] \mchip.top.switch19.data.D ;
	wire \mchip.top.switch19.data.clock ;
	wire \mchip.top.switch19.data.reset ;
	wire [11:0] \mchip.top.switch19.inputs ;
	wire \mchip.top.switch19.out ;
	wire \mchip.top.switch19.reset ;
	wire [3:0] \mchip.top.switch19.selectConfig ;
	wire \mchip.top.switch20.clock ;
	wire [3:0] \mchip.top.switch20.data.D ;
	wire \mchip.top.switch20.data.clock ;
	wire \mchip.top.switch20.data.reset ;
	wire [11:0] \mchip.top.switch20.inputs ;
	wire \mchip.top.switch20.out ;
	wire \mchip.top.switch20.reset ;
	wire [3:0] \mchip.top.switch20.selectConfig ;
	wire \mchip.top.switch21.clock ;
	wire [3:0] \mchip.top.switch21.data.D ;
	wire \mchip.top.switch21.data.clock ;
	wire \mchip.top.switch21.data.reset ;
	wire [11:0] \mchip.top.switch21.inputs ;
	wire \mchip.top.switch21.out ;
	wire \mchip.top.switch21.reset ;
	wire [3:0] \mchip.top.switch21.selectConfig ;
	wire \mchip.top.switch22.clock ;
	wire [3:0] \mchip.top.switch22.data.D ;
	wire \mchip.top.switch22.data.clock ;
	wire \mchip.top.switch22.data.reset ;
	wire [11:0] \mchip.top.switch22.inputs ;
	wire \mchip.top.switch22.out ;
	wire \mchip.top.switch22.reset ;
	wire [3:0] \mchip.top.switch22.selectConfig ;
	wire \mchip.top.switch23.clock ;
	wire [3:0] \mchip.top.switch23.data.D ;
	wire \mchip.top.switch23.data.clock ;
	wire \mchip.top.switch23.data.reset ;
	wire [11:0] \mchip.top.switch23.inputs ;
	wire \mchip.top.switch23.out ;
	wire \mchip.top.switch23.reset ;
	wire [3:0] \mchip.top.switch23.selectConfig ;
	wire \mchip.top.switch24.clock ;
	wire [3:0] \mchip.top.switch24.data.D ;
	wire \mchip.top.switch24.data.clock ;
	wire \mchip.top.switch24.data.reset ;
	wire [11:0] \mchip.top.switch24.inputs ;
	wire \mchip.top.switch24.out ;
	wire \mchip.top.switch24.reset ;
	wire [3:0] \mchip.top.switch24.selectConfig ;
	wire \mchip.top.switch25.clock ;
	wire [3:0] \mchip.top.switch25.data.D ;
	wire \mchip.top.switch25.data.clock ;
	wire \mchip.top.switch25.data.reset ;
	wire [11:0] \mchip.top.switch25.inputs ;
	wire \mchip.top.switch25.out ;
	wire \mchip.top.switch25.reset ;
	wire [3:0] \mchip.top.switch25.selectConfig ;
	wire \mchip.top.switch26.clock ;
	wire [3:0] \mchip.top.switch26.data.D ;
	wire \mchip.top.switch26.data.clock ;
	wire \mchip.top.switch26.data.reset ;
	wire [11:0] \mchip.top.switch26.inputs ;
	wire \mchip.top.switch26.out ;
	wire \mchip.top.switch26.reset ;
	wire [3:0] \mchip.top.switch26.selectConfig ;
	wire \mchip.top.switch27.clock ;
	wire [3:0] \mchip.top.switch27.data.D ;
	wire \mchip.top.switch27.data.clock ;
	wire \mchip.top.switch27.data.reset ;
	wire [11:0] \mchip.top.switch27.inputs ;
	wire \mchip.top.switch27.out ;
	wire \mchip.top.switch27.reset ;
	wire [3:0] \mchip.top.switch27.selectConfig ;
	wire \mchip.top.switch28.clock ;
	wire [3:0] \mchip.top.switch28.data.D ;
	wire \mchip.top.switch28.data.clock ;
	wire \mchip.top.switch28.data.reset ;
	wire [11:0] \mchip.top.switch28.inputs ;
	wire \mchip.top.switch28.out ;
	wire \mchip.top.switch28.reset ;
	wire [3:0] \mchip.top.switch28.selectConfig ;
	wire \mchip.top.switch29.clock ;
	wire [3:0] \mchip.top.switch29.data.D ;
	wire \mchip.top.switch29.data.clock ;
	wire \mchip.top.switch29.data.reset ;
	wire [11:0] \mchip.top.switch29.inputs ;
	wire \mchip.top.switch29.out ;
	wire \mchip.top.switch29.reset ;
	wire [3:0] \mchip.top.switch29.selectConfig ;
	wire \mchip.top.switch30.clock ;
	wire [3:0] \mchip.top.switch30.data.D ;
	wire \mchip.top.switch30.data.clock ;
	wire \mchip.top.switch30.data.reset ;
	wire [11:0] \mchip.top.switch30.inputs ;
	wire \mchip.top.switch30.out ;
	wire \mchip.top.switch30.reset ;
	wire [3:0] \mchip.top.switch30.selectConfig ;
	wire \mchip.top.switch31.clock ;
	wire [3:0] \mchip.top.switch31.data.D ;
	wire \mchip.top.switch31.data.clock ;
	wire \mchip.top.switch31.data.reset ;
	wire [11:0] \mchip.top.switch31.inputs ;
	wire \mchip.top.switch31.out ;
	wire \mchip.top.switch31.reset ;
	wire [3:0] \mchip.top.switch31.selectConfig ;
	wire \mchip.top.switch32.clock ;
	wire [3:0] \mchip.top.switch32.data.D ;
	wire \mchip.top.switch32.data.clock ;
	wire \mchip.top.switch32.data.reset ;
	wire [11:0] \mchip.top.switch32.inputs ;
	wire \mchip.top.switch32.out ;
	wire \mchip.top.switch32.reset ;
	wire [3:0] \mchip.top.switch32.selectConfig ;
	wire \mchip.top.switch33.clock ;
	wire [3:0] \mchip.top.switch33.data.D ;
	wire \mchip.top.switch33.data.clock ;
	wire \mchip.top.switch33.data.reset ;
	wire [11:0] \mchip.top.switch33.inputs ;
	wire \mchip.top.switch33.out ;
	wire \mchip.top.switch33.reset ;
	wire [3:0] \mchip.top.switch33.selectConfig ;
	wire \mchip.top.switch34.clock ;
	wire [3:0] \mchip.top.switch34.data.D ;
	wire \mchip.top.switch34.data.clock ;
	wire \mchip.top.switch34.data.reset ;
	wire [11:0] \mchip.top.switch34.inputs ;
	wire \mchip.top.switch34.out ;
	wire \mchip.top.switch34.reset ;
	wire [3:0] \mchip.top.switch34.selectConfig ;
	wire \mchip.top.switch35.clock ;
	wire [3:0] \mchip.top.switch35.data.D ;
	wire \mchip.top.switch35.data.clock ;
	wire \mchip.top.switch35.data.reset ;
	wire [11:0] \mchip.top.switch35.inputs ;
	wire \mchip.top.switch35.out ;
	wire \mchip.top.switch35.reset ;
	wire [3:0] \mchip.top.switch35.selectConfig ;
	wire \mchip.top.switch36.clock ;
	wire [3:0] \mchip.top.switch36.data.D ;
	wire \mchip.top.switch36.data.clock ;
	wire \mchip.top.switch36.data.reset ;
	wire [11:0] \mchip.top.switch36.inputs ;
	wire \mchip.top.switch36.out ;
	wire \mchip.top.switch36.reset ;
	wire [3:0] \mchip.top.switch36.selectConfig ;
	wire \mchip.top.switch37.clock ;
	wire [3:0] \mchip.top.switch37.data.D ;
	wire \mchip.top.switch37.data.clock ;
	wire \mchip.top.switch37.data.reset ;
	wire [11:0] \mchip.top.switch37.inputs ;
	wire \mchip.top.switch37.out ;
	wire \mchip.top.switch37.reset ;
	wire [3:0] \mchip.top.switch37.selectConfig ;
	wire \mchip.top.switch38.clock ;
	wire [3:0] \mchip.top.switch38.data.D ;
	wire \mchip.top.switch38.data.clock ;
	wire \mchip.top.switch38.data.reset ;
	wire [11:0] \mchip.top.switch38.inputs ;
	wire \mchip.top.switch38.out ;
	wire \mchip.top.switch38.reset ;
	wire [3:0] \mchip.top.switch38.selectConfig ;
	wire \mchip.top.switch39.clock ;
	wire [3:0] \mchip.top.switch39.data.D ;
	wire \mchip.top.switch39.data.clock ;
	wire \mchip.top.switch39.data.reset ;
	wire [11:0] \mchip.top.switch39.inputs ;
	wire \mchip.top.switch39.out ;
	wire \mchip.top.switch39.reset ;
	wire [3:0] \mchip.top.switch39.selectConfig ;
	wire [1:0] \mchip.top.switchOut10 ;
	wire [1:0] \mchip.top.switchOut11 ;
	wire [1:0] \mchip.top.switchOut12 ;
	wire [1:0] \mchip.top.switchOut13 ;
	wire [1:0] \mchip.top.switchOut14 ;
	wire [1:0] \mchip.top.switchOut15 ;
	wire [1:0] \mchip.top.switchOut4 ;
	wire [1:0] \mchip.top.switchOut5 ;
	wire [1:0] \mchip.top.switchOut6 ;
	wire [1:0] \mchip.top.switchOut7 ;
	wire [1:0] \mchip.top.switchOut8 ;
	wire [1:0] \mchip.top.switchOut9 ;
	assign _04_ = io_in[11] | ~io_in[0];
	assign _05_ = io_in[10] | ~io_in[0];
	assign _06_ = _05_ | _04_;
	assign _07_ = io_in[0] & ~io_in[9];
	assign _08_ = io_in[0] & ~io_in[8];
	assign _09_ = _08_ | _07_;
	assign _10_ = io_in[7] | ~io_in[0];
	assign _11_ = io_in[6] | ~io_in[0];
	assign _12_ = _11_ | _10_;
	assign _13_ = _12_ | _09_;
	assign _00_ = _13_ | _06_;
	assign _14_ = io_in[0] & ~io_in[6];
	assign _15_ = _14_ | _10_;
	assign _16_ = _15_ | _09_;
	assign _01_ = _16_ | _06_;
	assign _17_ = io_in[0] & ~io_in[7];
	assign _18_ = _11_ | _17_;
	assign _19_ = _18_ | _09_;
	assign _02_ = _19_ | _06_;
	assign _20_ = _14_ | _17_;
	assign _21_ = _20_ | _09_;
	assign _03_ = _21_ | _06_;
	assign \mchip.top.addr12.out  = (\mchip.top.addr12.dataSel.Q  ? \mchip.top.addr12.letVal.Q  : \mchip.top.addr12.data.Q [0]);
	assign \mchip.top.addr13.out  = (\mchip.top.addr13.dataSel.Q  ? \mchip.top.addr13.letVal.Q  : \mchip.top.addr13.data.Q [0]);
	assign \mchip.top.addr14.out  = (\mchip.top.addr14.dataSel.Q  ? \mchip.top.addr14.letVal.Q  : \mchip.top.addr14.data.Q [0]);
	assign \mchip.top.addr15.out  = (\mchip.top.addr15.dataSel.Q  ? \mchip.top.addr15.letVal.Q  : \mchip.top.addr15.data.Q [0]);
	assign \mchip.setData [0] = io_in[1] & io_in[0];
	assign \mchip.top.addr0.dataSel.D  = io_in[5] & io_in[0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.addr15.letVal.Q  <= 1'h0;
		else
			\mchip.top.addr15.letVal.Q  <= \mchip.top.addr15.data.Q [0];
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.addr12.dataSel.Q  <= 1'h0;
		else if (!_00_)
			\mchip.top.addr12.dataSel.Q  <= \mchip.top.addr0.dataSel.D ;
	reg \mchip.top.addr12.data.Q_reg[0] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.addr12.data.Q_reg[0]  <= 1'h0;
		else if (!_00_)
			\mchip.top.addr12.data.Q_reg[0]  <= \mchip.setData [0];
	assign \mchip.top.addr12.data.Q [0] = \mchip.top.addr12.data.Q_reg[0] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.addr13.dataSel.Q  <= 1'h0;
		else if (!_01_)
			\mchip.top.addr13.dataSel.Q  <= \mchip.top.addr0.dataSel.D ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.addr12.letVal.Q  <= 1'h0;
		else
			\mchip.top.addr12.letVal.Q  <= \mchip.top.addr12.data.Q [0];
	reg \mchip.top.addr13.data.Q_reg[0] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.addr13.data.Q_reg[0]  <= 1'h0;
		else if (!_01_)
			\mchip.top.addr13.data.Q_reg[0]  <= \mchip.setData [0];
	assign \mchip.top.addr13.data.Q [0] = \mchip.top.addr13.data.Q_reg[0] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.addr14.dataSel.Q  <= 1'h0;
		else if (!_02_)
			\mchip.top.addr14.dataSel.Q  <= \mchip.top.addr0.dataSel.D ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.addr13.letVal.Q  <= 1'h0;
		else
			\mchip.top.addr13.letVal.Q  <= \mchip.top.addr13.data.Q [0];
	reg \mchip.top.addr14.data.Q_reg[0] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.addr14.data.Q_reg[0]  <= 1'h0;
		else if (!_02_)
			\mchip.top.addr14.data.Q_reg[0]  <= \mchip.setData [0];
	assign \mchip.top.addr14.data.Q [0] = \mchip.top.addr14.data.Q_reg[0] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.addr15.dataSel.Q  <= 1'h0;
		else if (!_03_)
			\mchip.top.addr15.dataSel.Q  <= \mchip.top.addr0.dataSel.D ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.addr14.letVal.Q  <= 1'h0;
		else
			\mchip.top.addr14.letVal.Q  <= \mchip.top.addr14.data.Q [0];
	reg \mchip.top.addr15.data.Q_reg[0] ;
	always @(posedge io_in[12])
		if (io_in[13])
			\mchip.top.addr15.data.Q_reg[0]  <= 1'h0;
		else if (!_03_)
			\mchip.top.addr15.data.Q_reg[0]  <= \mchip.setData [0];
	assign \mchip.top.addr15.data.Q [0] = \mchip.top.addr15.data.Q_reg[0] ;
	assign io_out = {10'h000, \mchip.top.addr15.out , \mchip.top.addr14.out , \mchip.top.addr13.out , \mchip.top.addr12.out };
	assign \mchip.clock  = io_in[12];
	assign \mchip.io_in  = io_in[11:0];
	assign \mchip.io_out  = {8'h00, \mchip.top.addr15.out , \mchip.top.addr14.out , \mchip.top.addr13.out , \mchip.top.addr12.out };
	assign \mchip.reset  = io_in[13];
	assign \mchip.setData [4:1] = {\mchip.top.addr0.dataSel.D , 3'h0};
	assign \mchip.top.CLBOut  = {\mchip.top.addr15.out , \mchip.top.addr14.out , \mchip.top.addr13.out , \mchip.top.addr12.out , 12'h000};
	assign \mchip.top.addr0.LUTConfig  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.addr0.clock  = io_in[12];
	assign \mchip.top.addr0.data.D  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.addr0.data.clock  = io_in[12];
	assign \mchip.top.addr0.data.reset  = io_in[13];
	assign \mchip.top.addr0.dataSel.clock  = io_in[12];
	assign \mchip.top.addr0.dataSel.reset  = io_in[13];
	assign \mchip.top.addr0.letVal.clock  = io_in[12];
	assign \mchip.top.addr0.letVal.en  = 1'h1;
	assign \mchip.top.addr0.letVal.reset  = io_in[13];
	assign \mchip.top.addr0.memSel_in  = \mchip.top.addr0.dataSel.D ;
	assign \mchip.top.addr0.out  = 1'h0;
	assign \mchip.top.addr0.reset  = io_in[13];
	assign \mchip.top.addr1.LUTConfig  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.addr1.clock  = io_in[12];
	assign \mchip.top.addr1.data.D  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.addr1.data.clock  = io_in[12];
	assign \mchip.top.addr1.data.reset  = io_in[13];
	assign \mchip.top.addr1.dataSel.D  = \mchip.top.addr0.dataSel.D ;
	assign \mchip.top.addr1.dataSel.clock  = io_in[12];
	assign \mchip.top.addr1.dataSel.reset  = io_in[13];
	assign \mchip.top.addr1.letVal.clock  = io_in[12];
	assign \mchip.top.addr1.letVal.en  = 1'h1;
	assign \mchip.top.addr1.letVal.reset  = io_in[13];
	assign \mchip.top.addr1.memSel_in  = \mchip.top.addr0.dataSel.D ;
	assign \mchip.top.addr1.out  = 1'h0;
	assign \mchip.top.addr1.reset  = io_in[13];
	assign \mchip.top.addr10.LUTConfig  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.addr10.clock  = io_in[12];
	assign \mchip.top.addr10.data.D  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.addr10.data.clock  = io_in[12];
	assign \mchip.top.addr10.data.reset  = io_in[13];
	assign \mchip.top.addr10.dataSel.D  = \mchip.top.addr0.dataSel.D ;
	assign \mchip.top.addr10.dataSel.clock  = io_in[12];
	assign \mchip.top.addr10.dataSel.reset  = io_in[13];
	assign \mchip.top.addr10.letVal.clock  = io_in[12];
	assign \mchip.top.addr10.letVal.en  = 1'h1;
	assign \mchip.top.addr10.letVal.reset  = io_in[13];
	assign \mchip.top.addr10.memSel_in  = \mchip.top.addr0.dataSel.D ;
	assign \mchip.top.addr10.out  = 1'h0;
	assign \mchip.top.addr10.reset  = io_in[13];
	assign \mchip.top.addr10.sel  = {\mchip.top.addr12.out , \mchip.top.addr12.out };
	assign \mchip.top.addr11.LUTConfig  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.addr11.clock  = io_in[12];
	assign \mchip.top.addr11.data.D  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.addr11.data.clock  = io_in[12];
	assign \mchip.top.addr11.data.reset  = io_in[13];
	assign \mchip.top.addr11.dataSel.D  = \mchip.top.addr0.dataSel.D ;
	assign \mchip.top.addr11.dataSel.clock  = io_in[12];
	assign \mchip.top.addr11.dataSel.reset  = io_in[13];
	assign \mchip.top.addr11.letVal.clock  = io_in[12];
	assign \mchip.top.addr11.letVal.en  = 1'h1;
	assign \mchip.top.addr11.letVal.reset  = io_in[13];
	assign \mchip.top.addr11.memSel_in  = \mchip.top.addr0.dataSel.D ;
	assign \mchip.top.addr11.out  = 1'h0;
	assign \mchip.top.addr11.reset  = io_in[13];
	assign \mchip.top.addr11.sel  = {\mchip.top.addr12.out , \mchip.top.addr12.out };
	assign \mchip.top.addr12.LUTConfig  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.addr12.LUTData  = {3'h0, \mchip.top.addr12.data.Q [0]};
	assign \mchip.top.addr12.clock  = io_in[12];
	assign \mchip.top.addr12.data.D  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.addr12.data.Q [3:1] = 3'h0;
	assign \mchip.top.addr12.data.clock  = io_in[12];
	assign \mchip.top.addr12.data.reset  = io_in[13];
	assign \mchip.top.addr12.dataSel.D  = \mchip.top.addr0.dataSel.D ;
	assign \mchip.top.addr12.dataSel.clock  = io_in[12];
	assign \mchip.top.addr12.dataSel.reset  = io_in[13];
	assign \mchip.top.addr12.letVal.D  = \mchip.top.addr12.data.Q [0];
	assign \mchip.top.addr12.letVal.clock  = io_in[12];
	assign \mchip.top.addr12.letVal.en  = 1'h1;
	assign \mchip.top.addr12.letVal.reset  = io_in[13];
	assign \mchip.top.addr12.memSel_in  = \mchip.top.addr0.dataSel.D ;
	assign \mchip.top.addr12.memSel_mem  = \mchip.top.addr12.dataSel.Q ;
	assign \mchip.top.addr12.regData  = \mchip.top.addr12.letVal.Q ;
	assign \mchip.top.addr12.reset  = io_in[13];
	assign \mchip.top.addr12.sel  = 2'h0;
	assign \mchip.top.addr13.LUTConfig  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.addr13.LUTData  = {3'h0, \mchip.top.addr13.data.Q [0]};
	assign \mchip.top.addr13.clock  = io_in[12];
	assign \mchip.top.addr13.data.D  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.addr13.data.Q [3:1] = 3'h0;
	assign \mchip.top.addr13.data.clock  = io_in[12];
	assign \mchip.top.addr13.data.reset  = io_in[13];
	assign \mchip.top.addr13.dataSel.D  = \mchip.top.addr0.dataSel.D ;
	assign \mchip.top.addr13.dataSel.clock  = io_in[12];
	assign \mchip.top.addr13.dataSel.reset  = io_in[13];
	assign \mchip.top.addr13.letVal.D  = \mchip.top.addr13.data.Q [0];
	assign \mchip.top.addr13.letVal.clock  = io_in[12];
	assign \mchip.top.addr13.letVal.en  = 1'h1;
	assign \mchip.top.addr13.letVal.reset  = io_in[13];
	assign \mchip.top.addr13.memSel_in  = \mchip.top.addr0.dataSel.D ;
	assign \mchip.top.addr13.memSel_mem  = \mchip.top.addr13.dataSel.Q ;
	assign \mchip.top.addr13.regData  = \mchip.top.addr13.letVal.Q ;
	assign \mchip.top.addr13.reset  = io_in[13];
	assign \mchip.top.addr13.sel  = 2'h0;
	assign \mchip.top.addr14.LUTConfig  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.addr14.LUTData  = {3'h0, \mchip.top.addr14.data.Q [0]};
	assign \mchip.top.addr14.clock  = io_in[12];
	assign \mchip.top.addr14.data.D  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.addr14.data.Q [3:1] = 3'h0;
	assign \mchip.top.addr14.data.clock  = io_in[12];
	assign \mchip.top.addr14.data.reset  = io_in[13];
	assign \mchip.top.addr14.dataSel.D  = \mchip.top.addr0.dataSel.D ;
	assign \mchip.top.addr14.dataSel.clock  = io_in[12];
	assign \mchip.top.addr14.dataSel.reset  = io_in[13];
	assign \mchip.top.addr14.letVal.D  = \mchip.top.addr14.data.Q [0];
	assign \mchip.top.addr14.letVal.clock  = io_in[12];
	assign \mchip.top.addr14.letVal.en  = 1'h1;
	assign \mchip.top.addr14.letVal.reset  = io_in[13];
	assign \mchip.top.addr14.memSel_in  = \mchip.top.addr0.dataSel.D ;
	assign \mchip.top.addr14.memSel_mem  = \mchip.top.addr14.dataSel.Q ;
	assign \mchip.top.addr14.regData  = \mchip.top.addr14.letVal.Q ;
	assign \mchip.top.addr14.reset  = io_in[13];
	assign \mchip.top.addr14.sel  = 2'h0;
	assign \mchip.top.addr15.LUTConfig  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.addr15.LUTData  = {3'h0, \mchip.top.addr15.data.Q [0]};
	assign \mchip.top.addr15.clock  = io_in[12];
	assign \mchip.top.addr15.data.D  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.addr15.data.Q [3:1] = 3'h0;
	assign \mchip.top.addr15.data.clock  = io_in[12];
	assign \mchip.top.addr15.data.reset  = io_in[13];
	assign \mchip.top.addr15.dataSel.D  = \mchip.top.addr0.dataSel.D ;
	assign \mchip.top.addr15.dataSel.clock  = io_in[12];
	assign \mchip.top.addr15.dataSel.reset  = io_in[13];
	assign \mchip.top.addr15.letVal.D  = \mchip.top.addr15.data.Q [0];
	assign \mchip.top.addr15.letVal.clock  = io_in[12];
	assign \mchip.top.addr15.letVal.en  = 1'h1;
	assign \mchip.top.addr15.letVal.reset  = io_in[13];
	assign \mchip.top.addr15.memSel_in  = \mchip.top.addr0.dataSel.D ;
	assign \mchip.top.addr15.memSel_mem  = \mchip.top.addr15.dataSel.Q ;
	assign \mchip.top.addr15.regData  = \mchip.top.addr15.letVal.Q ;
	assign \mchip.top.addr15.reset  = io_in[13];
	assign \mchip.top.addr15.sel  = 2'h0;
	assign \mchip.top.addr2.LUTConfig  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.addr2.clock  = io_in[12];
	assign \mchip.top.addr2.data.D  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.addr2.data.clock  = io_in[12];
	assign \mchip.top.addr2.data.reset  = io_in[13];
	assign \mchip.top.addr2.dataSel.D  = \mchip.top.addr0.dataSel.D ;
	assign \mchip.top.addr2.dataSel.clock  = io_in[12];
	assign \mchip.top.addr2.dataSel.reset  = io_in[13];
	assign \mchip.top.addr2.letVal.clock  = io_in[12];
	assign \mchip.top.addr2.letVal.en  = 1'h1;
	assign \mchip.top.addr2.letVal.reset  = io_in[13];
	assign \mchip.top.addr2.memSel_in  = \mchip.top.addr0.dataSel.D ;
	assign \mchip.top.addr2.out  = 1'h0;
	assign \mchip.top.addr2.reset  = io_in[13];
	assign \mchip.top.addr3.LUTConfig  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.addr3.clock  = io_in[12];
	assign \mchip.top.addr3.data.D  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.addr3.data.clock  = io_in[12];
	assign \mchip.top.addr3.data.reset  = io_in[13];
	assign \mchip.top.addr3.dataSel.D  = \mchip.top.addr0.dataSel.D ;
	assign \mchip.top.addr3.dataSel.clock  = io_in[12];
	assign \mchip.top.addr3.dataSel.reset  = io_in[13];
	assign \mchip.top.addr3.letVal.clock  = io_in[12];
	assign \mchip.top.addr3.letVal.en  = 1'h1;
	assign \mchip.top.addr3.letVal.reset  = io_in[13];
	assign \mchip.top.addr3.memSel_in  = \mchip.top.addr0.dataSel.D ;
	assign \mchip.top.addr3.out  = 1'h0;
	assign \mchip.top.addr3.reset  = io_in[13];
	assign \mchip.top.addr4.LUTConfig  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.addr4.clock  = io_in[12];
	assign \mchip.top.addr4.data.D  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.addr4.data.clock  = io_in[12];
	assign \mchip.top.addr4.data.reset  = io_in[13];
	assign \mchip.top.addr4.dataSel.D  = \mchip.top.addr0.dataSel.D ;
	assign \mchip.top.addr4.dataSel.clock  = io_in[12];
	assign \mchip.top.addr4.dataSel.reset  = io_in[13];
	assign \mchip.top.addr4.letVal.clock  = io_in[12];
	assign \mchip.top.addr4.letVal.en  = 1'h1;
	assign \mchip.top.addr4.letVal.reset  = io_in[13];
	assign \mchip.top.addr4.memSel_in  = \mchip.top.addr0.dataSel.D ;
	assign \mchip.top.addr4.out  = 1'h0;
	assign \mchip.top.addr4.reset  = io_in[13];
	assign \mchip.top.addr4.sel  = 2'h0;
	assign \mchip.top.addr5.LUTConfig  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.addr5.clock  = io_in[12];
	assign \mchip.top.addr5.data.D  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.addr5.data.clock  = io_in[12];
	assign \mchip.top.addr5.data.reset  = io_in[13];
	assign \mchip.top.addr5.dataSel.D  = \mchip.top.addr0.dataSel.D ;
	assign \mchip.top.addr5.dataSel.clock  = io_in[12];
	assign \mchip.top.addr5.dataSel.reset  = io_in[13];
	assign \mchip.top.addr5.letVal.clock  = io_in[12];
	assign \mchip.top.addr5.letVal.en  = 1'h1;
	assign \mchip.top.addr5.letVal.reset  = io_in[13];
	assign \mchip.top.addr5.memSel_in  = \mchip.top.addr0.dataSel.D ;
	assign \mchip.top.addr5.out  = 1'h0;
	assign \mchip.top.addr5.reset  = io_in[13];
	assign \mchip.top.addr5.sel  = 2'h0;
	assign \mchip.top.addr6.LUTConfig  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.addr6.clock  = io_in[12];
	assign \mchip.top.addr6.data.D  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.addr6.data.clock  = io_in[12];
	assign \mchip.top.addr6.data.reset  = io_in[13];
	assign \mchip.top.addr6.dataSel.D  = \mchip.top.addr0.dataSel.D ;
	assign \mchip.top.addr6.dataSel.clock  = io_in[12];
	assign \mchip.top.addr6.dataSel.reset  = io_in[13];
	assign \mchip.top.addr6.letVal.clock  = io_in[12];
	assign \mchip.top.addr6.letVal.en  = 1'h1;
	assign \mchip.top.addr6.letVal.reset  = io_in[13];
	assign \mchip.top.addr6.memSel_in  = \mchip.top.addr0.dataSel.D ;
	assign \mchip.top.addr6.out  = 1'h0;
	assign \mchip.top.addr6.reset  = io_in[13];
	assign \mchip.top.addr6.sel  = 2'h0;
	assign \mchip.top.addr7.LUTConfig  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.addr7.clock  = io_in[12];
	assign \mchip.top.addr7.data.D  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.addr7.data.clock  = io_in[12];
	assign \mchip.top.addr7.data.reset  = io_in[13];
	assign \mchip.top.addr7.dataSel.D  = \mchip.top.addr0.dataSel.D ;
	assign \mchip.top.addr7.dataSel.clock  = io_in[12];
	assign \mchip.top.addr7.dataSel.reset  = io_in[13];
	assign \mchip.top.addr7.letVal.clock  = io_in[12];
	assign \mchip.top.addr7.letVal.en  = 1'h1;
	assign \mchip.top.addr7.letVal.reset  = io_in[13];
	assign \mchip.top.addr7.memSel_in  = \mchip.top.addr0.dataSel.D ;
	assign \mchip.top.addr7.out  = 1'h0;
	assign \mchip.top.addr7.reset  = io_in[13];
	assign \mchip.top.addr7.sel  = 2'h0;
	assign \mchip.top.addr8.LUTConfig  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.addr8.clock  = io_in[12];
	assign \mchip.top.addr8.data.D  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.addr8.data.clock  = io_in[12];
	assign \mchip.top.addr8.data.reset  = io_in[13];
	assign \mchip.top.addr8.dataSel.D  = \mchip.top.addr0.dataSel.D ;
	assign \mchip.top.addr8.dataSel.clock  = io_in[12];
	assign \mchip.top.addr8.dataSel.reset  = io_in[13];
	assign \mchip.top.addr8.letVal.clock  = io_in[12];
	assign \mchip.top.addr8.letVal.en  = 1'h1;
	assign \mchip.top.addr8.letVal.reset  = io_in[13];
	assign \mchip.top.addr8.memSel_in  = \mchip.top.addr0.dataSel.D ;
	assign \mchip.top.addr8.out  = 1'h0;
	assign \mchip.top.addr8.reset  = io_in[13];
	assign \mchip.top.addr8.sel  = {\mchip.top.addr12.out , \mchip.top.addr12.out };
	assign \mchip.top.addr9.LUTConfig  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.addr9.clock  = io_in[12];
	assign \mchip.top.addr9.data.D  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.addr9.data.clock  = io_in[12];
	assign \mchip.top.addr9.data.reset  = io_in[13];
	assign \mchip.top.addr9.dataSel.D  = \mchip.top.addr0.dataSel.D ;
	assign \mchip.top.addr9.dataSel.clock  = io_in[12];
	assign \mchip.top.addr9.dataSel.reset  = io_in[13];
	assign \mchip.top.addr9.letVal.clock  = io_in[12];
	assign \mchip.top.addr9.letVal.en  = 1'h1;
	assign \mchip.top.addr9.letVal.reset  = io_in[13];
	assign \mchip.top.addr9.memSel_in  = \mchip.top.addr0.dataSel.D ;
	assign \mchip.top.addr9.out  = 1'h0;
	assign \mchip.top.addr9.reset  = io_in[13];
	assign \mchip.top.addr9.sel  = {\mchip.top.addr12.out , \mchip.top.addr12.out };
	assign \mchip.top.clock  = io_in[12];
	assign \mchip.top.inputSel0.clock  = io_in[12];
	assign \mchip.top.inputSel0.regInput.D  = {1'h0, \mchip.setData [0]};
	assign \mchip.top.inputSel0.regInput.clock  = io_in[12];
	assign \mchip.top.inputSel0.regInput.reset  = io_in[13];
	assign \mchip.top.inputSel0.reset  = io_in[13];
	assign \mchip.top.inputSel0.selConfig  = {1'h0, \mchip.setData [0]};
	assign \mchip.top.inputSel1.clock  = io_in[12];
	assign \mchip.top.inputSel1.regInput.D  = {1'h0, \mchip.setData [0]};
	assign \mchip.top.inputSel1.regInput.clock  = io_in[12];
	assign \mchip.top.inputSel1.regInput.reset  = io_in[13];
	assign \mchip.top.inputSel1.reset  = io_in[13];
	assign \mchip.top.inputSel1.selConfig  = {1'h0, \mchip.setData [0]};
	assign \mchip.top.inputSel2.clock  = io_in[12];
	assign \mchip.top.inputSel2.regInput.D  = {1'h0, \mchip.setData [0]};
	assign \mchip.top.inputSel2.regInput.clock  = io_in[12];
	assign \mchip.top.inputSel2.regInput.reset  = io_in[13];
	assign \mchip.top.inputSel2.reset  = io_in[13];
	assign \mchip.top.inputSel2.selConfig  = {1'h0, \mchip.setData [0]};
	assign \mchip.top.inputSel3.clock  = io_in[12];
	assign \mchip.top.inputSel3.regInput.D  = {1'h0, \mchip.setData [0]};
	assign \mchip.top.inputSel3.regInput.clock  = io_in[12];
	assign \mchip.top.inputSel3.regInput.reset  = io_in[13];
	assign \mchip.top.inputSel3.reset  = io_in[13];
	assign \mchip.top.inputSel3.selConfig  = {1'h0, \mchip.setData [0]};
	assign \mchip.top.inputSel4.clock  = io_in[12];
	assign \mchip.top.inputSel4.regInput.D  = {1'h0, \mchip.setData [0]};
	assign \mchip.top.inputSel4.regInput.clock  = io_in[12];
	assign \mchip.top.inputSel4.regInput.reset  = io_in[13];
	assign \mchip.top.inputSel4.reset  = io_in[13];
	assign \mchip.top.inputSel4.selConfig  = {1'h0, \mchip.setData [0]};
	assign \mchip.top.inputSel5.clock  = io_in[12];
	assign \mchip.top.inputSel5.regInput.D  = {1'h0, \mchip.setData [0]};
	assign \mchip.top.inputSel5.regInput.clock  = io_in[12];
	assign \mchip.top.inputSel5.regInput.reset  = io_in[13];
	assign \mchip.top.inputSel5.reset  = io_in[13];
	assign \mchip.top.inputSel5.selConfig  = {1'h0, \mchip.setData [0]};
	assign \mchip.top.inputSel6.clock  = io_in[12];
	assign \mchip.top.inputSel6.regInput.D  = {1'h0, \mchip.setData [0]};
	assign \mchip.top.inputSel6.regInput.clock  = io_in[12];
	assign \mchip.top.inputSel6.regInput.reset  = io_in[13];
	assign \mchip.top.inputSel6.reset  = io_in[13];
	assign \mchip.top.inputSel6.selConfig  = {1'h0, \mchip.setData [0]};
	assign \mchip.top.inputSel7.clock  = io_in[12];
	assign \mchip.top.inputSel7.regInput.D  = {1'h0, \mchip.setData [0]};
	assign \mchip.top.inputSel7.regInput.clock  = io_in[12];
	assign \mchip.top.inputSel7.regInput.reset  = io_in[13];
	assign \mchip.top.inputSel7.reset  = io_in[13];
	assign \mchip.top.inputSel7.selConfig  = {1'h0, \mchip.setData [0]};
	assign \mchip.top.out  = {\mchip.top.addr15.out , \mchip.top.addr14.out , \mchip.top.addr13.out , \mchip.top.addr12.out };
	assign \mchip.top.reset  = io_in[13];
	assign \mchip.top.setData  = {\mchip.top.addr0.dataSel.D , 3'h0, \mchip.setData [0]};
	assign \mchip.top.switch16.clock  = io_in[12];
	assign \mchip.top.switch16.data.D  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.switch16.data.clock  = io_in[12];
	assign \mchip.top.switch16.data.reset  = io_in[13];
	assign \mchip.top.switch16.inputs  = 12'h000;
	assign \mchip.top.switch16.out  = 1'h0;
	assign \mchip.top.switch16.reset  = io_in[13];
	assign \mchip.top.switch16.selectConfig  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.switch17.clock  = io_in[12];
	assign \mchip.top.switch17.data.D  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.switch17.data.clock  = io_in[12];
	assign \mchip.top.switch17.data.reset  = io_in[13];
	assign \mchip.top.switch17.inputs  = 12'h000;
	assign \mchip.top.switch17.out  = 1'h0;
	assign \mchip.top.switch17.reset  = io_in[13];
	assign \mchip.top.switch17.selectConfig  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.switch18.clock  = io_in[12];
	assign \mchip.top.switch18.data.D  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.switch18.data.clock  = io_in[12];
	assign \mchip.top.switch18.data.reset  = io_in[13];
	assign \mchip.top.switch18.inputs  = 12'h000;
	assign \mchip.top.switch18.out  = 1'h0;
	assign \mchip.top.switch18.reset  = io_in[13];
	assign \mchip.top.switch18.selectConfig  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.switch19.clock  = io_in[12];
	assign \mchip.top.switch19.data.D  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.switch19.data.clock  = io_in[12];
	assign \mchip.top.switch19.data.reset  = io_in[13];
	assign \mchip.top.switch19.inputs  = 12'h000;
	assign \mchip.top.switch19.out  = 1'h0;
	assign \mchip.top.switch19.reset  = io_in[13];
	assign \mchip.top.switch19.selectConfig  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.switch20.clock  = io_in[12];
	assign \mchip.top.switch20.data.D  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.switch20.data.clock  = io_in[12];
	assign \mchip.top.switch20.data.reset  = io_in[13];
	assign \mchip.top.switch20.inputs  = 12'h000;
	assign \mchip.top.switch20.out  = 1'h0;
	assign \mchip.top.switch20.reset  = io_in[13];
	assign \mchip.top.switch20.selectConfig  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.switch21.clock  = io_in[12];
	assign \mchip.top.switch21.data.D  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.switch21.data.clock  = io_in[12];
	assign \mchip.top.switch21.data.reset  = io_in[13];
	assign \mchip.top.switch21.inputs  = 12'h000;
	assign \mchip.top.switch21.out  = 1'h0;
	assign \mchip.top.switch21.reset  = io_in[13];
	assign \mchip.top.switch21.selectConfig  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.switch22.clock  = io_in[12];
	assign \mchip.top.switch22.data.D  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.switch22.data.clock  = io_in[12];
	assign \mchip.top.switch22.data.reset  = io_in[13];
	assign \mchip.top.switch22.inputs  = 12'h000;
	assign \mchip.top.switch22.out  = 1'h0;
	assign \mchip.top.switch22.reset  = io_in[13];
	assign \mchip.top.switch22.selectConfig  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.switch23.clock  = io_in[12];
	assign \mchip.top.switch23.data.D  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.switch23.data.clock  = io_in[12];
	assign \mchip.top.switch23.data.reset  = io_in[13];
	assign \mchip.top.switch23.inputs  = 12'h000;
	assign \mchip.top.switch23.out  = 1'h0;
	assign \mchip.top.switch23.reset  = io_in[13];
	assign \mchip.top.switch23.selectConfig  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.switch24.clock  = io_in[12];
	assign \mchip.top.switch24.data.D  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.switch24.data.clock  = io_in[12];
	assign \mchip.top.switch24.data.reset  = io_in[13];
	assign \mchip.top.switch24.inputs  = {\mchip.top.addr15.out , \mchip.top.addr14.out , \mchip.top.addr13.out , \mchip.top.addr12.out , 8'h00};
	assign \mchip.top.switch24.out  = \mchip.top.addr12.out ;
	assign \mchip.top.switch24.reset  = io_in[13];
	assign \mchip.top.switch24.selectConfig  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.switch25.clock  = io_in[12];
	assign \mchip.top.switch25.data.D  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.switch25.data.clock  = io_in[12];
	assign \mchip.top.switch25.data.reset  = io_in[13];
	assign \mchip.top.switch25.inputs  = {\mchip.top.addr15.out , \mchip.top.addr14.out , \mchip.top.addr13.out , \mchip.top.addr12.out , 8'h00};
	assign \mchip.top.switch25.out  = \mchip.top.addr12.out ;
	assign \mchip.top.switch25.reset  = io_in[13];
	assign \mchip.top.switch25.selectConfig  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.switch26.clock  = io_in[12];
	assign \mchip.top.switch26.data.D  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.switch26.data.clock  = io_in[12];
	assign \mchip.top.switch26.data.reset  = io_in[13];
	assign \mchip.top.switch26.inputs  = {\mchip.top.addr15.out , \mchip.top.addr14.out , \mchip.top.addr13.out , \mchip.top.addr12.out , 8'h00};
	assign \mchip.top.switch26.out  = \mchip.top.addr12.out ;
	assign \mchip.top.switch26.reset  = io_in[13];
	assign \mchip.top.switch26.selectConfig  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.switch27.clock  = io_in[12];
	assign \mchip.top.switch27.data.D  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.switch27.data.clock  = io_in[12];
	assign \mchip.top.switch27.data.reset  = io_in[13];
	assign \mchip.top.switch27.inputs  = {\mchip.top.addr15.out , \mchip.top.addr14.out , \mchip.top.addr13.out , \mchip.top.addr12.out , 8'h00};
	assign \mchip.top.switch27.out  = \mchip.top.addr12.out ;
	assign \mchip.top.switch27.reset  = io_in[13];
	assign \mchip.top.switch27.selectConfig  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.switch28.clock  = io_in[12];
	assign \mchip.top.switch28.data.D  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.switch28.data.clock  = io_in[12];
	assign \mchip.top.switch28.data.reset  = io_in[13];
	assign \mchip.top.switch28.inputs  = {\mchip.top.addr15.out , \mchip.top.addr14.out , \mchip.top.addr13.out , \mchip.top.addr12.out , 8'h00};
	assign \mchip.top.switch28.out  = \mchip.top.addr12.out ;
	assign \mchip.top.switch28.reset  = io_in[13];
	assign \mchip.top.switch28.selectConfig  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.switch29.clock  = io_in[12];
	assign \mchip.top.switch29.data.D  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.switch29.data.clock  = io_in[12];
	assign \mchip.top.switch29.data.reset  = io_in[13];
	assign \mchip.top.switch29.inputs  = {\mchip.top.addr15.out , \mchip.top.addr14.out , \mchip.top.addr13.out , \mchip.top.addr12.out , 8'h00};
	assign \mchip.top.switch29.out  = \mchip.top.addr12.out ;
	assign \mchip.top.switch29.reset  = io_in[13];
	assign \mchip.top.switch29.selectConfig  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.switch30.clock  = io_in[12];
	assign \mchip.top.switch30.data.D  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.switch30.data.clock  = io_in[12];
	assign \mchip.top.switch30.data.reset  = io_in[13];
	assign \mchip.top.switch30.inputs  = {\mchip.top.addr15.out , \mchip.top.addr14.out , \mchip.top.addr13.out , \mchip.top.addr12.out , 8'h00};
	assign \mchip.top.switch30.out  = \mchip.top.addr12.out ;
	assign \mchip.top.switch30.reset  = io_in[13];
	assign \mchip.top.switch30.selectConfig  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.switch31.clock  = io_in[12];
	assign \mchip.top.switch31.data.D  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.switch31.data.clock  = io_in[12];
	assign \mchip.top.switch31.data.reset  = io_in[13];
	assign \mchip.top.switch31.inputs  = {\mchip.top.addr15.out , \mchip.top.addr14.out , \mchip.top.addr13.out , \mchip.top.addr12.out , 8'h00};
	assign \mchip.top.switch31.out  = \mchip.top.addr12.out ;
	assign \mchip.top.switch31.reset  = io_in[13];
	assign \mchip.top.switch31.selectConfig  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.switch32.clock  = io_in[12];
	assign \mchip.top.switch32.data.D  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.switch32.data.clock  = io_in[12];
	assign \mchip.top.switch32.data.reset  = io_in[13];
	assign \mchip.top.switch32.inputs  = {4'h0, \mchip.top.addr15.out , \mchip.top.addr14.out , \mchip.top.addr13.out , \mchip.top.addr12.out , 4'h0};
	assign \mchip.top.switch32.out  = 1'h0;
	assign \mchip.top.switch32.reset  = io_in[13];
	assign \mchip.top.switch32.selectConfig  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.switch33.clock  = io_in[12];
	assign \mchip.top.switch33.data.D  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.switch33.data.clock  = io_in[12];
	assign \mchip.top.switch33.data.reset  = io_in[13];
	assign \mchip.top.switch33.inputs  = {4'h0, \mchip.top.addr15.out , \mchip.top.addr14.out , \mchip.top.addr13.out , \mchip.top.addr12.out , 4'h0};
	assign \mchip.top.switch33.out  = 1'h0;
	assign \mchip.top.switch33.reset  = io_in[13];
	assign \mchip.top.switch33.selectConfig  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.switch34.clock  = io_in[12];
	assign \mchip.top.switch34.data.D  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.switch34.data.clock  = io_in[12];
	assign \mchip.top.switch34.data.reset  = io_in[13];
	assign \mchip.top.switch34.inputs  = {4'h0, \mchip.top.addr15.out , \mchip.top.addr14.out , \mchip.top.addr13.out , \mchip.top.addr12.out , 4'h0};
	assign \mchip.top.switch34.out  = 1'h0;
	assign \mchip.top.switch34.reset  = io_in[13];
	assign \mchip.top.switch34.selectConfig  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.switch35.clock  = io_in[12];
	assign \mchip.top.switch35.data.D  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.switch35.data.clock  = io_in[12];
	assign \mchip.top.switch35.data.reset  = io_in[13];
	assign \mchip.top.switch35.inputs  = {4'h0, \mchip.top.addr15.out , \mchip.top.addr14.out , \mchip.top.addr13.out , \mchip.top.addr12.out , 4'h0};
	assign \mchip.top.switch35.out  = 1'h0;
	assign \mchip.top.switch35.reset  = io_in[13];
	assign \mchip.top.switch35.selectConfig  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.switch36.clock  = io_in[12];
	assign \mchip.top.switch36.data.D  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.switch36.data.clock  = io_in[12];
	assign \mchip.top.switch36.data.reset  = io_in[13];
	assign \mchip.top.switch36.inputs  = {4'h0, \mchip.top.addr15.out , \mchip.top.addr14.out , \mchip.top.addr13.out , \mchip.top.addr12.out , 4'h0};
	assign \mchip.top.switch36.out  = 1'h0;
	assign \mchip.top.switch36.reset  = io_in[13];
	assign \mchip.top.switch36.selectConfig  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.switch37.clock  = io_in[12];
	assign \mchip.top.switch37.data.D  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.switch37.data.clock  = io_in[12];
	assign \mchip.top.switch37.data.reset  = io_in[13];
	assign \mchip.top.switch37.inputs  = {4'h0, \mchip.top.addr15.out , \mchip.top.addr14.out , \mchip.top.addr13.out , \mchip.top.addr12.out , 4'h0};
	assign \mchip.top.switch37.out  = 1'h0;
	assign \mchip.top.switch37.reset  = io_in[13];
	assign \mchip.top.switch37.selectConfig  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.switch38.clock  = io_in[12];
	assign \mchip.top.switch38.data.D  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.switch38.data.clock  = io_in[12];
	assign \mchip.top.switch38.data.reset  = io_in[13];
	assign \mchip.top.switch38.inputs  = {4'h0, \mchip.top.addr15.out , \mchip.top.addr14.out , \mchip.top.addr13.out , \mchip.top.addr12.out , 4'h0};
	assign \mchip.top.switch38.out  = 1'h0;
	assign \mchip.top.switch38.reset  = io_in[13];
	assign \mchip.top.switch38.selectConfig  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.switch39.clock  = io_in[12];
	assign \mchip.top.switch39.data.D  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.switch39.data.clock  = io_in[12];
	assign \mchip.top.switch39.data.reset  = io_in[13];
	assign \mchip.top.switch39.inputs  = {4'h0, \mchip.top.addr15.out , \mchip.top.addr14.out , \mchip.top.addr13.out , \mchip.top.addr12.out , 4'h0};
	assign \mchip.top.switch39.out  = 1'h0;
	assign \mchip.top.switch39.reset  = io_in[13];
	assign \mchip.top.switch39.selectConfig  = {3'h0, \mchip.setData [0]};
	assign \mchip.top.switchOut10  = {\mchip.top.addr12.out , \mchip.top.addr12.out };
	assign \mchip.top.switchOut11  = {\mchip.top.addr12.out , \mchip.top.addr12.out };
	assign \mchip.top.switchOut12  = 2'h0;
	assign \mchip.top.switchOut13  = 2'h0;
	assign \mchip.top.switchOut14  = 2'h0;
	assign \mchip.top.switchOut15  = 2'h0;
	assign \mchip.top.switchOut4  = 2'h0;
	assign \mchip.top.switchOut5  = 2'h0;
	assign \mchip.top.switchOut6  = 2'h0;
	assign \mchip.top.switchOut7  = 2'h0;
	assign \mchip.top.switchOut8  = {\mchip.top.addr12.out , \mchip.top.addr12.out };
	assign \mchip.top.switchOut9  = {\mchip.top.addr12.out , \mchip.top.addr12.out };
endmodule
module d31_mdhamank_lfsr (
	io_in,
	io_out
);
	wire _00_;
	wire _01_;
	wire _02_;
	input wire [13:0] io_in;
	output wire [13:0] io_out;
	wire \mchip.flipflop1.clk ;
	wire \mchip.flipflop1.d ;
	reg \mchip.flipflop1.q ;
	wire \mchip.flipflop10.clk ;
	reg \mchip.flipflop10.q ;
	wire \mchip.flipflop11.clk ;
	reg \mchip.flipflop11.q ;
	wire \mchip.flipflop12.clk ;
	reg \mchip.flipflop12.q ;
	wire \mchip.flipflop13.clk ;
	reg \mchip.flipflop13.q ;
	wire \mchip.flipflop14.clk ;
	reg \mchip.flipflop14.q ;
	wire \mchip.flipflop15.clk ;
	reg \mchip.flipflop15.q ;
	wire \mchip.flipflop16.clk ;
	reg \mchip.flipflop16.q ;
	wire \mchip.flipflop2.clk ;
	wire \mchip.flipflop2.d ;
	reg \mchip.flipflop2.q ;
	wire \mchip.flipflop3.clk ;
	wire \mchip.flipflop3.d ;
	reg \mchip.flipflop3.q ;
	wire \mchip.flipflop4.clk ;
	wire \mchip.flipflop4.d ;
	wire \mchip.flipflop4.notq ;
	reg \mchip.flipflop4.q ;
	wire \mchip.flipflop5.clk ;
	wire \mchip.flipflop5.d ;
	reg \mchip.flipflop5.q ;
	wire \mchip.flipflop6.clk ;
	wire \mchip.flipflop6.d ;
	wire \mchip.flipflop6.notq ;
	reg \mchip.flipflop6.q ;
	wire \mchip.flipflop7.clk ;
	wire \mchip.flipflop7.d ;
	reg \mchip.flipflop7.q ;
	wire \mchip.flipflop8.clk ;
	wire \mchip.flipflop8.d ;
	reg \mchip.flipflop8.q ;
	wire \mchip.flipflop9.clk ;
	reg \mchip.flipflop9.q ;
	wire \mchip.gate5.in ;
	wire [7:0] \mchip.io_in ;
	wire [7:0] \mchip.io_out ;
	wire \mchip.mux1.out ;
	wire \mchip.mux1.sel ;
	wire \mchip.mux2.a ;
	wire \mchip.mux2.b ;
	wire \mchip.mux2.sel ;
	wire \mchip.mux3.a ;
	wire \mchip.mux3.b ;
	wire \mchip.mux3.sel ;
	wire \mchip.mux4.a ;
	wire \mchip.mux4.b ;
	wire \mchip.mux4.sel ;
	wire \mchip.mux5.a ;
	wire \mchip.mux5.b ;
	wire \mchip.mux5.sel ;
	wire \mchip.mux6.a ;
	wire \mchip.mux6.b ;
	wire \mchip.mux6.sel ;
	wire \mchip.mux7.a ;
	wire \mchip.mux7.b ;
	wire \mchip.mux7.sel ;
	wire \mchip.mux8.a ;
	wire \mchip.mux8.b ;
	wire \mchip.mux8.sel ;
	wire \mchip.mux9.a ;
	wire \mchip.mux9.b ;
	wire \mchip.mux9.sel ;
	wire \mchip.net1 ;
	wire \mchip.net10 ;
	wire \mchip.net11 ;
	wire \mchip.net12 ;
	wire \mchip.net13 ;
	wire \mchip.net15 ;
	wire \mchip.net16 ;
	wire \mchip.net17 ;
	wire \mchip.net18 ;
	wire \mchip.net19 ;
	wire \mchip.net2 ;
	wire \mchip.net20 ;
	wire \mchip.net21 ;
	wire \mchip.net22 ;
	wire \mchip.net23 ;
	wire \mchip.net24 ;
	wire \mchip.net25 ;
	wire \mchip.net26 ;
	wire \mchip.net3 ;
	wire \mchip.net4 ;
	wire \mchip.net5 ;
	wire \mchip.net6 ;
	wire \mchip.net7 ;
	wire \mchip.net8 ;
	wire \mchip.net9 ;
	wire \mchip.xor2.a ;
	wire \mchip.xor2.b ;
	wire \mchip.xor3.a ;
	wire \mchip.xor3.b ;
	assign \mchip.flipflop8.d  = ~\mchip.flipflop6.q ;
	assign \mchip.flipflop5.d  = ~\mchip.flipflop4.q ;
	assign _00_ = \mchip.flipflop7.q  ^ \mchip.flipflop8.q ;
	assign _01_ = \mchip.flipflop5.q  ^ \mchip.flipflop4.q ;
	assign _02_ = ~(_01_ ^ _00_);
	assign \mchip.flipflop2.d  = ~(_02_ & io_in[1]);
	always @(posedge io_in[0])
		if (!io_in[2])
			\mchip.flipflop14.q  <= \mchip.flipflop6.q ;
	always @(posedge io_in[0])
		if (!io_in[2])
			\mchip.flipflop13.q  <= \mchip.flipflop5.q ;
	always @(posedge io_in[0])
		if (!io_in[2])
			\mchip.flipflop12.q  <= \mchip.flipflop4.q ;
	always @(posedge io_in[0])
		if (!io_in[2])
			\mchip.flipflop11.q  <= \mchip.flipflop3.q ;
	always @(posedge io_in[0])
		if (!io_in[2])
			\mchip.flipflop10.q  <= \mchip.flipflop1.q ;
	always @(posedge io_in[0])
		if (!io_in[2])
			\mchip.flipflop16.q  <= \mchip.flipflop8.q ;
	always @(posedge io_in[0]) \mchip.flipflop8.q  <= \mchip.flipflop8.d ;
	always @(posedge io_in[0]) \mchip.flipflop7.q  <= \mchip.flipflop5.q ;
	always @(posedge io_in[0]) \mchip.flipflop6.q  <= \mchip.flipflop7.q ;
	always @(posedge io_in[0]) \mchip.flipflop5.q  <= \mchip.flipflop5.d ;
	always @(posedge io_in[0]) \mchip.flipflop4.q  <= \mchip.flipflop1.q ;
	always @(posedge io_in[0]) \mchip.flipflop3.q  <= \mchip.flipflop2.q ;
	always @(posedge io_in[0]) \mchip.flipflop1.q  <= \mchip.flipflop3.q ;
	always @(posedge io_in[0]) \mchip.flipflop2.q  <= \mchip.flipflop2.d ;
	always @(posedge io_in[0])
		if (!io_in[2])
			\mchip.flipflop9.q  <= \mchip.flipflop2.q ;
	always @(posedge io_in[0])
		if (!io_in[2])
			\mchip.flipflop15.q  <= \mchip.flipflop7.q ;
	assign io_out = {6'h00, \mchip.flipflop16.q , \mchip.flipflop14.q , \mchip.flipflop15.q , \mchip.flipflop13.q , \mchip.flipflop12.q , \mchip.flipflop10.q , \mchip.flipflop11.q , \mchip.flipflop9.q };
	assign \mchip.flipflop1.clk  = io_in[0];
	assign \mchip.flipflop1.d  = \mchip.flipflop3.q ;
	assign \mchip.flipflop10.clk  = io_in[0];
	assign \mchip.flipflop11.clk  = io_in[0];
	assign \mchip.flipflop12.clk  = io_in[0];
	assign \mchip.flipflop13.clk  = io_in[0];
	assign \mchip.flipflop14.clk  = io_in[0];
	assign \mchip.flipflop15.clk  = io_in[0];
	assign \mchip.flipflop16.clk  = io_in[0];
	assign \mchip.flipflop2.clk  = io_in[0];
	assign \mchip.flipflop3.clk  = io_in[0];
	assign \mchip.flipflop3.d  = \mchip.flipflop2.q ;
	assign \mchip.flipflop4.clk  = io_in[0];
	assign \mchip.flipflop4.d  = \mchip.flipflop1.q ;
	assign \mchip.flipflop4.notq  = \mchip.flipflop5.d ;
	assign \mchip.flipflop5.clk  = io_in[0];
	assign \mchip.flipflop6.clk  = io_in[0];
	assign \mchip.flipflop6.d  = \mchip.flipflop7.q ;
	assign \mchip.flipflop6.notq  = \mchip.flipflop8.d ;
	assign \mchip.flipflop7.clk  = io_in[0];
	assign \mchip.flipflop7.d  = \mchip.flipflop5.q ;
	assign \mchip.flipflop8.clk  = io_in[0];
	assign \mchip.flipflop9.clk  = io_in[0];
	assign \mchip.gate5.in  = io_in[1];
	assign \mchip.io_in  = io_in[7:0];
	assign \mchip.io_out  = {\mchip.flipflop16.q , \mchip.flipflop14.q , \mchip.flipflop15.q , \mchip.flipflop13.q , \mchip.flipflop12.q , \mchip.flipflop10.q , \mchip.flipflop11.q , \mchip.flipflop9.q };
	assign \mchip.mux1.out  = \mchip.flipflop2.d ;
	assign \mchip.mux1.sel  = io_in[1];
	assign \mchip.mux2.a  = \mchip.flipflop2.q ;
	assign \mchip.mux2.b  = \mchip.flipflop9.q ;
	assign \mchip.mux2.sel  = io_in[2];
	assign \mchip.mux3.a  = \mchip.flipflop3.q ;
	assign \mchip.mux3.b  = \mchip.flipflop11.q ;
	assign \mchip.mux3.sel  = io_in[2];
	assign \mchip.mux4.a  = \mchip.flipflop1.q ;
	assign \mchip.mux4.b  = \mchip.flipflop10.q ;
	assign \mchip.mux4.sel  = io_in[2];
	assign \mchip.mux5.a  = \mchip.flipflop4.q ;
	assign \mchip.mux5.b  = \mchip.flipflop12.q ;
	assign \mchip.mux5.sel  = io_in[2];
	assign \mchip.mux6.a  = \mchip.flipflop5.q ;
	assign \mchip.mux6.b  = \mchip.flipflop13.q ;
	assign \mchip.mux6.sel  = io_in[2];
	assign \mchip.mux7.a  = \mchip.flipflop7.q ;
	assign \mchip.mux7.b  = \mchip.flipflop15.q ;
	assign \mchip.mux7.sel  = io_in[2];
	assign \mchip.mux8.a  = \mchip.flipflop6.q ;
	assign \mchip.mux8.b  = \mchip.flipflop14.q ;
	assign \mchip.mux8.sel  = io_in[2];
	assign \mchip.mux9.a  = \mchip.flipflop8.q ;
	assign \mchip.mux9.b  = \mchip.flipflop16.q ;
	assign \mchip.mux9.sel  = io_in[2];
	assign \mchip.net1  = io_in[0];
	assign \mchip.net10  = \mchip.flipflop14.q ;
	assign \mchip.net11  = \mchip.flipflop16.q ;
	assign \mchip.net12  = 1'h0;
	assign \mchip.net13  = 1'h1;
	assign \mchip.net15  = 1'h1;
	assign \mchip.net16  = \mchip.flipflop2.d ;
	assign \mchip.net17  = \mchip.flipflop2.q ;
	assign \mchip.net18  = \mchip.flipflop3.q ;
	assign \mchip.net19  = \mchip.flipflop1.q ;
	assign \mchip.net2  = io_in[1];
	assign \mchip.net20  = \mchip.flipflop4.q ;
	assign \mchip.net21  = \mchip.flipflop5.d ;
	assign \mchip.net22  = \mchip.flipflop5.q ;
	assign \mchip.net23  = \mchip.flipflop7.q ;
	assign \mchip.net24  = \mchip.flipflop6.q ;
	assign \mchip.net25  = \mchip.flipflop8.d ;
	assign \mchip.net26  = \mchip.flipflop8.q ;
	assign \mchip.net3  = io_in[2];
	assign \mchip.net4  = \mchip.flipflop9.q ;
	assign \mchip.net5  = \mchip.flipflop11.q ;
	assign \mchip.net6  = \mchip.flipflop10.q ;
	assign \mchip.net7  = \mchip.flipflop12.q ;
	assign \mchip.net8  = \mchip.flipflop13.q ;
	assign \mchip.net9  = \mchip.flipflop15.q ;
	assign \mchip.xor2.a  = \mchip.flipflop7.q ;
	assign \mchip.xor2.b  = \mchip.flipflop8.q ;
	assign \mchip.xor3.a  = \mchip.flipflop4.q ;
	assign \mchip.xor3.b  = \mchip.flipflop5.q ;
endmodule
module d32_ngaertne_cpu (
	io_in,
	io_out
);
	wire _0000_;
	wire _0001_;
	wire _0002_;
	wire _0003_;
	wire _0004_;
	wire _0005_;
	wire _0006_;
	wire _0007_;
	wire _0008_;
	wire _0009_;
	wire _0010_;
	wire _0011_;
	wire _0012_;
	wire _0013_;
	wire _0014_;
	wire _0015_;
	wire _0016_;
	wire _0017_;
	wire _0018_;
	wire _0019_;
	wire _0020_;
	wire _0021_;
	wire _0022_;
	wire _0023_;
	wire _0024_;
	wire _0025_;
	wire _0026_;
	wire _0027_;
	wire _0028_;
	wire _0029_;
	wire _0030_;
	wire _0031_;
	wire _0032_;
	wire _0033_;
	wire _0034_;
	wire _0035_;
	wire _0036_;
	wire _0037_;
	wire _0038_;
	wire _0039_;
	wire _0040_;
	wire _0041_;
	wire _0042_;
	wire _0043_;
	wire _0044_;
	wire _0045_;
	wire _0046_;
	wire _0047_;
	wire _0048_;
	wire _0049_;
	wire _0050_;
	wire _0051_;
	wire _0052_;
	wire _0053_;
	wire _0054_;
	wire _0055_;
	wire _0056_;
	wire _0057_;
	wire _0058_;
	wire _0059_;
	wire _0060_;
	wire _0061_;
	wire _0062_;
	wire _0063_;
	wire _0064_;
	wire _0065_;
	wire _0066_;
	wire _0067_;
	wire _0068_;
	wire _0069_;
	wire _0070_;
	wire _0071_;
	wire _0072_;
	wire _0073_;
	wire _0074_;
	wire _0075_;
	wire _0076_;
	wire _0077_;
	wire _0078_;
	wire _0079_;
	wire _0080_;
	wire _0081_;
	wire _0082_;
	wire _0083_;
	wire _0084_;
	wire _0085_;
	wire _0086_;
	wire _0087_;
	wire _0088_;
	wire _0089_;
	wire _0090_;
	wire _0091_;
	wire _0092_;
	wire _0093_;
	wire _0094_;
	wire _0095_;
	wire _0096_;
	wire _0097_;
	wire _0098_;
	wire _0099_;
	wire _0100_;
	wire _0101_;
	wire _0102_;
	wire _0103_;
	wire _0104_;
	wire _0105_;
	wire _0106_;
	wire _0107_;
	wire _0108_;
	wire _0109_;
	wire _0110_;
	wire _0111_;
	wire _0112_;
	wire _0113_;
	wire _0114_;
	wire _0115_;
	wire _0116_;
	wire _0117_;
	wire _0118_;
	wire _0119_;
	wire _0120_;
	wire _0121_;
	wire _0122_;
	wire _0123_;
	wire _0124_;
	wire _0125_;
	wire _0126_;
	wire _0127_;
	wire _0128_;
	wire _0129_;
	wire _0130_;
	wire _0131_;
	wire _0132_;
	wire _0133_;
	wire _0134_;
	wire _0135_;
	wire _0136_;
	wire _0137_;
	wire _0138_;
	wire _0139_;
	wire _0140_;
	wire _0141_;
	wire _0142_;
	wire _0143_;
	wire _0144_;
	wire _0145_;
	wire _0146_;
	wire _0147_;
	wire _0148_;
	wire _0149_;
	wire _0150_;
	wire _0151_;
	wire _0152_;
	wire _0153_;
	wire _0154_;
	wire _0155_;
	wire _0156_;
	wire _0157_;
	wire _0158_;
	wire _0159_;
	wire _0160_;
	wire _0161_;
	wire _0162_;
	wire _0163_;
	wire _0164_;
	wire _0165_;
	wire _0166_;
	wire _0167_;
	wire _0168_;
	wire _0169_;
	wire _0170_;
	wire _0171_;
	wire _0172_;
	wire _0173_;
	wire _0174_;
	wire _0175_;
	wire _0176_;
	wire _0177_;
	wire _0178_;
	wire _0179_;
	wire _0180_;
	wire _0181_;
	wire _0182_;
	wire _0183_;
	wire _0184_;
	wire _0185_;
	wire _0186_;
	wire _0187_;
	wire _0188_;
	wire _0189_;
	wire _0190_;
	wire _0191_;
	wire _0192_;
	wire _0193_;
	wire _0194_;
	wire _0195_;
	wire _0196_;
	wire _0197_;
	wire _0198_;
	wire _0199_;
	wire _0200_;
	wire _0201_;
	wire _0202_;
	wire _0203_;
	wire _0204_;
	wire _0205_;
	wire _0206_;
	wire _0207_;
	wire _0208_;
	wire _0209_;
	wire _0210_;
	wire _0211_;
	wire _0212_;
	wire _0213_;
	wire _0214_;
	wire _0215_;
	wire _0216_;
	wire _0217_;
	wire _0218_;
	wire _0219_;
	wire _0220_;
	wire _0221_;
	wire _0222_;
	wire _0223_;
	wire _0224_;
	wire _0225_;
	wire _0226_;
	wire _0227_;
	wire _0228_;
	wire _0229_;
	wire _0230_;
	wire _0231_;
	wire _0232_;
	wire _0233_;
	wire _0234_;
	wire _0235_;
	wire _0236_;
	wire _0237_;
	wire _0238_;
	wire _0239_;
	wire _0240_;
	wire _0241_;
	wire _0242_;
	wire _0243_;
	wire _0244_;
	wire _0245_;
	wire _0246_;
	wire _0247_;
	wire _0248_;
	wire _0249_;
	wire _0250_;
	wire _0251_;
	wire _0252_;
	wire _0253_;
	wire _0254_;
	wire _0255_;
	wire _0256_;
	wire _0257_;
	wire _0258_;
	wire _0259_;
	wire _0260_;
	wire _0261_;
	wire _0262_;
	wire _0263_;
	wire _0264_;
	wire _0265_;
	wire _0266_;
	wire _0267_;
	wire _0268_;
	wire _0269_;
	wire _0270_;
	wire _0271_;
	wire _0272_;
	wire _0273_;
	wire _0274_;
	wire _0275_;
	wire _0276_;
	wire _0277_;
	wire _0278_;
	wire _0279_;
	wire _0280_;
	wire _0281_;
	wire _0282_;
	wire _0283_;
	wire _0284_;
	wire _0285_;
	wire _0286_;
	wire _0287_;
	wire _0288_;
	wire _0289_;
	wire _0290_;
	wire _0291_;
	wire _0292_;
	wire _0293_;
	wire _0294_;
	wire _0295_;
	wire _0296_;
	wire _0297_;
	wire _0298_;
	wire _0299_;
	wire _0300_;
	wire _0301_;
	wire _0302_;
	wire _0303_;
	wire _0304_;
	wire _0305_;
	wire _0306_;
	wire _0307_;
	wire _0308_;
	wire _0309_;
	wire _0310_;
	wire _0311_;
	wire _0312_;
	wire _0313_;
	wire _0314_;
	wire _0315_;
	wire _0316_;
	wire _0317_;
	wire _0318_;
	wire _0319_;
	wire _0320_;
	wire _0321_;
	wire _0322_;
	wire _0323_;
	wire _0324_;
	wire _0325_;
	wire _0326_;
	wire _0327_;
	wire _0328_;
	wire _0329_;
	wire _0330_;
	wire _0331_;
	wire _0332_;
	wire _0333_;
	wire _0334_;
	wire _0335_;
	wire _0336_;
	wire _0337_;
	wire _0338_;
	wire _0339_;
	wire _0340_;
	wire _0341_;
	wire _0342_;
	wire _0343_;
	wire _0344_;
	wire _0345_;
	wire _0346_;
	wire _0347_;
	wire _0348_;
	wire _0349_;
	wire _0350_;
	wire _0351_;
	wire _0352_;
	wire _0353_;
	wire _0354_;
	wire _0355_;
	wire _0356_;
	wire _0357_;
	wire _0358_;
	wire _0359_;
	wire _0360_;
	wire _0361_;
	wire _0362_;
	wire _0363_;
	wire _0364_;
	wire _0365_;
	wire _0366_;
	wire _0367_;
	wire _0368_;
	wire _0369_;
	wire _0370_;
	wire _0371_;
	wire _0372_;
	wire _0373_;
	wire _0374_;
	wire _0375_;
	wire _0376_;
	wire _0377_;
	wire _0378_;
	wire _0379_;
	wire _0380_;
	wire _0381_;
	wire _0382_;
	wire _0383_;
	wire _0384_;
	wire _0385_;
	wire _0386_;
	wire _0387_;
	wire _0388_;
	wire _0389_;
	wire _0390_;
	wire _0391_;
	wire _0392_;
	wire _0393_;
	wire _0394_;
	wire _0395_;
	wire _0396_;
	wire _0397_;
	wire _0398_;
	wire _0399_;
	wire _0400_;
	wire _0401_;
	wire _0402_;
	wire _0403_;
	wire _0404_;
	wire _0405_;
	wire _0406_;
	wire _0407_;
	wire _0408_;
	wire _0409_;
	wire _0410_;
	wire _0411_;
	wire _0412_;
	wire _0413_;
	wire _0414_;
	wire _0415_;
	wire _0416_;
	wire _0417_;
	wire _0418_;
	wire _0419_;
	wire _0420_;
	wire _0421_;
	wire _0422_;
	wire _0423_;
	wire _0424_;
	wire _0425_;
	wire _0426_;
	wire _0427_;
	wire _0428_;
	wire _0429_;
	wire _0430_;
	wire _0431_;
	wire _0432_;
	wire _0433_;
	wire _0434_;
	wire _0435_;
	wire _0436_;
	wire _0437_;
	wire _0438_;
	wire _0439_;
	wire _0440_;
	wire _0441_;
	wire _0442_;
	wire _0443_;
	wire _0444_;
	wire _0445_;
	wire _0446_;
	wire _0447_;
	wire _0448_;
	wire _0449_;
	wire _0450_;
	wire _0451_;
	wire _0452_;
	wire _0453_;
	wire _0454_;
	wire _0455_;
	wire _0456_;
	wire _0457_;
	wire _0458_;
	wire _0459_;
	wire _0460_;
	wire _0461_;
	wire _0462_;
	wire _0463_;
	wire _0464_;
	wire _0465_;
	wire _0466_;
	wire _0467_;
	wire _0468_;
	wire _0469_;
	wire _0470_;
	wire _0471_;
	wire _0472_;
	wire _0473_;
	wire _0474_;
	wire _0475_;
	wire _0476_;
	wire _0477_;
	wire _0478_;
	wire _0479_;
	wire _0480_;
	wire _0481_;
	wire _0482_;
	wire _0483_;
	wire _0484_;
	wire _0485_;
	wire _0486_;
	wire _0487_;
	wire _0488_;
	wire _0489_;
	wire _0490_;
	wire _0491_;
	wire _0492_;
	wire _0493_;
	wire _0494_;
	wire _0495_;
	wire [3:0] _0496_;
	wire [3:0] _0497_;
	input wire [13:0] io_in;
	output wire [13:0] io_out;
	wire \mchip.clock ;
	reg [3:0] \mchip.data[0] ;
	reg [3:0] \mchip.data[10] ;
	reg [3:0] \mchip.data[11] ;
	reg [3:0] \mchip.data[12] ;
	reg [3:0] \mchip.data[13] ;
	reg [3:0] \mchip.data[14] ;
	reg [3:0] \mchip.data[15] ;
	reg [3:0] \mchip.data[1] ;
	reg [3:0] \mchip.data[2] ;
	reg [3:0] \mchip.data[3] ;
	reg [3:0] \mchip.data[4] ;
	reg [3:0] \mchip.data[5] ;
	reg [3:0] \mchip.data[6] ;
	reg [3:0] \mchip.data[7] ;
	reg [3:0] \mchip.data[8] ;
	reg [3:0] \mchip.data[9] ;
	wire [3:0] \mchip.inputdata ;
	wire [1:0] \mchip.instruction ;
	wire [7:0] \mchip.io_in ;
	wire [7:0] \mchip.io_out ;
	reg \mchip.lastdata3 ;
	reg [3:0] \mchip.pc ;
	reg [3:0] \mchip.prog[0] ;
	reg [3:0] \mchip.prog[10] ;
	reg [3:0] \mchip.prog[11] ;
	reg [3:0] \mchip.prog[12] ;
	reg [3:0] \mchip.prog[13] ;
	reg [3:0] \mchip.prog[14] ;
	reg [3:0] \mchip.prog[15] ;
	reg [3:0] \mchip.prog[1] ;
	reg [3:0] \mchip.prog[2] ;
	reg [3:0] \mchip.prog[3] ;
	reg [3:0] \mchip.prog[4] ;
	reg [3:0] \mchip.prog[5] ;
	reg [3:0] \mchip.prog[6] ;
	reg [3:0] \mchip.prog[7] ;
	reg [3:0] \mchip.prog[8] ;
	reg [3:0] \mchip.prog[9] ;
	reg [3:0] \mchip.regval ;
	wire \mchip.reset ;
	assign _0037_ = io_in[2] & io_in[3];
	assign _0038_ = ~\mchip.pc [3];
	assign _0039_ = ~\mchip.pc [2];
	assign _0040_ = ~\mchip.pc [1];
	assign _0041_ = (\mchip.pc [0] ? \mchip.prog[1] [1] : \mchip.prog[0] [1]);
	assign _0042_ = (\mchip.pc [0] ? \mchip.prog[3] [1] : \mchip.prog[2] [1]);
	assign _0043_ = (\mchip.pc [1] ? _0042_ : _0041_);
	assign _0044_ = (\mchip.pc [0] ? \mchip.prog[5] [1] : \mchip.prog[4] [1]);
	assign _0045_ = (\mchip.pc [0] ? \mchip.prog[7] [1] : \mchip.prog[6] [1]);
	assign _0046_ = (\mchip.pc [1] ? _0045_ : _0044_);
	assign _0047_ = (\mchip.pc [2] ? _0046_ : _0043_);
	assign _0048_ = (\mchip.pc [0] ? \mchip.prog[9] [1] : \mchip.prog[8] [1]);
	assign _0049_ = (\mchip.pc [0] ? \mchip.prog[11] [1] : \mchip.prog[10] [1]);
	assign _0050_ = (\mchip.pc [1] ? _0049_ : _0048_);
	assign _0051_ = (\mchip.pc [0] ? \mchip.prog[13] [1] : \mchip.prog[12] [1]);
	assign _0052_ = (\mchip.pc [0] ? \mchip.prog[15] [1] : \mchip.prog[14] [1]);
	assign _0053_ = (\mchip.pc [1] ? _0052_ : _0051_);
	assign _0054_ = (\mchip.pc [2] ? _0053_ : _0050_);
	assign _0055_ = (\mchip.pc [3] ? _0054_ : _0047_);
	assign _0056_ = (\mchip.pc [0] ? \mchip.prog[1] [0] : \mchip.prog[0] [0]);
	assign _0057_ = (\mchip.pc [0] ? \mchip.prog[3] [0] : \mchip.prog[2] [0]);
	assign _0058_ = (\mchip.pc [1] ? _0057_ : _0056_);
	assign _0059_ = (\mchip.pc [0] ? \mchip.prog[5] [0] : \mchip.prog[4] [0]);
	assign _0060_ = (\mchip.pc [0] ? \mchip.prog[7] [0] : \mchip.prog[6] [0]);
	assign _0061_ = (\mchip.pc [1] ? _0060_ : _0059_);
	assign _0062_ = (\mchip.pc [2] ? _0061_ : _0058_);
	assign _0063_ = (\mchip.pc [0] ? \mchip.prog[9] [0] : \mchip.prog[8] [0]);
	assign _0064_ = (\mchip.pc [0] ? \mchip.prog[11] [0] : \mchip.prog[10] [0]);
	assign _0065_ = (\mchip.pc [1] ? _0064_ : _0063_);
	assign _0066_ = (\mchip.pc [0] ? \mchip.prog[13] [0] : \mchip.prog[12] [0]);
	assign _0067_ = (\mchip.pc [0] ? \mchip.prog[15] [0] : \mchip.prog[14] [0]);
	assign _0068_ = (\mchip.pc [1] ? _0067_ : _0066_);
	assign _0069_ = (\mchip.pc [2] ? _0068_ : _0065_);
	assign _0070_ = (\mchip.pc [3] ? _0069_ : _0062_);
	assign _0071_ = ~(_0070_ | _0055_);
	assign _0072_ = (\mchip.pc [0] ? \mchip.prog[1] [2] : \mchip.prog[0] [2]);
	assign _0073_ = (\mchip.pc [0] ? \mchip.prog[3] [2] : \mchip.prog[2] [2]);
	assign _0074_ = (\mchip.pc [1] ? _0073_ : _0072_);
	assign _0075_ = (\mchip.pc [0] ? \mchip.prog[5] [2] : \mchip.prog[4] [2]);
	assign _0076_ = (\mchip.pc [0] ? \mchip.prog[7] [2] : \mchip.prog[6] [2]);
	assign _0077_ = (\mchip.pc [1] ? _0076_ : _0075_);
	assign _0078_ = (\mchip.pc [2] ? _0077_ : _0074_);
	assign _0079_ = (\mchip.pc [0] ? \mchip.prog[9] [2] : \mchip.prog[8] [2]);
	assign _0080_ = (\mchip.pc [0] ? \mchip.prog[11] [2] : \mchip.prog[10] [2]);
	assign _0081_ = (\mchip.pc [1] ? _0080_ : _0079_);
	assign _0082_ = (\mchip.pc [0] ? \mchip.prog[13] [2] : \mchip.prog[12] [2]);
	assign _0083_ = (\mchip.pc [0] ? \mchip.prog[15] [2] : \mchip.prog[14] [2]);
	assign _0084_ = (\mchip.pc [1] ? _0083_ : _0082_);
	assign _0085_ = (\mchip.pc [2] ? _0084_ : _0081_);
	assign _0086_ = (\mchip.pc [3] ? _0085_ : _0078_);
	assign _0087_ = (\mchip.pc [0] ? \mchip.prog[1] [3] : \mchip.prog[0] [3]);
	assign _0088_ = (\mchip.pc [0] ? \mchip.prog[3] [3] : \mchip.prog[2] [3]);
	assign _0089_ = (\mchip.pc [1] ? _0088_ : _0087_);
	assign _0090_ = (\mchip.pc [0] ? \mchip.prog[5] [3] : \mchip.prog[4] [3]);
	assign _0091_ = (\mchip.pc [0] ? \mchip.prog[7] [3] : \mchip.prog[6] [3]);
	assign _0092_ = (\mchip.pc [1] ? _0091_ : _0090_);
	assign _0093_ = (\mchip.pc [2] ? _0092_ : _0089_);
	assign _0094_ = (\mchip.pc [0] ? \mchip.prog[9] [3] : \mchip.prog[8] [3]);
	assign _0095_ = (\mchip.pc [0] ? \mchip.prog[11] [3] : \mchip.prog[10] [3]);
	assign _0096_ = (\mchip.pc [1] ? _0095_ : _0094_);
	assign _0097_ = (\mchip.pc [0] ? \mchip.prog[13] [3] : \mchip.prog[12] [3]);
	assign _0098_ = (\mchip.pc [0] ? \mchip.prog[15] [3] : \mchip.prog[14] [3]);
	assign _0099_ = (\mchip.pc [1] ? _0098_ : _0097_);
	assign _0100_ = (\mchip.pc [2] ? _0099_ : _0096_);
	assign _0101_ = (\mchip.pc [3] ? _0100_ : _0093_);
	assign _0102_ = _0101_ & ~_0086_;
	assign _0103_ = _0102_ & _0071_;
	assign _0104_ = _0070_ & ~_0055_;
	assign _0105_ = _0104_ & _0102_;
	assign _0106_ = ~(_0105_ | _0103_);
	assign _0107_ = _0101_ | ~_0086_;
	assign _0108_ = _0104_ & ~_0107_;
	assign _0109_ = _0086_ & ~_0101_;
	assign _0110_ = _0070_ | ~_0055_;
	assign _0111_ = _0109_ & ~_0110_;
	assign _0112_ = _0111_ | _0108_;
	assign _0113_ = _0106_ & ~_0112_;
	assign _0114_ = _0071_ & ~_0107_;
	assign _0115_ = ~(_0070_ & _0055_);
	assign _0116_ = _0101_ | _0086_;
	assign _0117_ = ~(_0116_ | _0115_);
	assign _0118_ = _0117_ | _0114_;
	assign _0119_ = _0055_ & ~_0070_;
	assign _0120_ = _0119_ & ~_0116_;
	assign _0121_ = _0071_ & ~_0116_;
	assign _0122_ = _0121_ | _0120_;
	assign _0123_ = _0122_ | _0118_;
	assign _0124_ = _0113_ & ~_0123_;
	assign _0125_ = ~(_0101_ & _0086_);
	assign _0126_ = _0104_ & ~_0125_;
	assign _0127_ = _0119_ & ~_0125_;
	assign _0128_ = ~(_0127_ | _0126_);
	assign _0129_ = _0102_ & ~_0110_;
	assign _0130_ = _0102_ & ~_0115_;
	assign _0131_ = _0130_ | _0129_;
	assign _0132_ = _0125_ | _0115_;
	assign _0133_ = _0071_ & ~_0125_;
	assign _0134_ = _0133_ | ~_0132_;
	assign _0135_ = ~(_0134_ | _0131_);
	assign _0136_ = ~(_0135_ & _0128_);
	assign _0137_ = _0124_ & ~_0136_;
	assign _0000_ = _0037_ & ~_0137_;
	assign _0138_ = _0126_ | ~_0132_;
	assign _0139_ = _0138_ | _0127_;
	assign _0140_ = _0133_ | _0130_;
	assign _0141_ = _0129_ | _0105_;
	assign _0142_ = _0141_ | _0140_;
	assign _0143_ = _0142_ | _0139_;
	assign _0144_ = _0109_ & ~_0115_;
	assign _0145_ = _0144_ | _0103_;
	assign _0146_ = _0145_ | _0112_;
	assign _0147_ = _0146_ | _0123_;
	assign _0148_ = _0147_ | _0143_;
	assign _0149_ = _0148_ | ~_0037_;
	assign _0150_ = _0149_ | io_in[1];
	assign _0001_ = (_0150_ ? io_in[4] : \mchip.regval [0]);
	assign _0002_ = (_0150_ ? io_in[5] : \mchip.regval [1]);
	assign _0003_ = (_0150_ ? io_in[6] : \mchip.regval [2]);
	assign _0004_ = (_0150_ ? io_in[7] : \mchip.regval [3]);
	assign _0151_ = (\mchip.pc [0] ? \mchip.data[1] [0] : \mchip.data[0] [0]);
	assign _0152_ = (\mchip.pc [0] ? \mchip.data[3] [0] : \mchip.data[2] [0]);
	assign _0153_ = (\mchip.pc [1] ? _0152_ : _0151_);
	assign _0154_ = (\mchip.pc [0] ? \mchip.data[5] [0] : \mchip.data[4] [0]);
	assign _0155_ = (\mchip.pc [0] ? \mchip.data[7] [0] : \mchip.data[6] [0]);
	assign _0156_ = (\mchip.pc [1] ? _0155_ : _0154_);
	assign _0157_ = (\mchip.pc [2] ? _0156_ : _0153_);
	assign _0158_ = (\mchip.pc [0] ? \mchip.data[9] [0] : \mchip.data[8] [0]);
	assign _0159_ = (\mchip.pc [0] ? \mchip.data[11] [0] : \mchip.data[10] [0]);
	assign _0160_ = (\mchip.pc [1] ? _0159_ : _0158_);
	assign _0161_ = (\mchip.pc [0] ? \mchip.data[13] [0] : \mchip.data[12] [0]);
	assign _0162_ = (\mchip.pc [0] ? \mchip.data[15] [0] : \mchip.data[14] [0]);
	assign _0163_ = (\mchip.pc [1] ? _0162_ : _0161_);
	assign _0164_ = (\mchip.pc [2] ? _0163_ : _0160_);
	assign _0165_ = (\mchip.pc [3] ? _0164_ : _0157_);
	assign _0166_ = ~\mchip.regval [0];
	assign _0167_ = _0165_ & ~_0166_;
	assign _0168_ = _0166_ & ~_0165_;
	assign _0169_ = ~(_0168_ | _0167_);
	assign _0170_ = _0169_ & _0120_;
	assign _0171_ = _0169_ & _0114_;
	assign _0172_ = ~_0167_;
	assign _0173_ = _0117_ & ~_0172_;
	assign _0174_ = _0173_ | _0171_;
	assign _0175_ = (\mchip.pc [0] ? \mchip.data[1] [3] : \mchip.data[0] [3]);
	assign _0176_ = (\mchip.pc [0] ? \mchip.data[3] [3] : \mchip.data[2] [3]);
	assign _0177_ = (\mchip.pc [1] ? _0176_ : _0175_);
	assign _0178_ = (\mchip.pc [0] ? \mchip.data[5] [3] : \mchip.data[4] [3]);
	assign _0179_ = (\mchip.pc [0] ? \mchip.data[7] [3] : \mchip.data[6] [3]);
	assign _0180_ = (\mchip.pc [1] ? _0179_ : _0178_);
	assign _0181_ = (\mchip.pc [2] ? _0180_ : _0177_);
	assign _0182_ = (\mchip.pc [0] ? \mchip.data[9] [3] : \mchip.data[8] [3]);
	assign _0183_ = (\mchip.pc [0] ? \mchip.data[11] [3] : \mchip.data[10] [3]);
	assign _0184_ = (\mchip.pc [1] ? _0183_ : _0182_);
	assign _0185_ = (\mchip.pc [0] ? \mchip.data[13] [3] : \mchip.data[12] [3]);
	assign _0186_ = (\mchip.pc [0] ? \mchip.data[15] [3] : \mchip.data[14] [3]);
	assign _0187_ = (\mchip.pc [1] ? _0186_ : _0185_);
	assign _0188_ = (\mchip.pc [2] ? _0187_ : _0184_);
	assign _0189_ = (\mchip.pc [3] ? _0188_ : _0181_);
	assign _0190_ = _0189_ | _0166_;
	assign _0191_ = _0190_ | _0165_;
	assign _0192_ = (\mchip.pc [0] ? \mchip.data[1] [1] : \mchip.data[0] [1]);
	assign _0193_ = (\mchip.pc [0] ? \mchip.data[3] [1] : \mchip.data[2] [1]);
	assign _0194_ = (\mchip.pc [1] ? _0193_ : _0192_);
	assign _0195_ = (\mchip.pc [0] ? \mchip.data[5] [1] : \mchip.data[4] [1]);
	assign _0196_ = (\mchip.pc [0] ? \mchip.data[7] [1] : \mchip.data[6] [1]);
	assign _0197_ = (\mchip.pc [1] ? _0196_ : _0195_);
	assign _0198_ = (\mchip.pc [2] ? _0197_ : _0194_);
	assign _0199_ = (\mchip.pc [0] ? \mchip.data[9] [1] : \mchip.data[8] [1]);
	assign _0200_ = (\mchip.pc [0] ? \mchip.data[11] [1] : \mchip.data[10] [1]);
	assign _0201_ = (\mchip.pc [1] ? _0200_ : _0199_);
	assign _0202_ = (\mchip.pc [0] ? \mchip.data[13] [1] : \mchip.data[12] [1]);
	assign _0203_ = (\mchip.pc [0] ? \mchip.data[15] [1] : \mchip.data[14] [1]);
	assign _0204_ = (\mchip.pc [1] ? _0203_ : _0202_);
	assign _0205_ = (\mchip.pc [2] ? _0204_ : _0201_);
	assign _0206_ = (\mchip.pc [3] ? _0205_ : _0198_);
	assign _0207_ = _0206_ | _0191_;
	assign _0208_ = (\mchip.pc [0] ? \mchip.data[1] [2] : \mchip.data[0] [2]);
	assign _0209_ = (\mchip.pc [0] ? \mchip.data[3] [2] : \mchip.data[2] [2]);
	assign _0210_ = (\mchip.pc [1] ? _0209_ : _0208_);
	assign _0211_ = (\mchip.pc [0] ? \mchip.data[5] [2] : \mchip.data[4] [2]);
	assign _0212_ = (\mchip.pc [0] ? \mchip.data[7] [2] : \mchip.data[6] [2]);
	assign _0213_ = (\mchip.pc [1] ? _0212_ : _0211_);
	assign _0214_ = (\mchip.pc [2] ? _0213_ : _0210_);
	assign _0215_ = (\mchip.pc [0] ? \mchip.data[9] [2] : \mchip.data[8] [2]);
	assign _0216_ = (\mchip.pc [0] ? \mchip.data[11] [2] : \mchip.data[10] [2]);
	assign _0217_ = (\mchip.pc [1] ? _0216_ : _0215_);
	assign _0218_ = (\mchip.pc [0] ? \mchip.data[13] [2] : \mchip.data[12] [2]);
	assign _0219_ = (\mchip.pc [0] ? \mchip.data[15] [2] : \mchip.data[14] [2]);
	assign _0220_ = (\mchip.pc [1] ? _0219_ : _0218_);
	assign _0221_ = (\mchip.pc [2] ? _0220_ : _0217_);
	assign _0222_ = (\mchip.pc [3] ? _0221_ : _0214_);
	assign _0223_ = _0222_ | _0207_;
	assign _0224_ = ~(_0222_ | _0189_);
	assign _0225_ = ~_0224_;
	assign _0226_ = _0225_ | _0223_;
	assign _0227_ = _0108_ & ~_0226_;
	assign _0228_ = ~\mchip.regval [3];
	assign _0229_ = ~\mchip.regval [1];
	assign _0230_ = _0189_ | _0229_;
	assign _0231_ = (_0165_ ? _0230_ : _0190_);
	assign _0232_ = ~\mchip.regval [2];
	assign _0233_ = _0189_ | _0232_;
	assign _0234_ = _0189_ | _0228_;
	assign _0235_ = (_0165_ ? _0234_ : _0233_);
	assign _0236_ = (_0206_ ? _0235_ : _0231_);
	assign _0237_ = _0236_ | _0222_;
	assign _0238_ = (_0224_ ? _0237_ : _0228_);
	assign _0239_ = _0111_ & ~_0238_;
	assign _0240_ = _0239_ | _0227_;
	assign _0241_ = _0240_ | _0174_;
	assign _0242_ = _0241_ | _0170_;
	assign _0243_ = _0206_ | _0165_;
	assign _0244_ = _0224_ & ~_0243_;
	assign _0245_ = ~(\mchip.regval [1] | \mchip.regval [0]);
	assign _0246_ = \mchip.regval [3] | \mchip.regval [2];
	assign _0247_ = _0245_ & ~_0246_;
	assign _0248_ = _0247_ | _0244_;
	assign _0249_ = _0103_ & ~_0248_;
	assign _0250_ = ~_0247_;
	assign _0251_ = _0244_ & ~_0250_;
	assign _0252_ = _0105_ & ~_0251_;
	assign _0253_ = _0252_ | _0249_;
	assign _0254_ = _0232_ & ~_0222_;
	assign _0255_ = _0222_ & ~_0232_;
	assign _0256_ = _0255_ | _0254_;
	assign _0257_ = _0228_ & ~_0189_;
	assign _0258_ = ~(_0189_ & \mchip.regval [3]);
	assign _0259_ = _0257_ | ~_0258_;
	assign _0260_ = _0259_ & _0256_;
	assign _0261_ = ~(_0206_ & \mchip.regval [1]);
	assign _0262_ = _0229_ & ~_0206_;
	assign _0263_ = _0261_ & ~_0262_;
	assign _0264_ = _0263_ | _0169_;
	assign _0265_ = _0260_ & ~_0264_;
	assign _0266_ = (_0265_ ? _0129_ : _0130_);
	assign _0267_ = _0266_ | _0253_;
	assign _0268_ = _0133_ & ~_0172_;
	assign _0269_ = _0166_ & ~_0132_;
	assign _0270_ = _0269_ | _0268_;
	assign _0271_ = _0126_ & ~_0168_;
	assign _0272_ = _0127_ & ~_0250_;
	assign _0273_ = _0272_ | _0271_;
	assign _0274_ = _0273_ | _0270_;
	assign _0275_ = _0274_ | _0267_;
	assign _0276_ = _0275_ | _0242_;
	assign _0277_ = _0128_ & ~_0134_;
	assign _0278_ = _0131_ | ~_0106_;
	assign _0279_ = _0277_ & ~_0278_;
	assign _0280_ = _0118_ | _0112_;
	assign _0281_ = _0280_ | _0120_;
	assign _0282_ = _0279_ & ~_0281_;
	assign _0497_[0] = (_0282_ ? _0165_ : _0276_);
	assign _0283_ = _0263_ ^ _0172_;
	assign _0284_ = _0120_ & ~_0283_;
	assign _0285_ = _0165_ & ~\mchip.regval [0];
	assign _0286_ = ~(_0285_ ^ _0263_);
	assign _0287_ = _0114_ & ~_0286_;
	assign _0288_ = ~(_0165_ & \mchip.regval [1]);
	assign _0289_ = ~(_0206_ & \mchip.regval [0]);
	assign _0290_ = ~(_0289_ ^ _0288_);
	assign _0291_ = _0117_ & ~_0290_;
	assign _0292_ = _0291_ | _0287_;
	assign _0293_ = (_0165_ ? _0190_ : _0230_);
	assign _0294_ = _0293_ | _0206_;
	assign _0295_ = _0294_ | _0222_;
	assign _0296_ = _0295_ | _0225_;
	assign _0297_ = _0108_ & ~_0296_;
	assign _0298_ = (_0165_ ? _0233_ : _0230_);
	assign _0299_ = _0234_ | _0165_;
	assign _0300_ = (_0206_ ? _0299_ : _0298_);
	assign _0301_ = _0300_ | _0222_;
	assign _0302_ = _0301_ | _0225_;
	assign _0303_ = _0111_ & ~_0302_;
	assign _0304_ = _0303_ | _0297_;
	assign _0305_ = _0304_ | _0292_;
	assign _0306_ = _0305_ | _0284_;
	assign _0307_ = _0133_ & ~_0261_;
	assign _0308_ = _0229_ & ~_0132_;
	assign _0309_ = _0308_ | _0307_;
	assign _0310_ = _0126_ & ~_0262_;
	assign _0311_ = _0310_ | _0309_;
	assign _0312_ = _0311_ | _0306_;
	assign _0497_[1] = (_0282_ ? _0206_ : _0312_);
	assign _0313_ = _0206_ & ~_0229_;
	assign _0314_ = _0263_ & ~_0172_;
	assign _0315_ = _0314_ | _0313_;
	assign _0316_ = _0222_ ^ _0232_;
	assign _0317_ = _0316_ ^ _0315_;
	assign _0318_ = _0120_ & ~_0317_;
	assign _0319_ = _0285_ | _0263_;
	assign _0320_ = \mchip.regval [1] & ~_0206_;
	assign _0321_ = _0319_ & ~_0320_;
	assign _0322_ = _0321_ ^ _0256_;
	assign _0323_ = _0114_ & ~_0322_;
	assign _0324_ = ~(_0289_ | _0288_);
	assign _0325_ = _0165_ & ~_0232_;
	assign _0326_ = ~(_0222_ & \mchip.regval [0]);
	assign _0327_ = _0326_ ^ _0313_;
	assign _0328_ = _0327_ ^ _0325_;
	assign _0329_ = _0328_ ^ _0324_;
	assign _0330_ = _0117_ & ~_0329_;
	assign _0331_ = _0330_ | _0323_;
	assign _0332_ = (_0165_ ? _0230_ : _0233_);
	assign _0333_ = (_0206_ ? _0191_ : _0332_);
	assign _0334_ = _0333_ | _0222_;
	assign _0335_ = _0334_ | _0225_;
	assign _0336_ = _0108_ & ~_0335_;
	assign _0337_ = _0235_ | _0206_;
	assign _0338_ = _0337_ | _0222_;
	assign _0339_ = _0338_ | _0225_;
	assign _0340_ = _0111_ & ~_0339_;
	assign _0341_ = _0340_ | _0336_;
	assign _0342_ = _0341_ | _0331_;
	assign _0343_ = _0342_ | _0318_;
	assign _0344_ = _0255_ & _0133_;
	assign _0345_ = _0232_ & ~_0132_;
	assign _0346_ = _0345_ | _0344_;
	assign _0347_ = _0126_ & ~_0254_;
	assign _0348_ = _0347_ | _0346_;
	assign _0349_ = _0348_ | _0343_;
	assign _0497_[2] = (_0282_ ? _0222_ : _0349_);
	assign _0350_ = _0315_ & ~_0316_;
	assign _0351_ = _0350_ | _0255_;
	assign _0352_ = _0189_ ^ _0228_;
	assign _0353_ = _0352_ ^ _0351_;
	assign _0354_ = _0120_ & ~_0353_;
	assign _0355_ = _0222_ | _0232_;
	assign _0356_ = _0256_ & ~_0321_;
	assign _0357_ = _0355_ & ~_0356_;
	assign _0358_ = _0357_ ^ _0259_;
	assign _0359_ = _0114_ & ~_0358_;
	assign _0360_ = _0328_ | ~_0324_;
	assign _0361_ = _0325_ & ~_0327_;
	assign _0362_ = _0165_ & ~_0228_;
	assign _0363_ = _0313_ & ~_0326_;
	assign _0364_ = _0206_ & ~_0232_;
	assign _0365_ = _0222_ & ~_0229_;
	assign _0366_ = _0189_ & ~_0166_;
	assign _0367_ = _0366_ ^ _0365_;
	assign _0368_ = _0367_ ^ _0364_;
	assign _0369_ = _0368_ ^ _0363_;
	assign _0370_ = _0369_ ^ _0362_;
	assign _0371_ = _0370_ ^ _0361_;
	assign _0372_ = _0371_ ^ _0360_;
	assign _0373_ = _0117_ & ~_0372_;
	assign _0374_ = _0373_ | _0359_;
	assign _0375_ = (_0165_ ? _0233_ : _0234_);
	assign _0376_ = (_0206_ ? _0293_ : _0375_);
	assign _0377_ = _0376_ | _0222_;
	assign _0378_ = (_0224_ ? _0377_ : _0166_);
	assign _0379_ = _0108_ & ~_0378_;
	assign _0380_ = _0299_ | _0206_;
	assign _0381_ = _0380_ | _0222_;
	assign _0382_ = _0381_ | _0225_;
	assign _0383_ = _0111_ & ~_0382_;
	assign _0384_ = _0383_ | _0379_;
	assign _0385_ = _0384_ | _0374_;
	assign _0386_ = _0385_ | _0354_;
	assign _0387_ = _0133_ & ~_0258_;
	assign _0388_ = _0228_ & ~_0132_;
	assign _0389_ = _0388_ | _0387_;
	assign _0390_ = _0126_ & ~_0257_;
	assign _0391_ = _0390_ | _0389_;
	assign _0392_ = _0391_ | _0386_;
	assign _0497_[3] = (_0282_ ? _0189_ : _0392_);
	assign _0393_ = ~\mchip.pc [0];
	assign _0394_ = io_in[3] & ~io_in[2];
	assign _0395_ = _0394_ & io_in[4];
	assign _0396_ = ~_0165_;
	assign _0397_ = (\mchip.lastdata3  ? _0396_ : \mchip.pc [0]);
	assign _0398_ = _0111_ | _0103_;
	assign _0399_ = _0117_ | _0108_;
	assign _0400_ = _0399_ | _0398_;
	assign _0401_ = _0120_ | _0114_;
	assign _0402_ = _0104_ & ~_0116_;
	assign _0403_ = _0402_ | _0121_;
	assign _0404_ = _0403_ | _0401_;
	assign _0405_ = _0404_ | _0400_;
	assign _0406_ = _0405_ | _0143_;
	assign _0407_ = (_0406_ ? \mchip.pc [0] : _0397_);
	assign _0408_ = _0037_ & ~_0407_;
	assign _0409_ = _0408_ | _0395_;
	assign _0410_ = ~(_0394_ | _0037_);
	assign _0496_[0] = (_0410_ ? _0393_ : _0409_);
	assign _0411_ = \mchip.pc [0] | ~\mchip.pc [1];
	assign _0412_ = \mchip.pc [1] | ~\mchip.pc [0];
	assign _0413_ = _0412_ & _0411_;
	assign _0414_ = ~_0413_;
	assign _0415_ = _0394_ & io_in[5];
	assign _0416_ = ~_0206_;
	assign _0417_ = (\mchip.lastdata3  ? _0416_ : _0413_);
	assign _0418_ = (_0406_ ? _0413_ : _0417_);
	assign _0419_ = _0037_ & ~_0418_;
	assign _0420_ = _0419_ | _0415_;
	assign _0496_[1] = (_0410_ ? _0414_ : _0420_);
	assign _0421_ = \mchip.pc [0] & \mchip.pc [1];
	assign _0422_ = _0421_ ^ \mchip.pc [2];
	assign _0423_ = _0394_ & io_in[6];
	assign _0424_ = (\mchip.lastdata3  ? _0222_ : _0422_);
	assign _0425_ = (_0406_ ? _0422_ : _0424_);
	assign _0426_ = _0425_ & _0037_;
	assign _0427_ = _0426_ | _0423_;
	assign _0496_[2] = (_0410_ ? _0422_ : _0427_);
	assign _0428_ = _0421_ & ~_0039_;
	assign _0429_ = _0428_ ^ \mchip.pc [3];
	assign _0430_ = _0394_ & io_in[7];
	assign _0431_ = (\mchip.lastdata3  ? _0189_ : _0429_);
	assign _0432_ = (_0406_ ? _0429_ : _0431_);
	assign _0433_ = _0432_ & _0037_;
	assign _0434_ = _0433_ | _0430_;
	assign _0496_[3] = (_0410_ ? _0429_ : _0434_);
	assign _0435_ = ~io_in[1];
	assign _0436_ = io_in[3] | ~io_in[2];
	assign _0437_ = _0435_ & ~_0436_;
	assign _0438_ = _0437_ | ~_0150_;
	assign _0439_ = ~_0189_;
	assign _0440_ = (_0150_ ? _0038_ : _0439_);
	assign _0441_ = ~_0222_;
	assign _0442_ = (_0150_ ? _0039_ : _0441_);
	assign _0443_ = _0442_ | _0440_;
	assign _0444_ = (_0150_ ? \mchip.pc [1] : _0206_);
	assign _0445_ = (_0150_ ? _0393_ : _0396_);
	assign _0446_ = _0445_ | _0444_;
	assign _0447_ = _0446_ | _0443_;
	assign _0009_ = _0438_ & ~_0447_;
	assign _0448_ = (_0150_ ? _0040_ : _0416_);
	assign _0449_ = (_0150_ ? \mchip.pc [0] : _0165_);
	assign _0450_ = _0449_ | _0448_;
	assign _0451_ = _0450_ | _0443_;
	assign _0010_ = _0438_ & ~_0451_;
	assign _0452_ = io_in[2] | io_in[3];
	assign _0453_ = _0435_ & ~_0452_;
	assign _0454_ = ~(\mchip.pc [2] & \mchip.pc [3]);
	assign _0455_ = _0454_ | _0412_;
	assign _0025_ = _0453_ & ~_0455_;
	assign _0456_ = _0448_ | _0445_;
	assign _0457_ = _0456_ | _0443_;
	assign _0011_ = _0438_ & ~_0457_;
	assign _0458_ = _0454_ | _0411_;
	assign _0026_ = _0453_ & ~_0458_;
	assign _0459_ = \mchip.pc [2] | \mchip.pc [3];
	assign _0460_ = \mchip.pc [0] | \mchip.pc [1];
	assign _0461_ = _0460_ | _0459_;
	assign _0021_ = _0453_ & ~_0461_;
	assign _0462_ = _0454_ | ~_0421_;
	assign _0027_ = _0453_ & ~_0462_;
	assign _0463_ = _0459_ | _0412_;
	assign _0028_ = _0453_ & ~_0463_;
	assign _0464_ = _0459_ | _0411_;
	assign _0029_ = _0453_ & ~_0464_;
	assign _0465_ = _0459_ | ~_0421_;
	assign _0030_ = _0453_ & ~_0465_;
	assign _0466_ = \mchip.pc [3] | ~\mchip.pc [2];
	assign _0467_ = _0466_ | _0460_;
	assign _0031_ = _0453_ & ~_0467_;
	assign _0468_ = _0466_ | _0412_;
	assign _0032_ = _0453_ & ~_0468_;
	assign _0469_ = _0466_ | _0411_;
	assign _0033_ = _0453_ & ~_0469_;
	assign _0470_ = _0466_ | ~_0421_;
	assign _0034_ = _0453_ & ~_0470_;
	assign _0471_ = \mchip.pc [2] | ~\mchip.pc [3];
	assign _0472_ = _0471_ | _0460_;
	assign _0035_ = _0453_ & ~_0472_;
	assign _0473_ = _0471_ | _0412_;
	assign _0036_ = _0453_ & ~_0473_;
	assign _0474_ = _0471_ | _0411_;
	assign _0022_ = _0453_ & ~_0474_;
	assign _0475_ = _0471_ | ~_0421_;
	assign _0023_ = _0453_ & ~_0475_;
	assign _0476_ = _0460_ | _0454_;
	assign _0024_ = _0453_ & ~_0476_;
	assign _0477_ = (_0150_ ? \mchip.pc [2] : _0222_);
	assign _0478_ = _0477_ | _0440_;
	assign _0479_ = _0478_ | _0456_;
	assign _0007_ = _0438_ & ~_0479_;
	assign _0480_ = _0478_ | _0450_;
	assign _0006_ = _0438_ & ~_0480_;
	assign _0481_ = _0478_ | _0446_;
	assign _0020_ = _0438_ & ~_0481_;
	assign _0482_ = _0449_ | _0444_;
	assign _0483_ = _0482_ | _0478_;
	assign _0019_ = _0438_ & ~_0483_;
	assign _0484_ = (_0150_ ? \mchip.pc [3] : _0189_);
	assign _0485_ = _0484_ | _0477_;
	assign _0486_ = _0485_ | _0482_;
	assign _0005_ = _0438_ & ~_0486_;
	assign _0487_ = _0484_ | _0442_;
	assign _0488_ = _0487_ | _0456_;
	assign _0018_ = _0438_ & ~_0488_;
	assign _0489_ = _0487_ | _0450_;
	assign _0017_ = _0438_ & ~_0489_;
	assign _0490_ = _0487_ | _0446_;
	assign _0016_ = _0438_ & ~_0490_;
	assign _0491_ = _0487_ | _0482_;
	assign _0015_ = _0438_ & ~_0491_;
	assign _0492_ = _0482_ | _0443_;
	assign _0008_ = _0438_ & ~_0492_;
	assign _0493_ = _0485_ | _0446_;
	assign _0012_ = _0438_ & ~_0493_;
	assign _0494_ = _0485_ | _0456_;
	assign _0014_ = _0438_ & ~_0494_;
	assign _0495_ = _0485_ | _0450_;
	assign _0013_ = _0438_ & ~_0495_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[0] [0] <= 1'h0;
		else if (_0021_)
			\mchip.prog[0] [0] <= io_in[4];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[0] [1] <= 1'h0;
		else if (_0021_)
			\mchip.prog[0] [1] <= io_in[5];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[0] [2] <= 1'h0;
		else if (_0021_)
			\mchip.prog[0] [2] <= io_in[6];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[0] [3] <= 1'h0;
		else if (_0021_)
			\mchip.prog[0] [3] <= io_in[7];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[1] [0] <= 1'h0;
		else if (_0028_)
			\mchip.prog[1] [0] <= io_in[4];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[1] [1] <= 1'h0;
		else if (_0028_)
			\mchip.prog[1] [1] <= io_in[5];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[1] [2] <= 1'h0;
		else if (_0028_)
			\mchip.prog[1] [2] <= io_in[6];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[1] [3] <= 1'h0;
		else if (_0028_)
			\mchip.prog[1] [3] <= io_in[7];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[2] [0] <= 1'h0;
		else if (_0029_)
			\mchip.prog[2] [0] <= io_in[4];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[2] [1] <= 1'h0;
		else if (_0029_)
			\mchip.prog[2] [1] <= io_in[5];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[2] [2] <= 1'h0;
		else if (_0029_)
			\mchip.prog[2] [2] <= io_in[6];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[2] [3] <= 1'h0;
		else if (_0029_)
			\mchip.prog[2] [3] <= io_in[7];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[3] [0] <= 1'h0;
		else if (_0030_)
			\mchip.prog[3] [0] <= io_in[4];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[3] [1] <= 1'h0;
		else if (_0030_)
			\mchip.prog[3] [1] <= io_in[5];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[3] [2] <= 1'h0;
		else if (_0030_)
			\mchip.prog[3] [2] <= io_in[6];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[3] [3] <= 1'h0;
		else if (_0030_)
			\mchip.prog[3] [3] <= io_in[7];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[4] [0] <= 1'h0;
		else if (_0031_)
			\mchip.prog[4] [0] <= io_in[4];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[4] [1] <= 1'h0;
		else if (_0031_)
			\mchip.prog[4] [1] <= io_in[5];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[4] [2] <= 1'h0;
		else if (_0031_)
			\mchip.prog[4] [2] <= io_in[6];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[4] [3] <= 1'h0;
		else if (_0031_)
			\mchip.prog[4] [3] <= io_in[7];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[5] [0] <= 1'h0;
		else if (_0032_)
			\mchip.prog[5] [0] <= io_in[4];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[5] [1] <= 1'h0;
		else if (_0032_)
			\mchip.prog[5] [1] <= io_in[5];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[5] [2] <= 1'h0;
		else if (_0032_)
			\mchip.prog[5] [2] <= io_in[6];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[5] [3] <= 1'h0;
		else if (_0032_)
			\mchip.prog[5] [3] <= io_in[7];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[6] [0] <= 1'h0;
		else if (_0033_)
			\mchip.prog[6] [0] <= io_in[4];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[6] [1] <= 1'h0;
		else if (_0033_)
			\mchip.prog[6] [1] <= io_in[5];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[6] [2] <= 1'h0;
		else if (_0033_)
			\mchip.prog[6] [2] <= io_in[6];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[6] [3] <= 1'h0;
		else if (_0033_)
			\mchip.prog[6] [3] <= io_in[7];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[7] [0] <= 1'h0;
		else if (_0034_)
			\mchip.prog[7] [0] <= io_in[4];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[7] [1] <= 1'h0;
		else if (_0034_)
			\mchip.prog[7] [1] <= io_in[5];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[7] [2] <= 1'h0;
		else if (_0034_)
			\mchip.prog[7] [2] <= io_in[6];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[7] [3] <= 1'h0;
		else if (_0034_)
			\mchip.prog[7] [3] <= io_in[7];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[8] [0] <= 1'h0;
		else if (_0035_)
			\mchip.prog[8] [0] <= io_in[4];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[8] [1] <= 1'h0;
		else if (_0035_)
			\mchip.prog[8] [1] <= io_in[5];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[8] [2] <= 1'h0;
		else if (_0035_)
			\mchip.prog[8] [2] <= io_in[6];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[8] [3] <= 1'h0;
		else if (_0035_)
			\mchip.prog[8] [3] <= io_in[7];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[9] [0] <= 1'h0;
		else if (_0036_)
			\mchip.prog[9] [0] <= io_in[4];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[9] [1] <= 1'h0;
		else if (_0036_)
			\mchip.prog[9] [1] <= io_in[5];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[9] [2] <= 1'h0;
		else if (_0036_)
			\mchip.prog[9] [2] <= io_in[6];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[9] [3] <= 1'h0;
		else if (_0036_)
			\mchip.prog[9] [3] <= io_in[7];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[10] [0] <= 1'h0;
		else if (_0022_)
			\mchip.prog[10] [0] <= io_in[4];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[10] [1] <= 1'h0;
		else if (_0022_)
			\mchip.prog[10] [1] <= io_in[5];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[10] [2] <= 1'h0;
		else if (_0022_)
			\mchip.prog[10] [2] <= io_in[6];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[10] [3] <= 1'h0;
		else if (_0022_)
			\mchip.prog[10] [3] <= io_in[7];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[11] [0] <= 1'h0;
		else if (_0023_)
			\mchip.prog[11] [0] <= io_in[4];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[11] [1] <= 1'h0;
		else if (_0023_)
			\mchip.prog[11] [1] <= io_in[5];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[11] [2] <= 1'h0;
		else if (_0023_)
			\mchip.prog[11] [2] <= io_in[6];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[11] [3] <= 1'h0;
		else if (_0023_)
			\mchip.prog[11] [3] <= io_in[7];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[12] [0] <= 1'h0;
		else if (_0024_)
			\mchip.prog[12] [0] <= io_in[4];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[12] [1] <= 1'h0;
		else if (_0024_)
			\mchip.prog[12] [1] <= io_in[5];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[12] [2] <= 1'h0;
		else if (_0024_)
			\mchip.prog[12] [2] <= io_in[6];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[12] [3] <= 1'h0;
		else if (_0024_)
			\mchip.prog[12] [3] <= io_in[7];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[13] [0] <= 1'h0;
		else if (_0025_)
			\mchip.prog[13] [0] <= io_in[4];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[13] [1] <= 1'h0;
		else if (_0025_)
			\mchip.prog[13] [1] <= io_in[5];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[13] [2] <= 1'h0;
		else if (_0025_)
			\mchip.prog[13] [2] <= io_in[6];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[13] [3] <= 1'h0;
		else if (_0025_)
			\mchip.prog[13] [3] <= io_in[7];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[14] [0] <= 1'h0;
		else if (_0026_)
			\mchip.prog[14] [0] <= io_in[4];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[14] [1] <= 1'h0;
		else if (_0026_)
			\mchip.prog[14] [1] <= io_in[5];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[14] [2] <= 1'h0;
		else if (_0026_)
			\mchip.prog[14] [2] <= io_in[6];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[14] [3] <= 1'h0;
		else if (_0026_)
			\mchip.prog[14] [3] <= io_in[7];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[15] [0] <= 1'h0;
		else if (_0027_)
			\mchip.prog[15] [0] <= io_in[4];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[15] [1] <= 1'h0;
		else if (_0027_)
			\mchip.prog[15] [1] <= io_in[5];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[15] [2] <= 1'h0;
		else if (_0027_)
			\mchip.prog[15] [2] <= io_in[6];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.prog[15] [3] <= 1'h0;
		else if (_0027_)
			\mchip.prog[15] [3] <= io_in[7];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.pc [0] <= 1'h0;
		else
			\mchip.pc [0] <= _0496_[0];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.pc [1] <= 1'h0;
		else
			\mchip.pc [1] <= _0496_[1];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.pc [2] <= 1'h0;
		else
			\mchip.pc [2] <= _0496_[2];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.pc [3] <= 1'h0;
		else
			\mchip.pc [3] <= _0496_[3];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[4] [0] <= 1'h0;
		else if (_0015_)
			\mchip.data[4] [0] <= _0001_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[4] [1] <= 1'h0;
		else if (_0015_)
			\mchip.data[4] [1] <= _0002_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[4] [2] <= 1'h0;
		else if (_0015_)
			\mchip.data[4] [2] <= _0003_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[4] [3] <= 1'h0;
		else if (_0015_)
			\mchip.data[4] [3] <= _0004_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[5] [0] <= 1'h0;
		else if (_0016_)
			\mchip.data[5] [0] <= _0001_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[5] [1] <= 1'h0;
		else if (_0016_)
			\mchip.data[5] [1] <= _0002_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[5] [2] <= 1'h0;
		else if (_0016_)
			\mchip.data[5] [2] <= _0003_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[5] [3] <= 1'h0;
		else if (_0016_)
			\mchip.data[5] [3] <= _0004_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.lastdata3  <= 1'h0;
		else
			\mchip.lastdata3  <= io_in[7];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[1] [0] <= 1'h0;
		else if (_0012_)
			\mchip.data[1] [0] <= _0001_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[1] [1] <= 1'h0;
		else if (_0012_)
			\mchip.data[1] [1] <= _0002_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[1] [2] <= 1'h0;
		else if (_0012_)
			\mchip.data[1] [2] <= _0003_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[1] [3] <= 1'h0;
		else if (_0012_)
			\mchip.data[1] [3] <= _0004_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[2] [0] <= 1'h0;
		else if (_0013_)
			\mchip.data[2] [0] <= _0001_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[2] [1] <= 1'h0;
		else if (_0013_)
			\mchip.data[2] [1] <= _0002_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[2] [2] <= 1'h0;
		else if (_0013_)
			\mchip.data[2] [2] <= _0003_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[2] [3] <= 1'h0;
		else if (_0013_)
			\mchip.data[2] [3] <= _0004_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[3] [0] <= 1'h0;
		else if (_0014_)
			\mchip.data[3] [0] <= _0001_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[3] [1] <= 1'h0;
		else if (_0014_)
			\mchip.data[3] [1] <= _0002_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[3] [2] <= 1'h0;
		else if (_0014_)
			\mchip.data[3] [2] <= _0003_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[3] [3] <= 1'h0;
		else if (_0014_)
			\mchip.data[3] [3] <= _0004_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[12] [0] <= 1'h0;
		else if (_0008_)
			\mchip.data[12] [0] <= _0001_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[12] [1] <= 1'h0;
		else if (_0008_)
			\mchip.data[12] [1] <= _0002_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[12] [2] <= 1'h0;
		else if (_0008_)
			\mchip.data[12] [2] <= _0003_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[12] [3] <= 1'h0;
		else if (_0008_)
			\mchip.data[12] [3] <= _0004_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[15] [0] <= 1'h0;
		else if (_0011_)
			\mchip.data[15] [0] <= _0001_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[15] [1] <= 1'h0;
		else if (_0011_)
			\mchip.data[15] [1] <= _0002_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[15] [2] <= 1'h0;
		else if (_0011_)
			\mchip.data[15] [2] <= _0003_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[15] [3] <= 1'h0;
		else if (_0011_)
			\mchip.data[15] [3] <= _0004_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[14] [0] <= 1'h0;
		else if (_0010_)
			\mchip.data[14] [0] <= _0001_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[14] [1] <= 1'h0;
		else if (_0010_)
			\mchip.data[14] [1] <= _0002_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[14] [2] <= 1'h0;
		else if (_0010_)
			\mchip.data[14] [2] <= _0003_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[14] [3] <= 1'h0;
		else if (_0010_)
			\mchip.data[14] [3] <= _0004_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.regval [0] <= 1'h0;
		else if (_0000_)
			\mchip.regval [0] <= _0497_[0];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.regval [1] <= 1'h0;
		else if (_0000_)
			\mchip.regval [1] <= _0497_[1];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.regval [2] <= 1'h0;
		else if (_0000_)
			\mchip.regval [2] <= _0497_[2];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.regval [3] <= 1'h0;
		else if (_0000_)
			\mchip.regval [3] <= _0497_[3];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[10] [0] <= 1'h0;
		else if (_0006_)
			\mchip.data[10] [0] <= _0001_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[10] [1] <= 1'h0;
		else if (_0006_)
			\mchip.data[10] [1] <= _0002_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[10] [2] <= 1'h0;
		else if (_0006_)
			\mchip.data[10] [2] <= _0003_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[10] [3] <= 1'h0;
		else if (_0006_)
			\mchip.data[10] [3] <= _0004_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[8] [0] <= 1'h0;
		else if (_0019_)
			\mchip.data[8] [0] <= _0001_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[8] [1] <= 1'h0;
		else if (_0019_)
			\mchip.data[8] [1] <= _0002_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[8] [2] <= 1'h0;
		else if (_0019_)
			\mchip.data[8] [2] <= _0003_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[8] [3] <= 1'h0;
		else if (_0019_)
			\mchip.data[8] [3] <= _0004_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[7] [0] <= 1'h0;
		else if (_0018_)
			\mchip.data[7] [0] <= _0001_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[7] [1] <= 1'h0;
		else if (_0018_)
			\mchip.data[7] [1] <= _0002_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[7] [2] <= 1'h0;
		else if (_0018_)
			\mchip.data[7] [2] <= _0003_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[7] [3] <= 1'h0;
		else if (_0018_)
			\mchip.data[7] [3] <= _0004_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[0] [0] <= 1'h0;
		else if (_0005_)
			\mchip.data[0] [0] <= _0001_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[0] [1] <= 1'h0;
		else if (_0005_)
			\mchip.data[0] [1] <= _0002_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[0] [2] <= 1'h0;
		else if (_0005_)
			\mchip.data[0] [2] <= _0003_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[0] [3] <= 1'h0;
		else if (_0005_)
			\mchip.data[0] [3] <= _0004_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[6] [0] <= 1'h0;
		else if (_0017_)
			\mchip.data[6] [0] <= _0001_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[6] [1] <= 1'h0;
		else if (_0017_)
			\mchip.data[6] [1] <= _0002_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[6] [2] <= 1'h0;
		else if (_0017_)
			\mchip.data[6] [2] <= _0003_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[6] [3] <= 1'h0;
		else if (_0017_)
			\mchip.data[6] [3] <= _0004_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[9] [0] <= 1'h0;
		else if (_0020_)
			\mchip.data[9] [0] <= _0001_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[9] [1] <= 1'h0;
		else if (_0020_)
			\mchip.data[9] [1] <= _0002_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[9] [2] <= 1'h0;
		else if (_0020_)
			\mchip.data[9] [2] <= _0003_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[9] [3] <= 1'h0;
		else if (_0020_)
			\mchip.data[9] [3] <= _0004_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[11] [0] <= 1'h0;
		else if (_0007_)
			\mchip.data[11] [0] <= _0001_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[11] [1] <= 1'h0;
		else if (_0007_)
			\mchip.data[11] [1] <= _0002_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[11] [2] <= 1'h0;
		else if (_0007_)
			\mchip.data[11] [2] <= _0003_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[11] [3] <= 1'h0;
		else if (_0007_)
			\mchip.data[11] [3] <= _0004_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[13] [0] <= 1'h0;
		else if (_0009_)
			\mchip.data[13] [0] <= _0001_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[13] [1] <= 1'h0;
		else if (_0009_)
			\mchip.data[13] [1] <= _0002_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[13] [2] <= 1'h0;
		else if (_0009_)
			\mchip.data[13] [2] <= _0003_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.data[13] [3] <= 1'h0;
		else if (_0009_)
			\mchip.data[13] [3] <= _0004_;
	assign io_out = {6'h00, \mchip.regval , \mchip.pc };
	assign \mchip.clock  = io_in[0];
	assign \mchip.inputdata  = io_in[7:4];
	assign \mchip.instruction  = io_in[3:2];
	assign \mchip.io_in  = io_in[7:0];
	assign \mchip.io_out  = {\mchip.regval , \mchip.pc };
	assign \mchip.reset  = io_in[1];
endmodule
module d33_mgee3_adder (
	io_in,
	io_out
);
	wire _00_;
	wire _01_;
	wire _02_;
	wire _03_;
	wire _04_;
	wire _05_;
	wire _06_;
	wire _07_;
	input wire [13:0] io_in;
	output wire [13:0] io_out;
	wire \mchip.gate10.a ;
	wire \mchip.gate10.b ;
	wire \mchip.gate12.a ;
	wire \mchip.gate12.b ;
	wire \mchip.gate13.out ;
	wire \mchip.gate15.a ;
	wire \mchip.gate15.b ;
	wire \mchip.gate16.out ;
	wire \mchip.gate17.a ;
	wire \mchip.gate17.b ;
	wire \mchip.gate18.a ;
	wire \mchip.gate18.b ;
	wire \mchip.gate18.out ;
	wire \mchip.gate7.a ;
	wire \mchip.gate7.b ;
	wire \mchip.gate8.out ;
	wire [7:0] \mchip.io_in ;
	wire [7:0] \mchip.io_out ;
	wire \mchip.net1 ;
	wire \mchip.net10 ;
	wire \mchip.net11 ;
	wire \mchip.net12 ;
	wire \mchip.net14 ;
	wire \mchip.net2 ;
	wire \mchip.net22 ;
	wire \mchip.net3 ;
	wire \mchip.net4 ;
	wire \mchip.net5 ;
	wire \mchip.net6 ;
	wire \mchip.net7 ;
	wire \mchip.net8 ;
	wire \mchip.net9 ;
	assign \mchip.gate18.out  = io_in[0] ^ io_in[3];
	assign _00_ = io_in[2] & io_in[5];
	assign _01_ = ~(io_in[0] & io_in[3]);
	assign _02_ = ~(io_in[1] ^ io_in[4]);
	assign _03_ = ~(_02_ | _01_);
	assign _04_ = io_in[1] & io_in[4];
	assign _05_ = _04_ | _03_;
	assign _06_ = io_in[2] ^ io_in[5];
	assign _07_ = _06_ & _05_;
	assign \mchip.gate16.out  = _07_ | _00_;
	assign \mchip.gate13.out  = _06_ ^ _05_;
	assign \mchip.gate8.out  = _02_ ^ _01_;
	assign io_out = {10'h000, \mchip.gate16.out , \mchip.gate13.out , \mchip.gate8.out , \mchip.gate18.out };
	assign \mchip.gate10.a  = io_in[1];
	assign \mchip.gate10.b  = io_in[4];
	assign \mchip.gate12.a  = io_in[2];
	assign \mchip.gate12.b  = io_in[5];
	assign \mchip.gate15.a  = io_in[2];
	assign \mchip.gate15.b  = io_in[5];
	assign \mchip.gate17.a  = io_in[0];
	assign \mchip.gate17.b  = io_in[3];
	assign \mchip.gate18.a  = io_in[0];
	assign \mchip.gate18.b  = io_in[3];
	assign \mchip.gate7.a  = io_in[1];
	assign \mchip.gate7.b  = io_in[4];
	assign \mchip.io_in  = io_in[7:0];
	assign \mchip.io_out  = {4'h0, \mchip.gate16.out , \mchip.gate13.out , \mchip.gate8.out , \mchip.gate18.out };
	assign \mchip.net1  = \mchip.gate18.out ;
	assign \mchip.net10  = io_in[5];
	assign \mchip.net11  = 1'h0;
	assign \mchip.net12  = 1'h1;
	assign \mchip.net14  = 1'h0;
	assign \mchip.net2  = \mchip.gate8.out ;
	assign \mchip.net22  = 1'h0;
	assign \mchip.net3  = \mchip.gate13.out ;
	assign \mchip.net4  = \mchip.gate16.out ;
	assign \mchip.net5  = io_in[0];
	assign \mchip.net6  = io_in[1];
	assign \mchip.net7  = io_in[2];
	assign \mchip.net8  = io_in[3];
	assign \mchip.net9  = io_in[4];
endmodule
module d34_hgrodin_collatz (
	io_in,
	io_out
);
	wire _00_;
	wire _01_;
	wire _02_;
	wire _03_;
	wire _04_;
	wire _05_;
	wire _06_;
	wire _07_;
	wire _08_;
	wire _09_;
	wire _10_;
	wire _11_;
	wire _12_;
	input wire [13:0] io_in;
	output wire [13:0] io_out;
	wire [3:0] \mchip.c.b ;
	wire [3:0] \mchip.c.inst2.in1 ;
	wire [3:0] \mchip.c.inst2.in2 ;
	wire [3:0] \mchip.c.inst2.out ;
	wire [3:0] \mchip.c.inst2.rem ;
	wire [3:0] \mchip.c.inst3.in1 ;
	wire [3:0] \mchip.c.inst3.in2 ;
	wire [3:0] \mchip.c.inst3.rem ;
	wire [3:0] \mchip.c.n ;
	wire [3:0] \mchip.c.out ;
	wire [3:0] \mchip.c.out_even ;
	wire [3:0] \mchip.c.tmp ;
	wire [3:0] \mchip.c.tmp2 ;
	wire [7:0] \mchip.io_in ;
	wire [7:0] \mchip.io_out ;
	assign io_out[0] = io_in[1] & ~io_in[0];
	assign _00_ = io_in[1] | ~io_in[0];
	assign _01_ = ~(io_in[2] ^ io_in[1]);
	assign _02_ = io_in[0] & io_in[1];
	assign _03_ = _02_ ^ _01_;
	assign _04_ = _03_ | _00_;
	assign _05_ = ~(io_in[2] & io_in[1]);
	assign _06_ = _05_ & ~_02_;
	assign _07_ = _02_ & io_in[2];
	assign _08_ = _06_ & ~_07_;
	assign _09_ = ~(io_in[2] ^ io_in[3]);
	assign _10_ = _09_ ^ _08_;
	assign _11_ = _10_ ^ _04_;
	assign io_out[3] = io_in[0] & ~_11_;
	assign io_out[1] = (io_in[0] ? io_in[1] : io_in[2]);
	assign _12_ = _03_ ^ _00_;
	assign io_out[2] = (io_in[0] ? _12_ : io_in[3]);
	assign io_out[13:4] = 10'h000;
	assign \mchip.c.b  = {io_in[0], io_in[0], io_in[0], io_in[0]};
	assign \mchip.c.inst2.in1  = {io_in[2:0], 1'h0};
	assign \mchip.c.inst2.in2  = io_in[3:0];
	assign \mchip.c.inst2.out  = {3'h0, io_in[0]};
	assign \mchip.c.inst2.rem  = 4'h0;
	assign \mchip.c.inst3.in1  = {3'h0, io_in[0]};
	assign \mchip.c.inst3.in2  = 4'h1;
	assign \mchip.c.inst3.rem  = {3'h0, io_in[0]};
	assign \mchip.c.n  = io_in[3:0];
	assign \mchip.c.out  = io_out[3:0];
	assign \mchip.c.out_even  = {1'h0, io_in[3:1]};
	assign \mchip.c.tmp  = {io_in[2:0], 1'h0};
	assign \mchip.c.tmp2  = {3'h0, io_in[0]};
	assign \mchip.io_in  = io_in[7:0];
	assign \mchip.io_out  = {4'h0, io_out[3:0]};
endmodule
module d35_ckasuba_comparator (
	io_in,
	io_out
);
	wire _00_;
	wire _01_;
	wire _02_;
	wire _03_;
	wire _04_;
	wire _05_;
	wire _06_;
	wire _07_;
	wire _08_;
	wire _09_;
	wire _10_;
	wire _11_;
	wire _12_;
	wire _13_;
	wire _14_;
	wire _15_;
	wire _16_;
	wire _17_;
	wire _18_;
	wire _19_;
	wire _20_;
	wire _21_;
	wire _22_;
	wire _23_;
	wire _24_;
	input wire [13:0] io_in;
	output wire [13:0] io_out;
	wire \mchip.and1.b ;
	wire \mchip.and2.a ;
	wire \mchip.and3.b ;
	wire \mchip.and4.a ;
	wire \mchip.and5.b ;
	wire \mchip.and6.a ;
	wire \mchip.and7.b ;
	wire \mchip.and8.a ;
	wire [7:0] \mchip.io_in ;
	wire [7:0] \mchip.io_out ;
	wire \mchip.net1 ;
	wire \mchip.net10 ;
	wire \mchip.net11 ;
	wire \mchip.net12 ;
	wire \mchip.net13 ;
	wire \mchip.net14 ;
	wire \mchip.net15 ;
	wire \mchip.net2 ;
	wire \mchip.net3 ;
	wire \mchip.net4 ;
	wire \mchip.net5 ;
	wire \mchip.net6 ;
	wire \mchip.net7 ;
	wire \mchip.net8 ;
	wire \mchip.net9 ;
	wire \mchip.not1.in ;
	wire \mchip.not10.in ;
	wire \mchip.not11.in ;
	wire \mchip.not2.in ;
	wire \mchip.not4.in ;
	wire \mchip.not5.in ;
	wire \mchip.not7.in ;
	wire \mchip.not8.in ;
	wire \mchip.or10.out ;
	wire \mchip.or11.a ;
	wire \mchip.or11.out ;
	wire \mchip.or12.a ;
	wire \mchip.or12.b ;
	wire \mchip.or12.out ;
	wire \mchip.or7.out ;
	assign _00_ = ~(io_in[0] ^ io_in[4]);
	assign _01_ = io_in[5] ^ io_in[1];
	assign _02_ = _00_ & ~_01_;
	assign _03_ = io_in[6] | ~io_in[2];
	assign _04_ = io_in[2] | ~io_in[6];
	assign _05_ = ~(_04_ & _03_);
	assign _06_ = _02_ & ~_05_;
	assign _07_ = io_in[3] | ~io_in[7];
	assign _08_ = _06_ & ~_07_;
	assign _09_ = _02_ & ~_04_;
	assign _10_ = _09_ | _08_;
	assign _11_ = io_in[1] | ~io_in[5];
	assign _12_ = _00_ & ~_11_;
	assign _13_ = io_in[4] & ~io_in[0];
	assign _14_ = _13_ | _12_;
	assign \mchip.net12  = _14_ | _10_;
	assign _15_ = io_in[7] | ~io_in[3];
	assign _16_ = _06_ & ~_15_;
	assign _17_ = _02_ & ~_03_;
	assign _18_ = _17_ | _16_;
	assign _19_ = io_in[5] | ~io_in[1];
	assign _20_ = _00_ & ~_19_;
	assign _21_ = io_in[0] & ~io_in[4];
	assign _22_ = _21_ | _20_;
	assign \mchip.net10  = _22_ | _18_;
	assign \mchip.net11  = \mchip.net10  | \mchip.net12 ;
	assign _23_ = ~(_15_ & _07_);
	assign _24_ = _06_ & ~_23_;
	assign \mchip.net9  = _24_ | \mchip.net10 ;
	assign io_out = {8'h01, \mchip.net11 , \mchip.net11 , \mchip.net12 , \mchip.net11 , \mchip.net10 , \mchip.net9 };
	assign \mchip.and1.b  = io_in[4];
	assign \mchip.and2.a  = io_in[0];
	assign \mchip.and3.b  = io_in[5];
	assign \mchip.and4.a  = io_in[1];
	assign \mchip.and5.b  = io_in[6];
	assign \mchip.and6.a  = io_in[2];
	assign \mchip.and7.b  = io_in[7];
	assign \mchip.and8.a  = io_in[3];
	assign \mchip.io_in  = io_in[7:0];
	assign \mchip.io_out  = {2'h1, \mchip.net11 , \mchip.net11 , \mchip.net12 , \mchip.net11 , \mchip.net10 , \mchip.net9 };
	assign \mchip.net1  = io_in[0];
	assign \mchip.net13  = 1'h1;
	assign \mchip.net14  = 1'h0;
	assign \mchip.net15  = 1'h1;
	assign \mchip.net2  = io_in[1];
	assign \mchip.net3  = io_in[2];
	assign \mchip.net4  = io_in[3];
	assign \mchip.net5  = io_in[4];
	assign \mchip.net6  = io_in[5];
	assign \mchip.net7  = io_in[6];
	assign \mchip.net8  = io_in[7];
	assign \mchip.not1.in  = io_in[0];
	assign \mchip.not10.in  = io_in[3];
	assign \mchip.not11.in  = io_in[7];
	assign \mchip.not2.in  = io_in[4];
	assign \mchip.not4.in  = io_in[1];
	assign \mchip.not5.in  = io_in[5];
	assign \mchip.not7.in  = io_in[2];
	assign \mchip.not8.in  = io_in[6];
	assign \mchip.or10.out  = \mchip.net10 ;
	assign \mchip.or11.a  = \mchip.net10 ;
	assign \mchip.or11.out  = \mchip.net9 ;
	assign \mchip.or12.a  = \mchip.net12 ;
	assign \mchip.or12.b  = \mchip.net10 ;
	assign \mchip.or12.out  = \mchip.net11 ;
	assign \mchip.or7.out  = \mchip.net12 ;
endmodule
module d36_jxli_fpmul (
	io_in,
	io_out
);
	wire _000_;
	wire _001_;
	wire _002_;
	wire _003_;
	wire _004_;
	wire _005_;
	wire _006_;
	wire _007_;
	wire _008_;
	wire _009_;
	wire _010_;
	wire _011_;
	wire _012_;
	wire _013_;
	wire _014_;
	wire _015_;
	wire _016_;
	wire _017_;
	wire _018_;
	wire _019_;
	wire _020_;
	wire _021_;
	wire _022_;
	wire _023_;
	wire _024_;
	wire _025_;
	wire _026_;
	wire _027_;
	wire _028_;
	wire _029_;
	wire _030_;
	wire _031_;
	wire _032_;
	wire _033_;
	wire _034_;
	wire _035_;
	wire _036_;
	wire _037_;
	wire _038_;
	wire _039_;
	wire _040_;
	wire _041_;
	wire _042_;
	wire _043_;
	wire _044_;
	wire _045_;
	wire _046_;
	wire _047_;
	wire _048_;
	wire _049_;
	wire _050_;
	wire _051_;
	wire _052_;
	wire _053_;
	wire _054_;
	wire _055_;
	wire _056_;
	wire _057_;
	wire _058_;
	wire _059_;
	wire _060_;
	wire _061_;
	wire _062_;
	wire _063_;
	wire _064_;
	wire _065_;
	wire _066_;
	wire _067_;
	wire _068_;
	wire _069_;
	wire _070_;
	wire _071_;
	wire _072_;
	wire _073_;
	wire _074_;
	wire _075_;
	wire _076_;
	wire _077_;
	wire _078_;
	wire _079_;
	wire _080_;
	wire _081_;
	wire _082_;
	wire _083_;
	wire _084_;
	wire _085_;
	wire _086_;
	wire _087_;
	wire _088_;
	wire _089_;
	wire _090_;
	wire _091_;
	wire _092_;
	wire _093_;
	wire _094_;
	wire _095_;
	wire _096_;
	wire _097_;
	wire _098_;
	wire _099_;
	wire _100_;
	wire _101_;
	wire _102_;
	wire _103_;
	wire _104_;
	wire _105_;
	wire _106_;
	wire _107_;
	wire _108_;
	wire _109_;
	wire _110_;
	wire _111_;
	wire _112_;
	wire _113_;
	wire _114_;
	wire _115_;
	wire _116_;
	wire _117_;
	wire _118_;
	wire _119_;
	wire _120_;
	wire _121_;
	wire _122_;
	wire _123_;
	wire _124_;
	wire _125_;
	wire _126_;
	wire _127_;
	wire _128_;
	wire _129_;
	wire _130_;
	wire _131_;
	wire _132_;
	wire _133_;
	wire _134_;
	wire _135_;
	wire _136_;
	wire _137_;
	wire _138_;
	wire _139_;
	wire _140_;
	wire _141_;
	wire _142_;
	wire _143_;
	wire _144_;
	wire _145_;
	wire _146_;
	wire _147_;
	wire _148_;
	wire _149_;
	wire _150_;
	wire _151_;
	wire _152_;
	wire _153_;
	wire _154_;
	wire _155_;
	wire _156_;
	wire _157_;
	wire _158_;
	wire _159_;
	wire _160_;
	wire _161_;
	wire _162_;
	wire _163_;
	wire _164_;
	wire _165_;
	wire _166_;
	wire _167_;
	wire _168_;
	wire _169_;
	wire _170_;
	wire _171_;
	wire _172_;
	wire _173_;
	wire _174_;
	wire _175_;
	wire _176_;
	wire _177_;
	wire _178_;
	wire _179_;
	wire _180_;
	wire _181_;
	wire _182_;
	wire _183_;
	wire _184_;
	wire _185_;
	wire _186_;
	wire _187_;
	wire _188_;
	wire _189_;
	wire _190_;
	wire _191_;
	wire _192_;
	wire _193_;
	wire _194_;
	wire _195_;
	wire _196_;
	wire _197_;
	wire _198_;
	wire _199_;
	wire _200_;
	wire _201_;
	wire _202_;
	wire _203_;
	wire _204_;
	wire _205_;
	wire _206_;
	wire _207_;
	wire _208_;
	wire _209_;
	wire _210_;
	wire _211_;
	wire _212_;
	wire _213_;
	wire _214_;
	wire _215_;
	wire _216_;
	wire _217_;
	wire _218_;
	wire _219_;
	wire _220_;
	wire _221_;
	wire _222_;
	wire _223_;
	wire _224_;
	wire _225_;
	wire _226_;
	wire _227_;
	wire _228_;
	wire _229_;
	wire _230_;
	wire _231_;
	wire _232_;
	wire _233_;
	wire _234_;
	wire _235_;
	wire _236_;
	wire _237_;
	wire _238_;
	wire _239_;
	wire _240_;
	wire _241_;
	wire _242_;
	wire _243_;
	wire _244_;
	wire _245_;
	wire _246_;
	wire _247_;
	wire _248_;
	wire _249_;
	wire _250_;
	wire _251_;
	wire _252_;
	wire _253_;
	wire _254_;
	wire _255_;
	wire _256_;
	wire _257_;
	wire _258_;
	wire _259_;
	wire _260_;
	wire _261_;
	wire _262_;
	wire _263_;
	wire _264_;
	wire _265_;
	wire _266_;
	wire _267_;
	wire _268_;
	wire _269_;
	wire _270_;
	wire _271_;
	wire _272_;
	wire _273_;
	wire _274_;
	wire _275_;
	wire _276_;
	wire _277_;
	wire _278_;
	wire _279_;
	wire _280_;
	wire _281_;
	wire _282_;
	wire _283_;
	wire _284_;
	wire _285_;
	wire _286_;
	wire _287_;
	wire _288_;
	wire _289_;
	wire _290_;
	wire _291_;
	wire _292_;
	wire _293_;
	wire _294_;
	wire _295_;
	wire _296_;
	wire _297_;
	wire _298_;
	wire _299_;
	wire _300_;
	wire _301_;
	wire _302_;
	wire _303_;
	wire _304_;
	wire _305_;
	wire _306_;
	wire _307_;
	wire _308_;
	wire _309_;
	wire _310_;
	wire _311_;
	wire _312_;
	wire _313_;
	wire _314_;
	wire _315_;
	wire _316_;
	wire _317_;
	wire _318_;
	wire _319_;
	wire _320_;
	wire _321_;
	wire _322_;
	wire _323_;
	wire _324_;
	wire _325_;
	wire _326_;
	wire _327_;
	wire _328_;
	wire _329_;
	wire _330_;
	wire _331_;
	wire _332_;
	wire _333_;
	wire _334_;
	wire _335_;
	wire _336_;
	wire _337_;
	wire _338_;
	wire _339_;
	wire _340_;
	wire _341_;
	wire _342_;
	wire _343_;
	wire _344_;
	wire _345_;
	wire _346_;
	wire _347_;
	wire _348_;
	wire _349_;
	wire _350_;
	wire _351_;
	wire _352_;
	wire _353_;
	wire _354_;
	wire _355_;
	wire _356_;
	wire _357_;
	wire _358_;
	wire _359_;
	wire _360_;
	wire [3:0] _361_;
	wire [4:0] _362_;
	wire [4:0] _363_;
	wire _364_;
	input wire [13:0] io_in;
	output wire [13:0] io_out;
	wire [6:0] \mchip.NaN ;
	reg [7:0] \mchip.a ;
	reg [4:0] \mchip.ae ;
	reg [3:0] \mchip.am ;
	reg [7:0] \mchip.b ;
	reg [4:0] \mchip.be ;
	reg [3:0] \mchip.bm ;
	reg [7:0] \mchip.c ;
	reg [4:0] \mchip.ce ;
	wire \mchip.clock ;
	reg [3:0] \mchip.cm ;
	wire [3:0] \mchip.data ;
	wire \mchip.enable ;
	wire [6:0] \mchip.infty ;
	wire [7:0] \mchip.io_in ;
	wire [7:0] \mchip.io_out ;
	wire [7:0] \mchip.product ;
	wire \mchip.reset ;
	wire [12:0] \mchip.state ;
	assign _042_ = ~(\mchip.state [8] & \mchip.cm [3]);
	assign _043_ = \mchip.ce [3] & ~\mchip.ce [2];
	assign _044_ = \mchip.ce [0] & \mchip.ce [1];
	assign _045_ = _043_ & ~_044_;
	assign _046_ = \mchip.ce [3] & ~_045_;
	assign _047_ = \mchip.ce [4] & ~_046_;
	assign _048_ = \mchip.ce [1] & ~\mchip.ce [0];
	assign _049_ = ~(_048_ & _043_);
	assign _050_ = \mchip.ce [4] & ~_049_;
	assign _051_ = _047_ & ~_050_;
	assign _052_ = \mchip.state [5] & ~_051_;
	assign _053_ = _042_ & ~_052_;
	assign _054_ = ~(\mchip.state [1] | \mchip.state [5]);
	assign _055_ = _054_ & ~\mchip.state [8];
	assign _018_ = _053_ & ~_055_;
	assign _017_ = ~(_055_ | _052_);
	assign _016_ = io_in[2] & \mchip.state [7];
	assign _015_ = \mchip.state [0] & io_in[2];
	assign _056_ = io_in[1] | io_in[2];
	assign _057_ = \mchip.state [0] & ~_056_;
	assign _004_ = _057_ | io_in[1];
	assign _014_ = \mchip.state [10] & io_in[2];
	assign _013_ = \mchip.state [4] & io_in[2];
	assign _058_ = \mchip.state [4] & ~_056_;
	assign _059_ = io_in[1] | ~io_in[2];
	assign _060_ = \mchip.state [7] & ~_059_;
	assign _007_ = _060_ | _058_;
	assign _061_ = ~\mchip.ae [4];
	assign _062_ = \mchip.ae [0] | \mchip.ae [1];
	assign _063_ = \mchip.ae [2] | ~\mchip.ae [3];
	assign _064_ = _063_ | _062_;
	assign _065_ = _061_ & ~_064_;
	assign _066_ = ~(\mchip.am [3] | \mchip.am [2]);
	assign _067_ = \mchip.am [0] | \mchip.am [1];
	assign _068_ = _067_ | ~_066_;
	assign _069_ = _065_ & ~_068_;
	assign _070_ = ~(\mchip.bm [3] | \mchip.bm [2]);
	assign _071_ = \mchip.bm [0] | \mchip.bm [1];
	assign _072_ = _070_ & ~_071_;
	assign _073_ = \mchip.be [0] | \mchip.be [1];
	assign _074_ = \mchip.be [2] | ~\mchip.be [3];
	assign _075_ = _074_ | _073_;
	assign _076_ = _075_ | \mchip.be [4];
	assign _077_ = ~(_076_ | _072_);
	assign _078_ = _068_ & _065_;
	assign _079_ = _078_ | _077_;
	assign _080_ = _072_ & ~_076_;
	assign _081_ = _080_ | _079_;
	assign _082_ = ~\mchip.state [9];
	assign _083_ = ~\mchip.be [4];
	assign _084_ = \mchip.be [1] | ~\mchip.be [0];
	assign _085_ = _084_ | _074_;
	assign _086_ = _085_ | _083_;
	assign _087_ = _072_ & ~_086_;
	assign _088_ = \mchip.ae [1] | ~\mchip.ae [0];
	assign _089_ = _088_ | _063_;
	assign _090_ = _089_ | _061_;
	assign _091_ = ~(_090_ | _068_);
	assign _092_ = _091_ | _087_;
	assign _093_ = _092_ | _082_;
	assign _094_ = _093_ | _081_;
	assign _095_ = _094_ | _069_;
	assign _096_ = ~(\mchip.state [11] | \mchip.state [9]);
	assign _012_ = _095_ & ~_096_;
	assign _097_ = \mchip.state [1] & ~io_in[1];
	assign _098_ = io_in[1] | \mchip.cm [3];
	assign _099_ = \mchip.state [8] & ~_098_;
	assign _011_ = _099_ | _097_;
	assign _100_ = \mchip.state [4] & ~_059_;
	assign _101_ = \mchip.state [10] & ~_056_;
	assign _005_ = _101_ | _100_;
	assign _102_ = \mchip.state [0] & ~_059_;
	assign _103_ = \mchip.state [7] & ~_056_;
	assign _010_ = _103_ | _102_;
	assign _104_ = io_in[1] | ~\mchip.am [3];
	assign _105_ = \mchip.state [6] & ~_104_;
	assign _106_ = \mchip.bm [3] | io_in[1];
	assign _107_ = \mchip.state [12] & ~_106_;
	assign _006_ = _107_ | _105_;
	assign _108_ = _080_ | _069_;
	assign _109_ = _092_ | _079_;
	assign _110_ = ~(_090_ & \mchip.state [9]);
	assign _111_ = _110_ | _109_;
	assign _112_ = _111_ | _108_;
	assign _113_ = \mchip.state [2] | \mchip.state [6];
	assign _114_ = _082_ & ~_113_;
	assign _115_ = _112_ & ~_114_;
	assign _116_ = _079_ & ~_082_;
	assign _117_ = \mchip.state [6] & \mchip.am [3];
	assign _118_ = _117_ | _116_;
	assign _119_ = _115_ & ~_118_;
	assign _120_ = ~(_092_ & \mchip.state [9]);
	assign _121_ = _120_ | _081_;
	assign _122_ = ~(_121_ | _069_);
	assign _123_ = _080_ & ~_069_;
	assign _124_ = _079_ | _082_;
	assign _125_ = _123_ & ~_124_;
	assign _126_ = _069_ & ~_124_;
	assign _127_ = _126_ | _125_;
	assign _128_ = _127_ | _122_;
	assign _024_ = _119_ & ~_128_;
	assign _129_ = ~(_086_ & \mchip.state [9]);
	assign _130_ = _129_ | _109_;
	assign _131_ = _130_ | _108_;
	assign _132_ = \mchip.state [12] & \mchip.bm [3];
	assign _133_ = _131_ & ~_132_;
	assign _134_ = _126_ | _116_;
	assign _135_ = _133_ & ~_134_;
	assign _136_ = ~(\mchip.state [2] | \mchip.state [9]);
	assign _137_ = _136_ & ~\mchip.state [12];
	assign _138_ = _125_ | _122_;
	assign _139_ = _138_ | _137_;
	assign _023_ = _135_ & ~_139_;
	assign _140_ = _092_ | io_in[1];
	assign _141_ = _140_ | _081_;
	assign _142_ = _141_ | _069_;
	assign _143_ = \mchip.state [9] & ~_142_;
	assign _144_ = \mchip.am [3] | io_in[1];
	assign _145_ = \mchip.state [6] & ~_144_;
	assign _009_ = _145_ | _143_;
	assign _146_ = io_in[1] | ~_051_;
	assign _147_ = \mchip.state [5] & ~_146_;
	assign _148_ = io_in[1] | ~\mchip.cm [3];
	assign _149_ = \mchip.state [8] & ~_148_;
	assign _008_ = _149_ | _147_;
	assign _150_ = _090_ | _082_;
	assign _151_ = _150_ | _109_;
	assign _152_ = ~(_151_ | _108_);
	assign _153_ = _152_ | _114_;
	assign _154_ = _153_ | _134_;
	assign _022_ = ~(_154_ | _138_);
	assign _021_ = _113_ & ~_117_;
	assign _155_ = ~\mchip.bm [3];
	assign _020_ = (\mchip.state [12] ? _155_ : \mchip.state [2]);
	assign _156_ = ~(_138_ | _134_);
	assign _157_ = _086_ | _082_;
	assign _158_ = _157_ | _109_;
	assign _159_ = ~(_158_ | _108_);
	assign _160_ = _159_ | _137_;
	assign _019_ = _156_ & ~_160_;
	assign _161_ = ~\mchip.ce [0];
	assign _162_ = \mchip.state [5] | \mchip.state [8];
	assign _163_ = ~(\mchip.be [0] ^ \mchip.ae [0]);
	assign _029_ = (_162_ ? _161_ : _163_);
	assign _164_ = ~(\mchip.state [5] ^ \mchip.ce [1]);
	assign _165_ = _164_ ^ \mchip.ce [0];
	assign _166_ = \mchip.be [0] | \mchip.ae [0];
	assign _167_ = \mchip.be [1] ^ \mchip.ae [1];
	assign _168_ = _167_ ^ _166_;
	assign _030_ = (_162_ ? _165_ : _168_);
	assign _169_ = \mchip.ce [1] & ~\mchip.state [5];
	assign _170_ = _164_ & ~_161_;
	assign _171_ = _170_ | _169_;
	assign _172_ = ~(\mchip.state [5] ^ \mchip.ce [2]);
	assign _173_ = _172_ ^ _171_;
	assign _174_ = \mchip.be [1] & \mchip.ae [1];
	assign _175_ = _167_ & _166_;
	assign _176_ = _175_ | _174_;
	assign _177_ = \mchip.be [2] ^ \mchip.ae [2];
	assign _178_ = _177_ ^ _176_;
	assign _031_ = (_162_ ? _173_ : _178_);
	assign _179_ = \mchip.ce [2] & ~\mchip.state [5];
	assign _180_ = _172_ & _171_;
	assign _181_ = _180_ | _179_;
	assign _182_ = ~(\mchip.state [5] ^ \mchip.ce [3]);
	assign _183_ = _182_ ^ _181_;
	assign _184_ = \mchip.be [2] & \mchip.ae [2];
	assign _185_ = _177_ & _176_;
	assign _186_ = _185_ | _184_;
	assign _187_ = \mchip.be [3] ^ \mchip.ae [3];
	assign _188_ = _187_ ^ _186_;
	assign _032_ = (_162_ ? _183_ : _188_);
	assign _189_ = \mchip.ce [3] & ~\mchip.state [5];
	assign _190_ = _182_ & _179_;
	assign _191_ = _190_ | _189_;
	assign _192_ = ~(_182_ & _172_);
	assign _193_ = _171_ & ~_192_;
	assign _194_ = _193_ | _191_;
	assign _195_ = ~(\mchip.state [5] ^ \mchip.ce [4]);
	assign _196_ = _195_ ^ _194_;
	assign _197_ = \mchip.be [3] & \mchip.ae [3];
	assign _198_ = _187_ & _184_;
	assign _199_ = _198_ | _197_;
	assign _200_ = ~(_187_ & _177_);
	assign _201_ = _176_ & ~_200_;
	assign _202_ = _201_ | _199_;
	assign _203_ = \mchip.be [4] ^ \mchip.ae [4];
	assign _204_ = _203_ ^ _202_;
	assign _033_ = (_162_ ? _196_ : _204_);
	assign _205_ = _108_ | _079_;
	assign _206_ = \mchip.cm [3] | ~_050_;
	assign _207_ = _206_ & ~\mchip.ce [0];
	assign _208_ = \mchip.ce [3] & ~\mchip.ce [4];
	assign _209_ = _208_ | _207_;
	assign _034_ = (\mchip.state [11] ? _209_ : _205_);
	assign _210_ = \mchip.ce [0] ^ \mchip.ce [1];
	assign _211_ = _206_ & ~_210_;
	assign _212_ = _211_ | _208_;
	assign _035_ = (\mchip.state [11] ? _212_ : _205_);
	assign _213_ = ~(\mchip.ce [0] | \mchip.ce [1]);
	assign _214_ = ~(_213_ ^ \mchip.ce [2]);
	assign _215_ = _206_ & ~_214_;
	assign _216_ = _215_ | _208_;
	assign _036_ = (\mchip.state [11] ? _216_ : _205_);
	assign _217_ = _213_ & ~\mchip.ce [2];
	assign _218_ = _217_ ^ \mchip.ce [3];
	assign _219_ = _206_ & ~_218_;
	assign _220_ = _219_ | _208_;
	assign _037_ = (\mchip.state [11] ? _220_ : _205_);
	assign _025_ = (\mchip.state [6] ? \mchip.am [0] : \mchip.a [1]);
	assign _026_ = (\mchip.state [6] ? \mchip.am [1] : \mchip.a [2]);
	assign _027_ = (\mchip.state [12] ? \mchip.bm [0] : \mchip.b [1]);
	assign _028_ = (\mchip.state [12] ? \mchip.bm [1] : \mchip.b [2]);
	assign _221_ = _091_ & _080_;
	assign _222_ = (_069_ ? _087_ : _221_);
	assign _223_ = _222_ | _079_;
	assign _224_ = \mchip.cm [0] & ~_208_;
	assign _038_ = (\mchip.state [11] ? _224_ : _223_);
	assign _225_ = \mchip.cm [1] & ~_208_;
	assign _039_ = (\mchip.state [11] ? _225_ : _223_);
	assign _226_ = \mchip.cm [2] & ~_208_;
	assign _040_ = (\mchip.state [11] ? _226_ : _223_);
	assign _227_ = ~\mchip.a [3];
	assign _228_ = \mchip.state [6] & ~\mchip.ae [0];
	assign _229_ = _228_ | \mchip.state [9];
	assign _230_ = ~(\mchip.state [6] | \mchip.state [9]);
	assign _363_[0] = (_230_ ? _227_ : _229_);
	assign _231_ = ~_230_;
	assign _232_ = \mchip.ae [0] ^ \mchip.ae [1];
	assign _233_ = \mchip.state [6] & ~_232_;
	assign _234_ = \mchip.a [4] ^ \mchip.a [3];
	assign _363_[1] = (_230_ ? _234_ : _233_);
	assign _235_ = _062_ ^ \mchip.ae [2];
	assign _236_ = \mchip.state [6] & ~_235_;
	assign _237_ = \mchip.a [4] & \mchip.a [3];
	assign _238_ = _237_ ^ \mchip.a [5];
	assign _363_[2] = (_230_ ? _238_ : _236_);
	assign _239_ = _062_ | \mchip.ae [2];
	assign _240_ = _239_ ^ \mchip.ae [3];
	assign _241_ = \mchip.state [6] & ~_240_;
	assign _242_ = _241_ | \mchip.state [9];
	assign _243_ = ~\mchip.a [6];
	assign _244_ = _237_ & \mchip.a [5];
	assign _245_ = _244_ ^ _243_;
	assign _363_[3] = (_230_ ? _245_ : _242_);
	assign _246_ = ~(\mchip.ae [3] | \mchip.ae [2]);
	assign _247_ = _246_ & ~_062_;
	assign _248_ = _247_ ^ _061_;
	assign _249_ = \mchip.state [6] & ~_248_;
	assign _250_ = _249_ | \mchip.state [9];
	assign _251_ = \mchip.a [6] | ~\mchip.a [5];
	assign _252_ = _237_ & ~_251_;
	assign _253_ = _243_ & ~_252_;
	assign _363_[4] = (_230_ ? _253_ : _250_);
	assign _254_ = ~\mchip.b [3];
	assign _255_ = \mchip.state [12] & ~\mchip.be [0];
	assign _256_ = _255_ | \mchip.state [9];
	assign _257_ = ~(\mchip.state [12] | \mchip.state [9]);
	assign _362_[0] = (_257_ ? _254_ : _256_);
	assign _258_ = ~_257_;
	assign _259_ = \mchip.be [0] ^ \mchip.be [1];
	assign _260_ = \mchip.state [12] & ~_259_;
	assign _261_ = \mchip.b [4] ^ \mchip.b [3];
	assign _362_[1] = (_257_ ? _261_ : _260_);
	assign _262_ = _073_ ^ \mchip.be [2];
	assign _263_ = \mchip.state [12] & ~_262_;
	assign _264_ = \mchip.b [4] & \mchip.b [3];
	assign _265_ = _264_ ^ \mchip.b [5];
	assign _362_[2] = (_257_ ? _265_ : _263_);
	assign _266_ = _073_ | \mchip.be [2];
	assign _267_ = _266_ ^ \mchip.be [3];
	assign _268_ = \mchip.state [12] & ~_267_;
	assign _269_ = _268_ | \mchip.state [9];
	assign _270_ = ~\mchip.b [6];
	assign _271_ = _264_ & \mchip.b [5];
	assign _272_ = _271_ ^ _270_;
	assign _362_[3] = (_257_ ? _272_ : _269_);
	assign _273_ = ~(\mchip.be [3] | \mchip.be [2]);
	assign _274_ = _273_ & ~_073_;
	assign _275_ = _274_ ^ _083_;
	assign _276_ = \mchip.state [12] & ~_275_;
	assign _277_ = _276_ | \mchip.state [9];
	assign _278_ = \mchip.b [6] | ~\mchip.b [5];
	assign _279_ = _264_ & ~_278_;
	assign _280_ = _270_ & ~_279_;
	assign _362_[4] = (_257_ ? _280_ : _277_);
	assign _281_ = \mchip.cm [1] & \mchip.state [5];
	assign _282_ = \mchip.bm [1] & \mchip.am [0];
	assign _283_ = ~(\mchip.bm [0] & \mchip.am [1]);
	assign _284_ = _282_ & ~_283_;
	assign _285_ = ~(\mchip.bm [1] & \mchip.am [1]);
	assign _286_ = \mchip.bm [0] & \mchip.am [2];
	assign _287_ = _286_ ^ _285_;
	assign _288_ = ~(\mchip.bm [2] & \mchip.am [0]);
	assign _289_ = ~_288_;
	assign _290_ = _289_ ^ _287_;
	assign _291_ = _284_ & ~_290_;
	assign _292_ = \mchip.bm [3] & \mchip.am [0];
	assign _293_ = _285_ | ~_286_;
	assign _294_ = _289_ & ~_287_;
	assign _295_ = _294_ | ~_293_;
	assign _296_ = ~(\mchip.bm [2] & \mchip.am [1]);
	assign _297_ = \mchip.bm [1] & \mchip.am [2];
	assign _298_ = ~(\mchip.bm [0] & \mchip.am [3]);
	assign _299_ = _298_ ^ _297_;
	assign _300_ = ~(_299_ ^ _296_);
	assign _301_ = _300_ ^ _295_;
	assign _302_ = _301_ ^ _292_;
	assign _303_ = ~(_302_ ^ _291_);
	assign _361_[0] = (_162_ ? _281_ : _303_);
	assign _304_ = \mchip.cm [3] | ~\mchip.cm [0];
	assign _305_ = \mchip.state [8] & ~_304_;
	assign _306_ = \mchip.cm [2] & \mchip.state [5];
	assign _307_ = _306_ | _305_;
	assign _308_ = _291_ & ~_302_;
	assign _309_ = _292_ & ~_301_;
	assign _310_ = _295_ & ~_300_;
	assign _311_ = _310_ | _309_;
	assign _312_ = \mchip.bm [3] & \mchip.am [1];
	assign _313_ = _299_ | _296_;
	assign _314_ = _297_ & ~_298_;
	assign _315_ = _314_ | ~_313_;
	assign _316_ = ~(\mchip.bm [2] & \mchip.am [2]);
	assign _317_ = \mchip.bm [1] & \mchip.am [3];
	assign _318_ = _317_ ^ _316_;
	assign _319_ = _318_ ^ _315_;
	assign _320_ = ~(_319_ ^ _312_);
	assign _321_ = ~(_320_ ^ _311_);
	assign _322_ = ~(_321_ ^ _308_);
	assign _361_[1] = (_162_ ? _307_ : _322_);
	assign _323_ = \mchip.cm [3] | ~\mchip.cm [1];
	assign _324_ = \mchip.state [8] & ~_323_;
	assign _325_ = \mchip.state [5] & \mchip.cm [3];
	assign _326_ = _325_ | _324_;
	assign _327_ = _320_ & _311_;
	assign _328_ = _308_ & ~_321_;
	assign _329_ = ~(_328_ | _327_);
	assign _330_ = _312_ & ~_319_;
	assign _331_ = _315_ & ~_318_;
	assign _332_ = _331_ | _330_;
	assign _333_ = \mchip.bm [3] & \mchip.am [2];
	assign _334_ = _316_ | ~_317_;
	assign _335_ = \mchip.bm [2] & \mchip.am [3];
	assign _336_ = _335_ ^ _334_;
	assign _337_ = ~(_336_ ^ _333_);
	assign _338_ = ~(_337_ ^ _332_);
	assign _339_ = _338_ ^ _329_;
	assign _361_[2] = (_162_ ? _326_ : _339_);
	assign _340_ = ~(\mchip.cm [2] | \mchip.cm [3]);
	assign _341_ = \mchip.state [8] & ~_340_;
	assign _342_ = _337_ & _332_;
	assign _343_ = _327_ & ~_338_;
	assign _344_ = _343_ | _342_;
	assign _345_ = _338_ | _321_;
	assign _346_ = _308_ & ~_345_;
	assign _347_ = _346_ | _344_;
	assign _348_ = _333_ & ~_336_;
	assign _349_ = _335_ & ~_334_;
	assign _350_ = _349_ | _348_;
	assign _351_ = \mchip.bm [3] & \mchip.am [3];
	assign _352_ = _351_ ^ _350_;
	assign _353_ = _352_ ^ _347_;
	assign _361_[3] = (_162_ ? _341_ : _353_);
	assign _354_ = \mchip.state [12] & ~_070_;
	assign _355_ = _082_ & ~_354_;
	assign _360_ = _258_ & ~_355_;
	assign _356_ = \mchip.state [6] & ~_066_;
	assign _357_ = _082_ & ~_356_;
	assign _364_ = _231_ & ~_357_;
	assign _002_ = \mchip.state [2] & ~io_in[1];
	assign _358_ = _051_ | io_in[1];
	assign _003_ = \mchip.state [5] & ~_358_;
	assign _041_ = \mchip.a [7] ^ \mchip.b [7];
	assign _001_ = \mchip.state [10] & ~_059_;
	assign _359_ = io_in[1] | ~\mchip.bm [3];
	assign _000_ = \mchip.state [12] & ~_359_;
	always @(posedge io_in[0])
		if (_013_)
			\mchip.b [4] <= io_in[3];
	always @(posedge io_in[0])
		if (_013_)
			\mchip.b [5] <= io_in[4];
	always @(posedge io_in[0])
		if (_013_)
			\mchip.b [6] <= io_in[5];
	always @(posedge io_in[0])
		if (_013_)
			\mchip.b [7] <= io_in[6];
	always @(posedge io_in[0])
		if (_018_)
			\mchip.cm [0] <= _361_[0];
	always @(posedge io_in[0])
		if (_018_)
			\mchip.cm [1] <= _361_[1];
	always @(posedge io_in[0])
		if (_018_)
			\mchip.cm [2] <= _361_[2];
	always @(posedge io_in[0])
		if (_016_)
			\mchip.a [0] <= io_in[3];
	always @(posedge io_in[0])
		if (_016_)
			\mchip.a [1] <= io_in[4];
	always @(posedge io_in[0])
		if (_016_)
			\mchip.a [2] <= io_in[5];
	always @(posedge io_in[0])
		if (_016_)
			\mchip.a [3] <= io_in[6];
	always @(posedge io_in[0])
		if (_014_)
			\mchip.b [0] <= io_in[3];
	always @(posedge io_in[0])
		if (_014_)
			\mchip.b [1] <= io_in[4];
	always @(posedge io_in[0])
		if (_014_)
			\mchip.b [2] <= io_in[5];
	always @(posedge io_in[0])
		if (_014_)
			\mchip.b [3] <= io_in[6];
	always @(posedge io_in[0])
		if (_020_)
			if (\mchip.state [12])
				\mchip.bm [0] <= 1'h0;
			else
				\mchip.bm [0] <= \mchip.b [0];
	always @(posedge io_in[0])
		if (_018_)
			\mchip.ce [0] <= _029_;
	always @(posedge io_in[0])
		if (_018_)
			\mchip.ce [1] <= _030_;
	always @(posedge io_in[0])
		if (_018_)
			\mchip.ce [2] <= _031_;
	always @(posedge io_in[0])
		if (_018_)
			\mchip.ce [3] <= _032_;
	always @(posedge io_in[0])
		if (_018_)
			\mchip.ce [4] <= _033_;
	always @(posedge io_in[0])
		if (_023_)
			\mchip.be [0] <= _362_[0];
	always @(posedge io_in[0])
		if (_023_)
			\mchip.be [1] <= _362_[1];
	always @(posedge io_in[0])
		if (_023_)
			\mchip.be [2] <= _362_[2];
	always @(posedge io_in[0])
		if (_023_)
			\mchip.be [3] <= _362_[3];
	always @(posedge io_in[0])
		if (_023_)
			\mchip.be [4] <= _362_[4];
	always @(posedge io_in[0])
		if (_024_)
			\mchip.ae [0] <= _363_[0];
	always @(posedge io_in[0])
		if (_024_)
			\mchip.ae [1] <= _363_[1];
	always @(posedge io_in[0])
		if (_024_)
			\mchip.ae [2] <= _363_[2];
	always @(posedge io_in[0])
		if (_024_)
			\mchip.ae [3] <= _363_[3];
	always @(posedge io_in[0])
		if (_024_)
			\mchip.ae [4] <= _363_[4];
	always @(posedge io_in[0])
		if (_019_)
			\mchip.bm [3] <= _360_;
	always @(posedge io_in[0])
		if (_017_)
			\mchip.cm [3] <= _361_[3];
	always @(posedge io_in[0])
		if (_015_)
			\mchip.a [4] <= io_in[3];
	always @(posedge io_in[0])
		if (_015_)
			\mchip.a [5] <= io_in[4];
	always @(posedge io_in[0])
		if (_015_)
			\mchip.a [6] <= io_in[5];
	always @(posedge io_in[0])
		if (_015_)
			\mchip.a [7] <= io_in[6];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.c [7] <= 1'h1;
		else if (\mchip.state [2])
			\mchip.c [7] <= _041_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.c [0] <= 1'h1;
		else if (_012_)
			\mchip.c [0] <= _038_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.c [1] <= 1'h1;
		else if (_012_)
			\mchip.c [1] <= _039_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.c [2] <= 1'h1;
		else if (_012_)
			\mchip.c [2] <= _040_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.c [3] <= 1'h1;
		else if (_012_)
			\mchip.c [3] <= _034_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.c [4] <= 1'h1;
		else if (_012_)
			\mchip.c [4] <= _035_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.c [5] <= 1'h1;
		else if (_012_)
			\mchip.c [5] <= _036_;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.c [6] <= 1'h1;
		else if (_012_)
			\mchip.c [6] <= _037_;
	reg \mchip.state_reg[0] ;
	always @(posedge io_in[0]) \mchip.state_reg[0]  <= _004_;
	assign \mchip.state [0] = \mchip.state_reg[0] ;
	reg \mchip.state_reg[1] ;
	always @(posedge io_in[0]) \mchip.state_reg[1]  <= _000_;
	assign \mchip.state [1] = \mchip.state_reg[1] ;
	reg \mchip.state_reg[2] ;
	always @(posedge io_in[0]) \mchip.state_reg[2]  <= _001_;
	assign \mchip.state [2] = \mchip.state_reg[2] ;
	reg \mchip.state_reg[4] ;
	always @(posedge io_in[0]) \mchip.state_reg[4]  <= _007_;
	assign \mchip.state [4] = \mchip.state_reg[4] ;
	reg \mchip.state_reg[5] ;
	always @(posedge io_in[0]) \mchip.state_reg[5]  <= _008_;
	assign \mchip.state [5] = \mchip.state_reg[5] ;
	reg \mchip.state_reg[6] ;
	always @(posedge io_in[0]) \mchip.state_reg[6]  <= _009_;
	assign \mchip.state [6] = \mchip.state_reg[6] ;
	reg \mchip.state_reg[7] ;
	always @(posedge io_in[0]) \mchip.state_reg[7]  <= _010_;
	assign \mchip.state [7] = \mchip.state_reg[7] ;
	reg \mchip.state_reg[8] ;
	always @(posedge io_in[0]) \mchip.state_reg[8]  <= _011_;
	assign \mchip.state [8] = \mchip.state_reg[8] ;
	reg \mchip.state_reg[9] ;
	always @(posedge io_in[0]) \mchip.state_reg[9]  <= _002_;
	assign \mchip.state [9] = \mchip.state_reg[9] ;
	reg \mchip.state_reg[10] ;
	always @(posedge io_in[0]) \mchip.state_reg[10]  <= _005_;
	assign \mchip.state [10] = \mchip.state_reg[10] ;
	reg \mchip.state_reg[11] ;
	always @(posedge io_in[0]) \mchip.state_reg[11]  <= _003_;
	assign \mchip.state [11] = \mchip.state_reg[11] ;
	reg \mchip.state_reg[12] ;
	always @(posedge io_in[0]) \mchip.state_reg[12]  <= _006_;
	assign \mchip.state [12] = \mchip.state_reg[12] ;
	always @(posedge io_in[0])
		if (_022_)
			\mchip.am [3] <= _364_;
	always @(posedge io_in[0])
		if (_020_)
			\mchip.bm [1] <= _027_;
	always @(posedge io_in[0])
		if (_020_)
			\mchip.bm [2] <= _028_;
	always @(posedge io_in[0])
		if (_021_)
			\mchip.am [1] <= _025_;
	always @(posedge io_in[0])
		if (_021_)
			\mchip.am [2] <= _026_;
	always @(posedge io_in[0])
		if (_021_)
			if (\mchip.state [6])
				\mchip.am [0] <= 1'h0;
			else
				\mchip.am [0] <= \mchip.a [0];
	assign io_out = {6'h00, \mchip.c };
	assign \mchip.NaN  = 7'h7f;
	assign \mchip.clock  = io_in[0];
	assign \mchip.data  = io_in[6:3];
	assign \mchip.enable  = io_in[2];
	assign \mchip.infty  = 7'h78;
	assign \mchip.io_in  = io_in[7:0];
	assign \mchip.io_out  = \mchip.c ;
	assign \mchip.product  = 8'h00;
	assign \mchip.reset  = io_in[1];
	assign \mchip.state [3] = 1'h0;
endmodule
module d37_sophiali_calculator (
	io_in,
	io_out
);
	wire _000_;
	wire _001_;
	wire _002_;
	wire _003_;
	wire _004_;
	wire _005_;
	wire _006_;
	wire _007_;
	wire _008_;
	wire _009_;
	wire _010_;
	wire _011_;
	wire _012_;
	wire _013_;
	wire _014_;
	wire _015_;
	wire _016_;
	wire _017_;
	wire _018_;
	wire _019_;
	wire _020_;
	wire _021_;
	wire _022_;
	wire _023_;
	wire _024_;
	wire _025_;
	wire _026_;
	wire _027_;
	wire _028_;
	wire _029_;
	wire _030_;
	wire _031_;
	wire _032_;
	wire _033_;
	wire _034_;
	wire _035_;
	wire _036_;
	wire _037_;
	wire _038_;
	wire _039_;
	wire _040_;
	wire _041_;
	wire _042_;
	wire _043_;
	wire _044_;
	wire _045_;
	wire _046_;
	wire _047_;
	wire _048_;
	wire _049_;
	wire _050_;
	wire _051_;
	wire _052_;
	wire _053_;
	wire _054_;
	wire _055_;
	wire _056_;
	wire _057_;
	wire _058_;
	wire _059_;
	wire _060_;
	wire _061_;
	wire _062_;
	wire _063_;
	wire _064_;
	wire _065_;
	wire _066_;
	wire _067_;
	wire _068_;
	wire _069_;
	wire _070_;
	wire _071_;
	wire _072_;
	wire _073_;
	wire _074_;
	wire _075_;
	wire _076_;
	wire _077_;
	wire _078_;
	wire _079_;
	wire _080_;
	wire _081_;
	wire _082_;
	wire _083_;
	wire _084_;
	wire _085_;
	wire _086_;
	wire _087_;
	wire _088_;
	wire _089_;
	wire _090_;
	wire _091_;
	wire _092_;
	wire _093_;
	wire _094_;
	wire [7:0] _095_;
	input wire [13:0] io_in;
	output wire [13:0] io_out;
	wire [1:0] \mchip.arithOp ;
	wire \mchip.clock ;
	wire \mchip.en ;
	wire \mchip.enable ;
	wire [2:0] \mchip.in ;
	wire [7:0] \mchip.io_in ;
	reg [7:0] \mchip.io_out ;
	wire \mchip.nextState ;
	wire \mchip.reset ;
	reg \mchip.state ;
	assign \mchip.enable  = io_in[2] & ~\mchip.state ;
	assign _028_ = io_in[7] & ~io_in[6];
	assign _000_ = \mchip.enable  & ~_028_;
	assign _029_ = ~(io_in[3] ^ \mchip.io_out [0]);
	assign _030_ = _028_ & ~_029_;
	assign _031_ = io_in[6] & io_in[7];
	assign _032_ = ~io_in[5];
	assign _033_ = \mchip.io_out [0] & ~io_in[3];
	assign _034_ = _033_ & ~io_in[4];
	assign _035_ = ~(_034_ & _032_);
	assign _036_ = _031_ & ~_035_;
	assign _037_ = _036_ | _030_;
	assign _038_ = _031_ | _028_;
	assign _039_ = \mchip.io_out [0] | ~io_in[3];
	assign _040_ = _033_ | ~_039_;
	assign _095_[0] = (_038_ ? _037_ : _040_);
	assign _041_ = ~(\mchip.io_out [1] ^ io_in[4]);
	assign _042_ = _028_ & ~_041_;
	assign _043_ = (io_in[3] ? \mchip.io_out [0] : \mchip.io_out [1]);
	assign _044_ = _043_ & ~io_in[4];
	assign _045_ = ~(_044_ & _032_);
	assign _046_ = _031_ & ~_045_;
	assign _047_ = _046_ | _042_;
	assign _048_ = io_in[4] ^ io_in[3];
	assign _049_ = io_in[6] & ~io_in[7];
	assign _050_ = (_049_ ? io_in[4] : _048_);
	assign _051_ = _050_ ^ \mchip.io_out [1];
	assign _052_ = ~(_051_ ^ _039_);
	assign _095_[1] = (_038_ ? _047_ : _052_);
	assign _053_ = ~(\mchip.io_out [2] ^ io_in[5]);
	assign _054_ = _028_ & ~_053_;
	assign _055_ = (io_in[3] ? \mchip.io_out [1] : \mchip.io_out [2]);
	assign _056_ = (io_in[4] ? _033_ : _055_);
	assign _057_ = ~(_056_ & _032_);
	assign _058_ = _031_ & ~_057_;
	assign _059_ = _058_ | _054_;
	assign _060_ = _039_ & ~_051_;
	assign _061_ = \mchip.io_out [1] & ~_050_;
	assign _062_ = _061_ | _060_;
	assign _063_ = ~(io_in[4] | io_in[3]);
	assign _064_ = _063_ ^ _032_;
	assign _065_ = (_049_ ? io_in[5] : _064_);
	assign _066_ = _065_ ^ \mchip.io_out [2];
	assign _067_ = ~(_066_ ^ _062_);
	assign _095_[2] = (_038_ ? _059_ : _067_);
	assign _068_ = (io_in[3] ? \mchip.io_out [2] : \mchip.io_out [3]);
	assign _069_ = (io_in[4] ? _043_ : _068_);
	assign _070_ = ~(_069_ & _032_);
	assign _071_ = _031_ & ~_070_;
	assign _072_ = \mchip.io_out [2] & ~_065_;
	assign _073_ = _062_ & ~_066_;
	assign _074_ = ~(_073_ | _072_);
	assign _075_ = _063_ & ~io_in[5];
	assign _076_ = ~(_075_ | _049_);
	assign _077_ = _076_ ^ \mchip.io_out [3];
	assign _078_ = _077_ ^ _074_;
	assign _095_[3] = (_038_ ? _071_ : _078_);
	assign _079_ = ~_031_;
	assign _080_ = (io_in[3] ? \mchip.io_out [3] : \mchip.io_out [4]);
	assign _081_ = (io_in[4] ? _055_ : _080_);
	assign _082_ = (io_in[5] ? _034_ : _081_);
	assign _083_ = _082_ & ~_079_;
	assign _084_ = \mchip.io_out [3] & ~_076_;
	assign _085_ = _072_ & ~_077_;
	assign _086_ = _085_ | _084_;
	assign _087_ = _077_ | _066_;
	assign _088_ = _062_ & ~_087_;
	assign _089_ = _088_ | _086_;
	assign _090_ = _076_ ^ \mchip.io_out [4];
	assign _091_ = ~(_090_ ^ _089_);
	assign _095_[4] = (_038_ ? _083_ : _091_);
	assign _092_ = (io_in[3] ? \mchip.io_out [4] : \mchip.io_out [5]);
	assign _093_ = (io_in[4] ? _068_ : _092_);
	assign _094_ = (io_in[5] ? _044_ : _093_);
	assign _001_ = _094_ & ~_079_;
	assign _002_ = \mchip.io_out [4] & ~_076_;
	assign _003_ = _089_ & ~_090_;
	assign _004_ = ~(_003_ | _002_);
	assign _005_ = _076_ ^ \mchip.io_out [5];
	assign _006_ = _005_ ^ _004_;
	assign _095_[5] = (_038_ ? _001_ : _006_);
	assign _007_ = (io_in[3] ? \mchip.io_out [5] : \mchip.io_out [6]);
	assign _008_ = (io_in[4] ? _080_ : _007_);
	assign _009_ = (io_in[5] ? _056_ : _008_);
	assign _010_ = _009_ & ~_079_;
	assign _011_ = \mchip.io_out [5] & ~_076_;
	assign _012_ = _002_ & ~_005_;
	assign _013_ = _012_ | _011_;
	assign _014_ = _005_ | _090_;
	assign _015_ = _089_ & ~_014_;
	assign _016_ = _015_ | _013_;
	assign _017_ = ~(_076_ ^ \mchip.io_out [6]);
	assign _018_ = _017_ ^ _016_;
	assign _095_[6] = (_038_ ? _010_ : _018_);
	assign _019_ = (io_in[3] ? \mchip.io_out [6] : \mchip.io_out [7]);
	assign _020_ = (io_in[4] ? _092_ : _019_);
	assign _021_ = (io_in[5] ? _069_ : _020_);
	assign _022_ = _021_ & _031_;
	assign _023_ = \mchip.io_out [6] & ~_076_;
	assign _024_ = _017_ & _016_;
	assign _025_ = _024_ | _023_;
	assign _026_ = ~(_076_ ^ \mchip.io_out [7]);
	assign _027_ = _026_ ^ _025_;
	assign _095_[7] = (_038_ ? _022_ : _027_);
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.io_out [0] <= 1'h0;
		else if (\mchip.enable )
			\mchip.io_out [0] <= _095_[0];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.io_out [1] <= 1'h0;
		else if (\mchip.enable )
			\mchip.io_out [1] <= _095_[1];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.io_out [2] <= 1'h0;
		else if (\mchip.enable )
			\mchip.io_out [2] <= _095_[2];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.state  <= 1'h0;
		else
			\mchip.state  <= io_in[2];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.io_out [3] <= 1'h0;
		else if (_000_)
			\mchip.io_out [3] <= _095_[3];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.io_out [4] <= 1'h0;
		else if (_000_)
			\mchip.io_out [4] <= _095_[4];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.io_out [5] <= 1'h0;
		else if (_000_)
			\mchip.io_out [5] <= _095_[5];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.io_out [6] <= 1'h0;
		else if (_000_)
			\mchip.io_out [6] <= _095_[6];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.io_out [7] <= 1'h0;
		else if (_000_)
			\mchip.io_out [7] <= _095_[7];
	assign io_out = {6'h00, \mchip.io_out };
	assign \mchip.arithOp  = io_in[7:6];
	assign \mchip.clock  = io_in[0];
	assign \mchip.en  = io_in[2];
	assign \mchip.in  = io_in[5:3];
	assign \mchip.io_in  = io_in[7:0];
	assign \mchip.nextState  = io_in[2];
	assign \mchip.reset  = io_in[1];
endmodule
module d38_jxlu_pwm (
	io_in,
	io_out
);
	wire _000_;
	wire _001_;
	wire _002_;
	wire _003_;
	wire _004_;
	wire _005_;
	wire _006_;
	wire _007_;
	wire _008_;
	wire _009_;
	wire _010_;
	wire _011_;
	wire _012_;
	wire _013_;
	wire _014_;
	wire _015_;
	wire _016_;
	wire _017_;
	wire _018_;
	wire _019_;
	wire _020_;
	wire _021_;
	wire _022_;
	wire _023_;
	wire _024_;
	wire _025_;
	wire _026_;
	wire _027_;
	wire _028_;
	wire _029_;
	wire _030_;
	wire _031_;
	wire _032_;
	wire _033_;
	wire _034_;
	wire _035_;
	wire _036_;
	wire _037_;
	wire _038_;
	wire _039_;
	wire _040_;
	wire _041_;
	wire _042_;
	wire [5:0] _043_;
	wire [5:0] _044_;
	wire [5:0] _045_;
	input wire [13:0] io_in;
	output wire [13:0] io_out;
	wire [7:0] \mchip.io_in ;
	wire [7:0] \mchip.io_out ;
	reg [5:0] \mchip.pwm.active_duty ;
	wire \mchip.pwm.clk ;
	reg [5:0] \mchip.pwm.counter ;
	wire [5:0] \mchip.pwm.duty ;
	reg \mchip.pwm.pwm_signal ;
	wire \mchip.pwm.reset ;
	assign _002_ = \mchip.pwm.counter [0] & ~\mchip.pwm.counter [1];
	assign _003_ = \mchip.pwm.counter [2] | \mchip.pwm.counter [3];
	assign _004_ = _002_ & ~_003_;
	assign _005_ = ~(\mchip.pwm.counter [5] & \mchip.pwm.counter [4]);
	assign _006_ = _004_ & ~_005_;
	assign _000_ = _006_ | io_in[1];
	assign _044_[0] = ~\mchip.pwm.counter [0];
	assign _007_ = ~(\mchip.pwm.active_duty [0] ^ \mchip.pwm.counter [0]);
	assign _008_ = ~(\mchip.pwm.active_duty [1] ^ \mchip.pwm.counter [1]);
	assign _009_ = _008_ & _007_;
	assign _010_ = ~(\mchip.pwm.active_duty [3] ^ \mchip.pwm.counter [3]);
	assign _011_ = \mchip.pwm.active_duty [2] ^ \mchip.pwm.counter [2];
	assign _012_ = _010_ & ~_011_;
	assign _013_ = _012_ & _009_;
	assign _014_ = ~(\mchip.pwm.active_duty [5] ^ \mchip.pwm.counter [5]);
	assign _015_ = \mchip.pwm.active_duty [4] ^ \mchip.pwm.counter [4];
	assign _016_ = _014_ & ~_015_;
	assign _017_ = ~(_016_ & _013_);
	assign _018_ = \mchip.pwm.active_duty [3] | ~\mchip.pwm.counter [3];
	assign _019_ = \mchip.pwm.active_duty [2] | ~\mchip.pwm.counter [2];
	assign _020_ = _010_ & ~_019_;
	assign _021_ = _018_ & ~_020_;
	assign _022_ = \mchip.pwm.active_duty [1] | ~\mchip.pwm.counter [1];
	assign _023_ = \mchip.pwm.active_duty [0] & ~\mchip.pwm.counter [0];
	assign _024_ = _008_ & ~_023_;
	assign _025_ = _022_ & ~_024_;
	assign _026_ = _012_ & ~_025_;
	assign _027_ = _021_ & ~_026_;
	assign _028_ = _016_ & ~_027_;
	assign _029_ = \mchip.pwm.active_duty [4] | ~\mchip.pwm.counter [4];
	assign _030_ = _014_ & ~_029_;
	assign _031_ = \mchip.pwm.counter [5] & ~\mchip.pwm.active_duty [5];
	assign _032_ = _031_ | _030_;
	assign _033_ = _032_ | _028_;
	assign _001_ = _017_ & ~_033_;
	assign _045_[1] = \mchip.pwm.counter [1] ^ \mchip.pwm.counter [0];
	assign _034_ = ~(\mchip.pwm.counter [1] & \mchip.pwm.counter [0]);
	assign _045_[2] = ~(_034_ ^ \mchip.pwm.counter [2]);
	assign _035_ = \mchip.pwm.counter [2] & ~_034_;
	assign _045_[3] = _035_ ^ \mchip.pwm.counter [3];
	assign _036_ = ~(\mchip.pwm.counter [2] & \mchip.pwm.counter [3]);
	assign _037_ = _036_ | _034_;
	assign _045_[4] = ~(_037_ ^ \mchip.pwm.counter [4]);
	assign _038_ = \mchip.pwm.counter [4] & ~_037_;
	assign _045_[5] = _038_ ^ \mchip.pwm.counter [5];
	assign _039_ = ~(io_in[6] & io_in[7]);
	assign _040_ = ~(io_in[2] & io_in[3]);
	assign _041_ = io_in[4] | io_in[5];
	assign _042_ = _040_ & ~_041_;
	assign _043_[5] = _042_ | _039_;
	always @(posedge io_in[0])
		if (_000_)
			\mchip.pwm.counter [0] <= 1'h0;
		else
			\mchip.pwm.counter [0] <= _044_[0];
	always @(posedge io_in[0])
		if (_000_)
			\mchip.pwm.counter [1] <= 1'h0;
		else
			\mchip.pwm.counter [1] <= _045_[1];
	always @(posedge io_in[0])
		if (_000_)
			\mchip.pwm.counter [2] <= 1'h0;
		else
			\mchip.pwm.counter [2] <= _045_[2];
	always @(posedge io_in[0])
		if (_000_)
			\mchip.pwm.counter [3] <= 1'h0;
		else
			\mchip.pwm.counter [3] <= _045_[3];
	always @(posedge io_in[0])
		if (_000_)
			\mchip.pwm.counter [4] <= 1'h0;
		else
			\mchip.pwm.counter [4] <= _045_[4];
	always @(posedge io_in[0])
		if (_000_)
			\mchip.pwm.counter [5] <= 1'h0;
		else
			\mchip.pwm.counter [5] <= _045_[5];
	always @(posedge io_in[0])
		if (!io_in[1])
			\mchip.pwm.pwm_signal  <= _001_;
	always @(posedge io_in[0])
		if (io_in[1])
			if (!_043_[5])
				\mchip.pwm.active_duty [0] <= 1'h0;
			else
				\mchip.pwm.active_duty [0] <= io_in[2];
	always @(posedge io_in[0])
		if (io_in[1])
			if (!_043_[5])
				\mchip.pwm.active_duty [1] <= 1'h1;
			else
				\mchip.pwm.active_duty [1] <= io_in[3];
	always @(posedge io_in[0])
		if (io_in[1])
			if (!_043_[5])
				\mchip.pwm.active_duty [2] <= 1'h0;
			else
				\mchip.pwm.active_duty [2] <= io_in[4];
	always @(posedge io_in[0])
		if (io_in[1])
			if (!_043_[5])
				\mchip.pwm.active_duty [3] <= 1'h0;
			else
				\mchip.pwm.active_duty [3] <= io_in[5];
	always @(posedge io_in[0])
		if (io_in[1])
			if (!_043_[5])
				\mchip.pwm.active_duty [4] <= 1'h1;
			else
				\mchip.pwm.active_duty [4] <= io_in[6];
	always @(posedge io_in[0])
		if (io_in[1])
			if (!_043_[5])
				\mchip.pwm.active_duty [5] <= 1'h1;
			else
				\mchip.pwm.active_duty [5] <= io_in[7];
	assign _043_[4:0] = 5'h00;
	assign _044_[5:1] = \mchip.pwm.counter [5:1];
	assign _045_[0] = _044_[0];
	assign io_out = {13'h0000, \mchip.pwm.pwm_signal };
	assign \mchip.io_in  = io_in[7:0];
	assign \mchip.io_out  = {7'h00, \mchip.pwm.pwm_signal };
	assign \mchip.pwm.clk  = io_in[0];
	assign \mchip.pwm.duty  = io_in[7:2];
	assign \mchip.pwm.reset  = io_in[1];
endmodule
module d39_oonyeado_sevenseg (
	io_in,
	io_out
);
	wire _000_;
	wire _001_;
	wire _002_;
	wire _003_;
	wire _004_;
	wire _005_;
	wire _006_;
	wire _007_;
	wire _008_;
	wire _009_;
	wire _010_;
	wire _011_;
	wire _012_;
	wire _013_;
	wire _014_;
	wire _015_;
	wire _016_;
	wire _017_;
	wire _018_;
	wire _019_;
	wire _020_;
	wire _021_;
	wire _022_;
	wire _023_;
	wire _024_;
	wire _025_;
	wire _026_;
	wire _027_;
	wire _028_;
	wire _029_;
	wire _030_;
	wire _031_;
	wire _032_;
	wire _033_;
	wire _034_;
	wire _035_;
	wire _036_;
	wire _037_;
	wire _038_;
	wire _039_;
	wire _040_;
	wire _041_;
	wire _042_;
	wire _043_;
	wire _044_;
	wire _045_;
	wire _046_;
	wire _047_;
	wire _048_;
	wire _049_;
	input wire [13:0] io_in;
	output wire [13:0] io_out;
	wire \mchip.gate1.b ;
	wire \mchip.gate11.out ;
	wire \mchip.gate15.out ;
	wire \mchip.gate19.out ;
	wire \mchip.gate22.out ;
	wire \mchip.gate26.out ;
	wire \mchip.gate30.out ;
	wire \mchip.gate32.out ;
	wire \mchip.gate37.a ;
	wire \mchip.gate37.b ;
	wire \mchip.gate39.a ;
	wire \mchip.gate40.b ;
	wire \mchip.gate41.a ;
	wire \mchip.gate41.b ;
	wire \mchip.gate43.b ;
	wire \mchip.gate45.a ;
	wire \mchip.gate46.b ;
	wire \mchip.gate47.b ;
	wire \mchip.gate48.b ;
	wire \mchip.gate49.b ;
	wire \mchip.gate5.in ;
	wire \mchip.gate50.b ;
	wire \mchip.gate53.a ;
	wire \mchip.gate55.a ;
	wire \mchip.gate55.b ;
	wire \mchip.gate56.a ;
	wire \mchip.gate56.b ;
	wire \mchip.gate58.b ;
	wire \mchip.gate59.a ;
	wire \mchip.gate60.a ;
	wire \mchip.gate60.b ;
	wire \mchip.gate64.b ;
	wire \mchip.gate65.b ;
	wire \mchip.gate66.b ;
	wire \mchip.gate67.a ;
	wire \mchip.gate68.a ;
	wire \mchip.gate69.a ;
	wire \mchip.gate7.in ;
	wire \mchip.gate72.a ;
	wire \mchip.gate73.a ;
	wire \mchip.gate74.a ;
	wire \mchip.gate74.b ;
	wire \mchip.gate75.a ;
	wire \mchip.gate76.a ;
	wire \mchip.gate76.b ;
	wire \mchip.gate77.b ;
	wire \mchip.gate78.a ;
	wire \mchip.gate8.in ;
	wire \mchip.gate9.in ;
	wire [7:0] \mchip.io_in ;
	wire [7:0] \mchip.io_out ;
	wire \mchip.net1 ;
	wire \mchip.net10 ;
	wire \mchip.net11 ;
	wire \mchip.net12 ;
	wire \mchip.net2 ;
	wire \mchip.net3 ;
	wire \mchip.net4 ;
	wire \mchip.net5 ;
	wire \mchip.net6 ;
	wire \mchip.net7 ;
	wire \mchip.net8 ;
	wire \mchip.net84 ;
	wire \mchip.net9 ;
	assign _000_ = ~(io_in[5] & io_in[6]);
	assign _001_ = io_in[4] | ~io_in[7];
	assign _002_ = ~(_001_ & _000_);
	assign _003_ = io_in[5] & ~io_in[7];
	assign _004_ = _003_ | _002_;
	assign _005_ = ~(io_in[4] | io_in[6]);
	assign _006_ = io_in[7] | ~io_in[6];
	assign _007_ = io_in[4] & ~_006_;
	assign _008_ = io_in[7] & ~io_in[6];
	assign _009_ = _008_ & ~io_in[5];
	assign _010_ = _009_ | _007_;
	assign _011_ = _010_ | _005_;
	assign \mchip.gate32.out  = _011_ | _004_;
	assign _012_ = _008_ | ~_006_;
	assign _013_ = io_in[4] & ~io_in[5];
	assign _014_ = _013_ | _012_;
	assign _015_ = io_in[4] & ~io_in[7];
	assign _016_ = ~(io_in[5] | io_in[7]);
	assign _017_ = _016_ | _015_;
	assign \mchip.gate30.out  = _017_ | _014_;
	assign _018_ = ~(io_in[5] | io_in[6]);
	assign _019_ = _018_ | _005_;
	assign _020_ = ~io_in[4];
	assign _021_ = io_in[7] & ~io_in[5];
	assign _022_ = _021_ & ~_020_;
	assign _023_ = _022_ | _019_;
	assign _024_ = (io_in[4] ? _003_ : _016_);
	assign \mchip.gate26.out  = _024_ | _023_;
	assign _025_ = io_in[5] & ~io_in[4];
	assign _026_ = io_in[5] & ~io_in[6];
	assign _027_ = _026_ | _025_;
	assign _028_ = io_in[4] & io_in[7];
	assign _029_ = _028_ | _027_;
	assign _030_ = ~(_006_ | io_in[5]);
	assign _031_ = _030_ | _008_;
	assign \mchip.gate22.out  = _031_ | _029_;
	assign _032_ = _025_ | _005_;
	assign _033_ = io_in[6] & io_in[7];
	assign _034_ = io_in[5] & io_in[7];
	assign _035_ = _034_ | _033_;
	assign \mchip.gate19.out  = _035_ | _032_;
	assign _036_ = _034_ | _008_;
	assign _037_ = io_in[6] & ~io_in[4];
	assign _038_ = _037_ | _036_;
	assign _039_ = ~(io_in[4] | io_in[5]);
	assign _040_ = _039_ | _030_;
	assign \mchip.gate15.out  = _040_ | _038_;
	assign _041_ = _020_ & ~_000_;
	assign _042_ = _041_ | _021_;
	assign _043_ = io_in[5] | ~io_in[6];
	assign _044_ = io_in[4] & ~_043_;
	assign _045_ = _044_ | _042_;
	assign _046_ = io_in[4] & io_in[5];
	assign _047_ = _046_ & ~io_in[6];
	assign _048_ = _005_ & ~io_in[7];
	assign _049_ = _048_ | _047_;
	assign \mchip.gate11.out  = _049_ | _045_;
	assign io_out = {6'h00, \mchip.gate22.out , \mchip.gate15.out , \mchip.gate19.out , \mchip.gate11.out , \mchip.gate30.out , \mchip.gate26.out , \mchip.gate32.out , 1'h0};
	assign \mchip.gate1.b  = io_in[6];
	assign \mchip.gate37.a  = io_in[4];
	assign \mchip.gate37.b  = io_in[5];
	assign \mchip.gate39.a  = io_in[6];
	assign \mchip.gate40.b  = io_in[4];
	assign \mchip.gate41.a  = io_in[6];
	assign \mchip.gate41.b  = io_in[5];
	assign \mchip.gate43.b  = io_in[6];
	assign \mchip.gate45.a  = io_in[7];
	assign \mchip.gate46.b  = io_in[4];
	assign \mchip.gate47.b  = io_in[5];
	assign \mchip.gate48.b  = io_in[4];
	assign \mchip.gate49.b  = io_in[6];
	assign \mchip.gate5.in  = io_in[7];
	assign \mchip.gate50.b  = io_in[4];
	assign \mchip.gate53.a  = io_in[7];
	assign \mchip.gate55.a  = io_in[7];
	assign \mchip.gate55.b  = io_in[5];
	assign \mchip.gate56.a  = io_in[7];
	assign \mchip.gate56.b  = io_in[6];
	assign \mchip.gate58.b  = io_in[5];
	assign \mchip.gate59.a  = io_in[7];
	assign \mchip.gate60.a  = io_in[6];
	assign \mchip.gate60.b  = io_in[5];
	assign \mchip.gate64.b  = io_in[4];
	assign \mchip.gate65.b  = io_in[4];
	assign \mchip.gate66.b  = io_in[6];
	assign \mchip.gate67.a  = io_in[7];
	assign \mchip.gate68.a  = io_in[5];
	assign \mchip.gate69.a  = io_in[7];
	assign \mchip.gate7.in  = io_in[6];
	assign \mchip.gate72.a  = io_in[6];
	assign \mchip.gate73.a  = io_in[7];
	assign \mchip.gate74.a  = io_in[7];
	assign \mchip.gate74.b  = io_in[5];
	assign \mchip.gate75.a  = io_in[7];
	assign \mchip.gate76.a  = io_in[7];
	assign \mchip.gate76.b  = io_in[4];
	assign \mchip.gate77.b  = io_in[5];
	assign \mchip.gate78.a  = io_in[5];
	assign \mchip.gate8.in  = io_in[5];
	assign \mchip.gate9.in  = io_in[4];
	assign \mchip.io_in  = io_in[7:0];
	assign \mchip.io_out  = {\mchip.gate22.out , \mchip.gate15.out , \mchip.gate19.out , \mchip.gate11.out , \mchip.gate30.out , \mchip.gate26.out , \mchip.gate32.out , 1'h0};
	assign \mchip.net1  = io_in[4];
	assign \mchip.net10  = \mchip.gate15.out ;
	assign \mchip.net11  = \mchip.gate22.out ;
	assign \mchip.net12  = 1'h1;
	assign \mchip.net2  = io_in[5];
	assign \mchip.net3  = io_in[6];
	assign \mchip.net4  = io_in[7];
	assign \mchip.net5  = \mchip.gate32.out ;
	assign \mchip.net6  = \mchip.gate26.out ;
	assign \mchip.net7  = \mchip.gate30.out ;
	assign \mchip.net8  = \mchip.gate11.out ;
	assign \mchip.net84  = 1'h0;
	assign \mchip.net9  = \mchip.gate19.out ;
endmodule
module d40_jrecta_asyncfifo (
	io_in,
	io_out
);
	wire _000_;
	wire _001_;
	wire _002_;
	wire _003_;
	wire _004_;
	wire _005_;
	wire _006_;
	wire _007_;
	wire _008_;
	wire _009_;
	wire _010_;
	wire _011_;
	wire _012_;
	wire _013_;
	wire _014_;
	wire _015_;
	wire _016_;
	wire _017_;
	wire _018_;
	wire _019_;
	wire _020_;
	wire _021_;
	wire _022_;
	wire _023_;
	wire _024_;
	wire _025_;
	wire _026_;
	wire _027_;
	wire _028_;
	wire _029_;
	wire _030_;
	wire _031_;
	wire _032_;
	wire _033_;
	wire _034_;
	wire _035_;
	wire _036_;
	wire _037_;
	wire _038_;
	wire _039_;
	wire _040_;
	wire _041_;
	wire _042_;
	wire _043_;
	wire _044_;
	wire _045_;
	wire _046_;
	wire _047_;
	wire _048_;
	wire _049_;
	wire _050_;
	wire _051_;
	wire _052_;
	wire _053_;
	wire _054_;
	input wire [13:0] io_in;
	output wire [13:0] io_out;
	wire [7:0] \mchip.io_in ;
	wire [7:0] \mchip.io_out ;
	wire \mchip.top.backend.empty ;
	wire \mchip.top.backend.rclk ;
	wire \mchip.top.backend.re ;
	wire [3:0] \mchip.top.backend.rptr ;
	wire [3:0] \mchip.top.backend.rptr_b2g.binary ;
	wire [3:0] \mchip.top.backend.rptr_b2g.gray ;
	wire [3:0] \mchip.top.backend.rptr_gray ;
	wire \mchip.top.backend.rptr_reg.clk ;
	wire [3:0] \mchip.top.backend.rptr_reg.d ;
	wire \mchip.top.backend.rptr_reg.en ;
	reg [3:0] \mchip.top.backend.rptr_reg.q ;
	wire \mchip.top.backend.rptr_reg.rst ;
	wire \mchip.top.backend.rst ;
	wire [3:0] \mchip.top.backend.wptr_gray ;
	wire [3:0] \mchip.top.backend.wptr_gray1 ;
	wire [3:0] \mchip.top.backend.wptr_gray2 ;
	wire \mchip.top.backend.wptr_gray_sync.clk ;
	wire [7:0] \mchip.top.backend.wptr_gray_sync.d ;
	wire \mchip.top.backend.wptr_gray_sync.en ;
	reg [7:0] \mchip.top.backend.wptr_gray_sync.q ;
	wire \mchip.top.backend.wptr_gray_sync.rst ;
	reg [2:0] \mchip.top.data[0] ;
	reg [2:0] \mchip.top.data[1] ;
	reg [2:0] \mchip.top.data[2] ;
	reg [2:0] \mchip.top.data[3] ;
	reg [2:0] \mchip.top.data[4] ;
	reg [2:0] \mchip.top.data[5] ;
	reg [2:0] \mchip.top.data[6] ;
	reg [2:0] \mchip.top.data[7] ;
	wire \mchip.top.empty ;
	wire \mchip.top.frontend.full ;
	wire [3:0] \mchip.top.frontend.rptr_gray ;
	wire [3:0] \mchip.top.frontend.rptr_gray1 ;
	wire [3:0] \mchip.top.frontend.rptr_gray2 ;
	wire \mchip.top.frontend.rptr_gray_sync.clk ;
	wire [7:0] \mchip.top.frontend.rptr_gray_sync.d ;
	wire \mchip.top.frontend.rptr_gray_sync.en ;
	reg [7:0] \mchip.top.frontend.rptr_gray_sync.q ;
	wire \mchip.top.frontend.rptr_gray_sync.rst ;
	wire \mchip.top.frontend.rst ;
	wire \mchip.top.frontend.wclk ;
	wire \mchip.top.frontend.we ;
	wire [3:0] \mchip.top.frontend.wptr ;
	wire [3:0] \mchip.top.frontend.wptr_b2g.binary ;
	wire [3:0] \mchip.top.frontend.wptr_b2g.gray ;
	wire [3:0] \mchip.top.frontend.wptr_gray ;
	wire \mchip.top.frontend.wptr_reg.clk ;
	wire [3:0] \mchip.top.frontend.wptr_reg.d ;
	wire \mchip.top.frontend.wptr_reg.en ;
	reg [3:0] \mchip.top.frontend.wptr_reg.q ;
	wire \mchip.top.frontend.wptr_reg.rst ;
	wire \mchip.top.full ;
	wire \mchip.top.rclk ;
	wire [2:0] \mchip.top.rdata ;
	wire \mchip.top.re ;
	wire [3:0] \mchip.top.rptr ;
	wire [3:0] \mchip.top.rptr_gray ;
	wire \mchip.top.rst ;
	wire \mchip.top.wclk ;
	wire [2:0] \mchip.top.wdata ;
	wire \mchip.top.we ;
	wire [3:0] \mchip.top.wptr ;
	wire [3:0] \mchip.top.wptr_gray ;
	assign \mchip.top.frontend.wptr_reg.d [0] = ~\mchip.top.frontend.wptr_reg.q [0];
	assign \mchip.top.backend.rptr_reg.d [0] = ~\mchip.top.backend.rptr_reg.q [0];
	assign \mchip.top.backend.rptr_gray [0] = \mchip.top.backend.rptr_reg.q [1] ^ \mchip.top.backend.rptr_reg.q [0];
	assign _036_ = ~(\mchip.top.backend.rptr_gray [0] ^ \mchip.top.backend.wptr_gray_sync.q [0]);
	assign \mchip.top.backend.rptr_gray [1] = \mchip.top.backend.rptr_reg.q [2] ^ \mchip.top.backend.rptr_reg.q [1];
	assign _037_ = \mchip.top.backend.rptr_gray [1] ^ \mchip.top.backend.wptr_gray_sync.q [1];
	assign _038_ = _036_ & ~_037_;
	assign _039_ = \mchip.top.backend.wptr_gray_sync.q [3] ^ \mchip.top.backend.rptr_reg.q [3];
	assign \mchip.top.backend.rptr_gray [2] = \mchip.top.backend.rptr_reg.q [3] ^ \mchip.top.backend.rptr_reg.q [2];
	assign _040_ = \mchip.top.backend.rptr_gray [2] ^ \mchip.top.backend.wptr_gray_sync.q [2];
	assign _041_ = _040_ | _039_;
	assign \mchip.top.backend.empty  = _038_ & ~_041_;
	assign \mchip.top.frontend.wptr_gray [2] = \mchip.top.frontend.wptr_reg.q [2] ^ \mchip.top.frontend.wptr_reg.q [3];
	assign _042_ = \mchip.top.frontend.wptr_gray [2] ^ \mchip.top.frontend.rptr_gray_sync.q [2];
	assign _043_ = ~(\mchip.top.frontend.rptr_gray_sync.q [3] ^ \mchip.top.frontend.wptr_reg.q [3]);
	assign _044_ = _042_ & ~_043_;
	assign \mchip.top.frontend.wptr_gray [1] = \mchip.top.frontend.wptr_reg.q [1] ^ \mchip.top.frontend.wptr_reg.q [2];
	assign _045_ = \mchip.top.frontend.wptr_gray [1] ^ \mchip.top.frontend.rptr_gray_sync.q [1];
	assign \mchip.top.frontend.wptr_gray [0] = \mchip.top.frontend.wptr_reg.q [1] ^ \mchip.top.frontend.wptr_reg.q [0];
	assign _046_ = \mchip.top.frontend.wptr_gray [0] ^ \mchip.top.frontend.rptr_gray_sync.q [0];
	assign _047_ = _046_ | _045_;
	assign \mchip.top.frontend.full  = _044_ & ~_047_;
	assign _048_ = ~\mchip.top.backend.rptr_reg.q [2];
	assign _049_ = (\mchip.top.backend.rptr_reg.q [0] ? \mchip.top.data[1] [0] : \mchip.top.data[0] [0]);
	assign _050_ = (\mchip.top.backend.rptr_reg.q [0] ? \mchip.top.data[3] [0] : \mchip.top.data[2] [0]);
	assign _051_ = (\mchip.top.backend.rptr_reg.q [1] ? _050_ : _049_);
	assign _052_ = (\mchip.top.backend.rptr_reg.q [0] ? \mchip.top.data[5] [0] : \mchip.top.data[4] [0]);
	assign _053_ = (\mchip.top.backend.rptr_reg.q [0] ? \mchip.top.data[7] [0] : \mchip.top.data[6] [0]);
	assign _054_ = (\mchip.top.backend.rptr_reg.q [1] ? _053_ : _052_);
	assign io_out[5] = (\mchip.top.backend.rptr_reg.q [2] ? _054_ : _051_);
	assign _008_ = (\mchip.top.backend.rptr_reg.q [0] ? \mchip.top.data[1] [1] : \mchip.top.data[0] [1]);
	assign _009_ = (\mchip.top.backend.rptr_reg.q [0] ? \mchip.top.data[3] [1] : \mchip.top.data[2] [1]);
	assign _010_ = (\mchip.top.backend.rptr_reg.q [1] ? _009_ : _008_);
	assign _011_ = (\mchip.top.backend.rptr_reg.q [0] ? \mchip.top.data[5] [1] : \mchip.top.data[4] [1]);
	assign _012_ = (\mchip.top.backend.rptr_reg.q [0] ? \mchip.top.data[7] [1] : \mchip.top.data[6] [1]);
	assign _013_ = (\mchip.top.backend.rptr_reg.q [1] ? _012_ : _011_);
	assign io_out[6] = (\mchip.top.backend.rptr_reg.q [2] ? _013_ : _010_);
	assign _014_ = (\mchip.top.backend.rptr_reg.q [0] ? \mchip.top.data[1] [2] : \mchip.top.data[0] [2]);
	assign _015_ = (\mchip.top.backend.rptr_reg.q [0] ? \mchip.top.data[3] [2] : \mchip.top.data[2] [2]);
	assign _016_ = (\mchip.top.backend.rptr_reg.q [1] ? _015_ : _014_);
	assign _017_ = (\mchip.top.backend.rptr_reg.q [0] ? \mchip.top.data[5] [2] : \mchip.top.data[4] [2]);
	assign _018_ = (\mchip.top.backend.rptr_reg.q [0] ? \mchip.top.data[7] [2] : \mchip.top.data[6] [2]);
	assign _019_ = (\mchip.top.backend.rptr_reg.q [1] ? _018_ : _017_);
	assign io_out[7] = (\mchip.top.backend.rptr_reg.q [2] ? _019_ : _016_);
	assign \mchip.top.frontend.wptr_reg.en  = io_in[3] & ~\mchip.top.frontend.full ;
	assign _020_ = \mchip.top.frontend.wptr_reg.q [2] | ~\mchip.top.frontend.wptr_reg.q [1];
	assign _021_ = _020_ | \mchip.top.frontend.wptr_reg.q [0];
	assign _002_ = \mchip.top.frontend.wptr_reg.en  & ~_021_;
	assign _022_ = _020_ | \mchip.top.frontend.wptr_reg.d [0];
	assign _003_ = \mchip.top.frontend.wptr_reg.en  & ~_022_;
	assign _023_ = \mchip.top.frontend.wptr_reg.q [1] | ~\mchip.top.frontend.wptr_reg.q [2];
	assign _024_ = _023_ | \mchip.top.frontend.wptr_reg.q [0];
	assign _004_ = \mchip.top.frontend.wptr_reg.en  & ~_024_;
	assign _025_ = _023_ | \mchip.top.frontend.wptr_reg.d [0];
	assign _005_ = \mchip.top.frontend.wptr_reg.en  & ~_025_;
	assign _026_ = ~(\mchip.top.frontend.wptr_reg.q [1] & \mchip.top.frontend.wptr_reg.q [2]);
	assign _027_ = _026_ | \mchip.top.frontend.wptr_reg.q [0];
	assign _006_ = \mchip.top.frontend.wptr_reg.en  & ~_027_;
	assign _028_ = _026_ | \mchip.top.frontend.wptr_reg.d [0];
	assign _007_ = \mchip.top.frontend.wptr_reg.en  & ~_028_;
	assign _029_ = \mchip.top.frontend.wptr_reg.q [1] | \mchip.top.frontend.wptr_reg.q [2];
	assign _030_ = _029_ | \mchip.top.frontend.wptr_reg.q [0];
	assign _000_ = \mchip.top.frontend.wptr_reg.en  & ~_030_;
	assign _031_ = _029_ | \mchip.top.frontend.wptr_reg.d [0];
	assign _001_ = \mchip.top.frontend.wptr_reg.en  & ~_031_;
	assign \mchip.top.backend.rptr_reg.en  = io_in[4] & ~\mchip.top.backend.empty ;
	assign _032_ = ~(\mchip.top.backend.rptr_reg.q [1] & \mchip.top.backend.rptr_reg.q [0]);
	assign \mchip.top.backend.rptr_reg.d [2] = _032_ ^ _048_;
	assign _033_ = \mchip.top.backend.rptr_reg.q [2] & ~_032_;
	assign \mchip.top.backend.rptr_reg.d [3] = _033_ ^ \mchip.top.backend.rptr_reg.q [3];
	assign _034_ = ~(\mchip.top.frontend.wptr_reg.q [1] & \mchip.top.frontend.wptr_reg.q [0]);
	assign \mchip.top.frontend.wptr_reg.d [2] = ~(_034_ ^ \mchip.top.frontend.wptr_reg.q [2]);
	assign _035_ = \mchip.top.frontend.wptr_reg.q [2] & ~_034_;
	assign \mchip.top.frontend.wptr_reg.d [3] = _035_ ^ \mchip.top.frontend.wptr_reg.q [3];
	always @(posedge io_in[0])
		if (_007_)
			\mchip.top.data[7] [0] <= io_in[5];
	always @(posedge io_in[0])
		if (_007_)
			\mchip.top.data[7] [1] <= io_in[6];
	always @(posedge io_in[0])
		if (_007_)
			\mchip.top.data[7] [2] <= io_in[7];
	always @(posedge io_in[0])
		if (_001_)
			\mchip.top.data[1] [0] <= io_in[5];
	always @(posedge io_in[0])
		if (_001_)
			\mchip.top.data[1] [1] <= io_in[6];
	always @(posedge io_in[0])
		if (_001_)
			\mchip.top.data[1] [2] <= io_in[7];
	always @(posedge io_in[0])
		if (io_in[2])
			\mchip.top.frontend.rptr_gray_sync.q [0] <= 1'h0;
		else
			\mchip.top.frontend.rptr_gray_sync.q [0] <= \mchip.top.frontend.rptr_gray_sync.q [4];
	always @(posedge io_in[0])
		if (io_in[2])
			\mchip.top.frontend.rptr_gray_sync.q [1] <= 1'h0;
		else
			\mchip.top.frontend.rptr_gray_sync.q [1] <= \mchip.top.frontend.rptr_gray_sync.q [5];
	always @(posedge io_in[0])
		if (io_in[2])
			\mchip.top.frontend.rptr_gray_sync.q [2] <= 1'h0;
		else
			\mchip.top.frontend.rptr_gray_sync.q [2] <= \mchip.top.frontend.rptr_gray_sync.q [6];
	always @(posedge io_in[0])
		if (io_in[2])
			\mchip.top.frontend.rptr_gray_sync.q [3] <= 1'h0;
		else
			\mchip.top.frontend.rptr_gray_sync.q [3] <= \mchip.top.frontend.rptr_gray_sync.q [7];
	always @(posedge io_in[0])
		if (io_in[2])
			\mchip.top.frontend.rptr_gray_sync.q [4] <= 1'h0;
		else
			\mchip.top.frontend.rptr_gray_sync.q [4] <= \mchip.top.backend.rptr_gray [0];
	always @(posedge io_in[0])
		if (io_in[2])
			\mchip.top.frontend.rptr_gray_sync.q [5] <= 1'h0;
		else
			\mchip.top.frontend.rptr_gray_sync.q [5] <= \mchip.top.backend.rptr_gray [1];
	always @(posedge io_in[0])
		if (io_in[2])
			\mchip.top.frontend.rptr_gray_sync.q [6] <= 1'h0;
		else
			\mchip.top.frontend.rptr_gray_sync.q [6] <= \mchip.top.backend.rptr_gray [2];
	always @(posedge io_in[0])
		if (io_in[2])
			\mchip.top.frontend.rptr_gray_sync.q [7] <= 1'h0;
		else
			\mchip.top.frontend.rptr_gray_sync.q [7] <= \mchip.top.backend.rptr_reg.q [3];
	always @(posedge io_in[0])
		if (_002_)
			\mchip.top.data[2] [0] <= io_in[5];
	always @(posedge io_in[0])
		if (_002_)
			\mchip.top.data[2] [1] <= io_in[6];
	always @(posedge io_in[0])
		if (_002_)
			\mchip.top.data[2] [2] <= io_in[7];
	always @(posedge io_in[0])
		if (_006_)
			\mchip.top.data[6] [0] <= io_in[5];
	always @(posedge io_in[0])
		if (_006_)
			\mchip.top.data[6] [1] <= io_in[6];
	always @(posedge io_in[0])
		if (_006_)
			\mchip.top.data[6] [2] <= io_in[7];
	always @(posedge io_in[0])
		if (_005_)
			\mchip.top.data[5] [0] <= io_in[5];
	always @(posedge io_in[0])
		if (_005_)
			\mchip.top.data[5] [1] <= io_in[6];
	always @(posedge io_in[0])
		if (_005_)
			\mchip.top.data[5] [2] <= io_in[7];
	always @(posedge io_in[0])
		if (_004_)
			\mchip.top.data[4] [0] <= io_in[5];
	always @(posedge io_in[0])
		if (_004_)
			\mchip.top.data[4] [1] <= io_in[6];
	always @(posedge io_in[0])
		if (_004_)
			\mchip.top.data[4] [2] <= io_in[7];
	always @(posedge io_in[0])
		if (_000_)
			\mchip.top.data[0] [0] <= io_in[5];
	always @(posedge io_in[0])
		if (_000_)
			\mchip.top.data[0] [1] <= io_in[6];
	always @(posedge io_in[0])
		if (_000_)
			\mchip.top.data[0] [2] <= io_in[7];
	always @(posedge io_in[1])
		if (io_in[2])
			\mchip.top.backend.wptr_gray_sync.q [0] <= 1'h0;
		else
			\mchip.top.backend.wptr_gray_sync.q [0] <= \mchip.top.backend.wptr_gray_sync.q [4];
	always @(posedge io_in[1])
		if (io_in[2])
			\mchip.top.backend.wptr_gray_sync.q [1] <= 1'h0;
		else
			\mchip.top.backend.wptr_gray_sync.q [1] <= \mchip.top.backend.wptr_gray_sync.q [5];
	always @(posedge io_in[1])
		if (io_in[2])
			\mchip.top.backend.wptr_gray_sync.q [2] <= 1'h0;
		else
			\mchip.top.backend.wptr_gray_sync.q [2] <= \mchip.top.backend.wptr_gray_sync.q [6];
	always @(posedge io_in[1])
		if (io_in[2])
			\mchip.top.backend.wptr_gray_sync.q [3] <= 1'h0;
		else
			\mchip.top.backend.wptr_gray_sync.q [3] <= \mchip.top.backend.wptr_gray_sync.q [7];
	always @(posedge io_in[1])
		if (io_in[2])
			\mchip.top.backend.wptr_gray_sync.q [4] <= 1'h0;
		else
			\mchip.top.backend.wptr_gray_sync.q [4] <= \mchip.top.frontend.wptr_gray [0];
	always @(posedge io_in[1])
		if (io_in[2])
			\mchip.top.backend.wptr_gray_sync.q [5] <= 1'h0;
		else
			\mchip.top.backend.wptr_gray_sync.q [5] <= \mchip.top.frontend.wptr_gray [1];
	always @(posedge io_in[1])
		if (io_in[2])
			\mchip.top.backend.wptr_gray_sync.q [6] <= 1'h0;
		else
			\mchip.top.backend.wptr_gray_sync.q [6] <= \mchip.top.frontend.wptr_gray [2];
	always @(posedge io_in[1])
		if (io_in[2])
			\mchip.top.backend.wptr_gray_sync.q [7] <= 1'h0;
		else
			\mchip.top.backend.wptr_gray_sync.q [7] <= \mchip.top.frontend.wptr_reg.q [3];
	always @(posedge io_in[0])
		if (_003_)
			\mchip.top.data[3] [0] <= io_in[5];
	always @(posedge io_in[0])
		if (_003_)
			\mchip.top.data[3] [1] <= io_in[6];
	always @(posedge io_in[0])
		if (_003_)
			\mchip.top.data[3] [2] <= io_in[7];
	always @(posedge io_in[0])
		if (io_in[2])
			\mchip.top.frontend.wptr_reg.q [0] <= 1'h0;
		else if (\mchip.top.frontend.wptr_reg.en )
			\mchip.top.frontend.wptr_reg.q [0] <= \mchip.top.frontend.wptr_reg.d [0];
	always @(posedge io_in[0])
		if (io_in[2])
			\mchip.top.frontend.wptr_reg.q [1] <= 1'h0;
		else if (\mchip.top.frontend.wptr_reg.en )
			\mchip.top.frontend.wptr_reg.q [1] <= \mchip.top.frontend.wptr_gray [0];
	always @(posedge io_in[0])
		if (io_in[2])
			\mchip.top.frontend.wptr_reg.q [2] <= 1'h0;
		else if (\mchip.top.frontend.wptr_reg.en )
			\mchip.top.frontend.wptr_reg.q [2] <= \mchip.top.frontend.wptr_reg.d [2];
	always @(posedge io_in[0])
		if (io_in[2])
			\mchip.top.frontend.wptr_reg.q [3] <= 1'h0;
		else if (\mchip.top.frontend.wptr_reg.en )
			\mchip.top.frontend.wptr_reg.q [3] <= \mchip.top.frontend.wptr_reg.d [3];
	always @(posedge io_in[1])
		if (io_in[2])
			\mchip.top.backend.rptr_reg.q [0] <= 1'h0;
		else if (\mchip.top.backend.rptr_reg.en )
			\mchip.top.backend.rptr_reg.q [0] <= \mchip.top.backend.rptr_reg.d [0];
	always @(posedge io_in[1])
		if (io_in[2])
			\mchip.top.backend.rptr_reg.q [1] <= 1'h0;
		else if (\mchip.top.backend.rptr_reg.en )
			\mchip.top.backend.rptr_reg.q [1] <= \mchip.top.backend.rptr_gray [0];
	always @(posedge io_in[1])
		if (io_in[2])
			\mchip.top.backend.rptr_reg.q [2] <= 1'h0;
		else if (\mchip.top.backend.rptr_reg.en )
			\mchip.top.backend.rptr_reg.q [2] <= \mchip.top.backend.rptr_reg.d [2];
	always @(posedge io_in[1])
		if (io_in[2])
			\mchip.top.backend.rptr_reg.q [3] <= 1'h0;
		else if (\mchip.top.backend.rptr_reg.en )
			\mchip.top.backend.rptr_reg.q [3] <= \mchip.top.backend.rptr_reg.d [3];
	assign {io_out[13:8], io_out[4:0]} = {6'h00, \mchip.top.backend.empty , \mchip.top.frontend.full , 3'h0};
	assign \mchip.io_in  = io_in[7:0];
	assign \mchip.io_out  = {io_out[7:5], \mchip.top.backend.empty , \mchip.top.frontend.full , 3'h0};
	assign \mchip.top.backend.rclk  = io_in[1];
	assign \mchip.top.backend.re  = io_in[4];
	assign \mchip.top.backend.rptr  = \mchip.top.backend.rptr_reg.q ;
	assign \mchip.top.backend.rptr_b2g.binary  = \mchip.top.backend.rptr_reg.q ;
	assign \mchip.top.backend.rptr_b2g.gray  = {\mchip.top.backend.rptr_reg.q [3], \mchip.top.backend.rptr_gray [2:0]};
	assign \mchip.top.backend.rptr_gray [3] = \mchip.top.backend.rptr_reg.q [3];
	assign \mchip.top.backend.rptr_reg.clk  = io_in[1];
	assign \mchip.top.backend.rptr_reg.d [1] = \mchip.top.backend.rptr_gray [0];
	assign \mchip.top.backend.rptr_reg.rst  = io_in[2];
	assign \mchip.top.backend.rst  = io_in[2];
	assign \mchip.top.backend.wptr_gray  = {\mchip.top.frontend.wptr_reg.q [3], \mchip.top.frontend.wptr_gray [2:0]};
	assign \mchip.top.backend.wptr_gray1  = \mchip.top.backend.wptr_gray_sync.q [7:4];
	assign \mchip.top.backend.wptr_gray2  = \mchip.top.backend.wptr_gray_sync.q [3:0];
	assign \mchip.top.backend.wptr_gray_sync.clk  = io_in[1];
	assign \mchip.top.backend.wptr_gray_sync.d  = {\mchip.top.frontend.wptr_reg.q [3], \mchip.top.frontend.wptr_gray [2:0], \mchip.top.backend.wptr_gray_sync.q [7:4]};
	assign \mchip.top.backend.wptr_gray_sync.en  = 1'h1;
	assign \mchip.top.backend.wptr_gray_sync.rst  = io_in[2];
	assign \mchip.top.empty  = \mchip.top.backend.empty ;
	assign \mchip.top.frontend.rptr_gray  = {\mchip.top.backend.rptr_reg.q [3], \mchip.top.backend.rptr_gray [2:0]};
	assign \mchip.top.frontend.rptr_gray1  = \mchip.top.frontend.rptr_gray_sync.q [7:4];
	assign \mchip.top.frontend.rptr_gray2  = \mchip.top.frontend.rptr_gray_sync.q [3:0];
	assign \mchip.top.frontend.rptr_gray_sync.clk  = io_in[0];
	assign \mchip.top.frontend.rptr_gray_sync.d  = {\mchip.top.backend.rptr_reg.q [3], \mchip.top.backend.rptr_gray [2:0], \mchip.top.frontend.rptr_gray_sync.q [7:4]};
	assign \mchip.top.frontend.rptr_gray_sync.en  = 1'h1;
	assign \mchip.top.frontend.rptr_gray_sync.rst  = io_in[2];
	assign \mchip.top.frontend.rst  = io_in[2];
	assign \mchip.top.frontend.wclk  = io_in[0];
	assign \mchip.top.frontend.we  = io_in[3];
	assign \mchip.top.frontend.wptr  = \mchip.top.frontend.wptr_reg.q ;
	assign \mchip.top.frontend.wptr_b2g.binary  = \mchip.top.frontend.wptr_reg.q ;
	assign \mchip.top.frontend.wptr_b2g.gray  = {\mchip.top.frontend.wptr_reg.q [3], \mchip.top.frontend.wptr_gray [2:0]};
	assign \mchip.top.frontend.wptr_gray [3] = \mchip.top.frontend.wptr_reg.q [3];
	assign \mchip.top.frontend.wptr_reg.clk  = io_in[0];
	assign \mchip.top.frontend.wptr_reg.d [1] = \mchip.top.frontend.wptr_gray [0];
	assign \mchip.top.frontend.wptr_reg.rst  = io_in[2];
	assign \mchip.top.full  = \mchip.top.frontend.full ;
	assign \mchip.top.rclk  = io_in[1];
	assign \mchip.top.rdata  = io_out[7:5];
	assign \mchip.top.re  = io_in[4];
	assign \mchip.top.rptr  = \mchip.top.backend.rptr_reg.q ;
	assign \mchip.top.rptr_gray  = {\mchip.top.backend.rptr_reg.q [3], \mchip.top.backend.rptr_gray [2:0]};
	assign \mchip.top.rst  = io_in[2];
	assign \mchip.top.wclk  = io_in[0];
	assign \mchip.top.wdata  = io_in[7:5];
	assign \mchip.top.we  = io_in[3];
	assign \mchip.top.wptr  = \mchip.top.frontend.wptr_reg.q ;
	assign \mchip.top.wptr_gray  = {\mchip.top.frontend.wptr_reg.q [3], \mchip.top.frontend.wptr_gray [2:0]};
endmodule
module d41_stroucki_corralgame (
	io_in,
	io_out
);
	wire _000_;
	wire _001_;
	wire _002_;
	wire _003_;
	wire _004_;
	wire _005_;
	wire _006_;
	wire _007_;
	wire _008_;
	wire _009_;
	wire _010_;
	wire _011_;
	wire _012_;
	wire _013_;
	wire _014_;
	wire _015_;
	wire _016_;
	wire _017_;
	wire _018_;
	wire _019_;
	wire _020_;
	wire _021_;
	wire _022_;
	wire _023_;
	wire _024_;
	wire _025_;
	wire _026_;
	wire _027_;
	wire _028_;
	wire _029_;
	wire _030_;
	wire _031_;
	wire _032_;
	wire _033_;
	wire _034_;
	wire _035_;
	wire _036_;
	wire _037_;
	wire _038_;
	wire _039_;
	wire _040_;
	wire _041_;
	wire _042_;
	wire _043_;
	wire _044_;
	wire _045_;
	wire _046_;
	wire _047_;
	wire _048_;
	wire _049_;
	wire _050_;
	wire _051_;
	wire _052_;
	wire _053_;
	wire _054_;
	wire _055_;
	wire _056_;
	wire _057_;
	wire _058_;
	wire _059_;
	wire _060_;
	wire _061_;
	wire _062_;
	wire _063_;
	wire _064_;
	wire _065_;
	wire _066_;
	wire _067_;
	wire _068_;
	wire _069_;
	wire _070_;
	wire _071_;
	wire _072_;
	wire _073_;
	wire _074_;
	wire _075_;
	wire _076_;
	wire _077_;
	wire _078_;
	wire _079_;
	wire _080_;
	wire _081_;
	wire _082_;
	wire _083_;
	wire _084_;
	wire _085_;
	wire _086_;
	wire _087_;
	wire _088_;
	wire _089_;
	wire _090_;
	wire _091_;
	wire _092_;
	wire _093_;
	wire _094_;
	wire _095_;
	wire _096_;
	wire _097_;
	wire [31:0] _098_;
	wire [2:0] _099_;
	wire [2:0] _100_;
	input wire [13:0] io_in;
	output wire [13:0] io_out;
	wire \mchip.clock ;
	wire [3:0] \mchip.cowboypos ;
	wire [3:0] \mchip.data ;
	wire \mchip.enter ;
	wire \mchip.gameenter ;
	wire \mchip.gamegameover ;
	wire [31:0] \mchip.gameinstance.boltDest$func$d41_stroucki_corralgame/src/game.sv:154$21.boltStrength ;
	wire \mchip.gameinstance.boltDest$func$d41_stroucki_corralgame/src/game.sv:154$21.cowboyLeftOfHorse ;
	wire [3:0] \mchip.gameinstance.boltDest$func$d41_stroucki_corralgame/src/game.sv:154$21.horsePos ;
	wire [31:0] \mchip.gameinstance.boundHorse$func$d41_stroucki_corralgame/src/game.sv:144$17.horsePos ;
	wire [31:0] \mchip.gameinstance.boundHorse$func$d41_stroucki_corralgame/src/game.sv:144$17.targetHorsePos ;
	wire [31:0] \mchip.gameinstance.boundHorse$func$d41_stroucki_corralgame/src/game.sv:146$18.horsePos ;
	wire [31:0] \mchip.gameinstance.boundHorse$func$d41_stroucki_corralgame/src/game.sv:146$18.targetHorsePos ;
	wire [31:0] \mchip.gameinstance.boundHorse$func$d41_stroucki_corralgame/src/game.sv:151$20.horsePos ;
	wire [31:0] \mchip.gameinstance.boundHorse$func$d41_stroucki_corralgame/src/game.sv:151$20.targetHorsePos ;
	wire [31:0] \mchip.gameinstance.boundHorse$func$d41_stroucki_corralgame/src/game.sv:154$22.horsePos ;
	wire [31:0] \mchip.gameinstance.boundHorse$func$d41_stroucki_corralgame/src/game.sv:154$22.targetHorsePos ;
	wire [31:0] \mchip.gameinstance.boundHorse$func$d41_stroucki_corralgame/src/game.sv:156$23.horsePos ;
	wire [31:0] \mchip.gameinstance.boundHorse$func$d41_stroucki_corralgame/src/game.sv:156$23.targetHorsePos ;
	wire [31:0] \mchip.gameinstance.boundHorse$func$d41_stroucki_corralgame/src/game.sv:175$24.horsePos ;
	wire [31:0] \mchip.gameinstance.boundHorse$func$d41_stroucki_corralgame/src/game.sv:175$24.targetHorsePos ;
	wire \mchip.gameinstance.clock ;
	wire \mchip.gameinstance.cowboyDest$func$d41_stroucki_corralgame/src/game.sv:150$19.cowboyLeftOfHorse ;
	wire [3:0] \mchip.gameinstance.cowboyDest$func$d41_stroucki_corralgame/src/game.sv:150$19.cowboyPos ;
	wire [3:0] \mchip.gameinstance.cowboyDest$func$d41_stroucki_corralgame/src/game.sv:150$19.move ;
	wire [2:0] \mchip.gameinstance.cowboyHitpoints ;
	wire \mchip.gameinstance.cowboyInBound$func$d41_stroucki_corralgame/src/game.sv:122$16.cowboyLeftOfHorse ;
	wire [3:0] \mchip.gameinstance.cowboyInBound$func$d41_stroucki_corralgame/src/game.sv:122$16.cowboyPos ;
	wire [31:0] \mchip.gameinstance.cowboyInBound$func$d41_stroucki_corralgame/src/game.sv:122$16.dest ;
	wire [3:0] \mchip.gameinstance.cowboyInBound$func$d41_stroucki_corralgame/src/game.sv:122$16.move ;
	wire [3:0] \mchip.gameinstance.cowboyPos ;
	reg [3:0] \mchip.gameinstance.cowboypos ;
	wire [3:0] \mchip.gameinstance.distance ;
	wire \mchip.gameinstance.enter ;
	wire \mchip.gameinstance.gameover ;
	wire [3:0] \mchip.gameinstance.horsepos ;
	reg [2:0] \mchip.gameinstance.kickcount ;
	reg [2:0] \mchip.gameinstance.kickflight ;
	wire \mchip.gameinstance.lfsrinstance.i_Clk ;
	wire \mchip.gameinstance.lfsrinstance.i_Enable ;
	wire [4:0] \mchip.gameinstance.lfsrinstance.o_LFSR_Data ;
	wire [5:1] \mchip.gameinstance.lfsrinstance.r_LFSR ;
	wire [4:0] \mchip.gameinstance.lfsrout ;
	reg \mchip.gameinstance.lostwon ;
	wire [2:0] \mchip.gameinstance.move ;
	wire [2:0] \mchip.gameinstance.nextState ;
	wire [30:0] \mchip.gameinstance.p ;
	wire [3:0] \mchip.gameinstance.pVal ;
	wire [30:0] \mchip.gameinstance.q ;
	wire [3:0] \mchip.gameinstance.qVal ;
	wire [4:0] \mchip.gameinstance.randomVal ;
	wire \mchip.gameinstance.ready ;
	reg [2:0] \mchip.gameinstance.state  = 3'h1;
	wire \mchip.gameinstance.targetGameover ;
	wire [3:0] \mchip.gameinstance.targetHorsepos ;
	wire [2:0] \mchip.gameinstance.targetKickflight ;
	wire \mchip.gameinstance.targetLostwon ;
	wire [2:0] \mchip.gameinstance.targetMove ;
	wire \mchip.gamelostwon ;
	wire [2:0] \mchip.gamemove ;
	wire \mchip.gameover ;
	wire \mchip.gameready ;
	wire [7:0] \mchip.io_in ;
	wire [7:0] \mchip.io_out ;
	reg \mchip.lostwon ;
	wire [2:0] \mchip.move ;
	wire \mchip.ready ;
	wire \mchip.reset ;
	wire [2:0] \mchip.state ;
	assign _099_[0] = ~\mchip.gameinstance.kickcount [0];
	assign _042_ = ~(\mchip.gameinstance.state [1] | \mchip.gameinstance.state [0]);
	assign _043_ = _042_ & ~\mchip.gameinstance.state [2];
	assign _044_ = ~\mchip.gameinstance.state [2];
	assign _045_ = ~(\mchip.gameinstance.state [1] & \mchip.gameinstance.state [0]);
	assign _046_ = _044_ & ~_045_;
	assign _047_ = \mchip.gameinstance.state [0] | ~\mchip.gameinstance.state [1];
	assign _048_ = _044_ & ~_047_;
	assign _049_ = ~(_048_ | _046_);
	assign _050_ = _049_ & ~_043_;
	assign _002_ = _050_ & ~io_in[1];
	assign \mchip.gameinstance.move [0] = io_in[2] & io_in[5];
	assign _051_ = _042_ & ~_044_;
	assign _052_ = ~\mchip.gameinstance.cowboypos [2];
	assign _053_ = \mchip.gameinstance.cowboypos [1] | ~\mchip.gameinstance.horsepos [1];
	assign _054_ = ~\mchip.gameinstance.cowboypos [0];
	assign _055_ = \mchip.gameinstance.cowboypos [1] ^ \mchip.gameinstance.horsepos [1];
	assign _056_ = _054_ & ~_055_;
	assign _057_ = _056_ | ~_053_;
	assign _058_ = ~(_057_ & _052_);
	assign _059_ = \mchip.gameinstance.horsepos [1] ^ \mchip.gameinstance.cowboypos [3];
	assign _060_ = _059_ ^ _058_;
	assign _061_ = \mchip.gameinstance.cowboypos [3] | ~\mchip.gameinstance.horsepos [1];
	assign _062_ = _059_ | \mchip.gameinstance.cowboypos [2];
	assign _063_ = _057_ & ~_062_;
	assign _064_ = _061_ & ~_063_;
	assign _065_ = _052_ & ~_053_;
	assign _066_ = _065_ ^ _059_;
	assign _067_ = (_064_ ? _066_ : _060_);
	assign _068_ = _055_ ^ \mchip.gameinstance.cowboypos [0];
	assign _069_ = (_064_ ? _055_ : _068_);
	assign _070_ = (_064_ ? _053_ : _057_);
	assign _071_ = _070_ ^ \mchip.gameinstance.cowboypos [2];
	assign _072_ = _069_ | ~_071_;
	assign _073_ = ~(_072_ | _067_);
	assign _074_ = io_in[5] & io_in[4];
	assign _075_ = ~_074_;
	assign _076_ = _075_ ^ _067_;
	assign _077_ = io_in[3] & io_in[5];
	assign _078_ = _077_ | _071_;
	assign _079_ = _077_ ^ _071_;
	assign _080_ = \mchip.gameinstance.move [0] & ~_069_;
	assign _081_ = _079_ & ~_080_;
	assign _082_ = _078_ & ~_081_;
	assign _083_ = _076_ & ~_082_;
	assign _084_ = _067_ & ~_074_;
	assign _085_ = _084_ | _083_;
	assign _086_ = _085_ | _073_;
	assign _087_ = _051_ & ~_086_;
	assign _088_ = _069_ & ~_054_;
	assign _089_ = _067_ | ~_071_;
	assign _090_ = _089_ | _088_;
	assign _091_ = ~(_090_ & _086_);
	assign _092_ = _051_ & ~_091_;
	assign _093_ = _092_ | _087_;
	assign _000_ = _002_ & ~_093_;
	assign _094_ = (\mchip.gameinstance.state [0] ? \mchip.gameinstance.state [2] : \mchip.gameinstance.state [1]);
	assign _095_ = ~(\mchip.gameinstance.kickcount [2] | \mchip.gameinstance.kickcount [1]);
	assign _096_ = ~_095_;
	assign _097_ = _048_ & ~_096_;
	assign _004_ = _094_ & ~_097_;
	assign _005_ = ~(_046_ | _043_);
	assign _006_ = _048_ & ~_095_;
	assign _007_ = _006_ | io_in[1];
	assign _003_ = _005_ & ~_007_;
	assign _008_ = _007_ | _093_;
	assign _001_ = _005_ & ~_008_;
	assign _009_ = \mchip.gameinstance.state [0] & ~\mchip.gameinstance.state [1];
	assign \mchip.gameinstance.targetHorsepos [3] = _009_ & ~\mchip.gameinstance.state [2];
	assign _010_ = _077_ ^ \mchip.gameinstance.move [0];
	assign _098_[1] = (_064_ ? _010_ : _077_);
	assign _011_ = ~(_077_ | \mchip.gameinstance.move [0]);
	assign _012_ = _011_ ^ _075_;
	assign _098_[2] = (_064_ ? _012_ : _074_);
	assign _013_ = _011_ & ~_074_;
	assign _098_[31] = _064_ & ~_013_;
	assign _014_ = ~\mchip.gameinstance.kickflight [0];
	assign _015_ = (\mchip.gameinstance.state [2] ? _042_ : _009_);
	assign \mchip.gameinstance.targetKickflight [0] = (_015_ ? _051_ : _014_);
	assign _016_ = ~(\mchip.gameinstance.kickflight [1] ^ \mchip.gameinstance.kickflight [0]);
	assign \mchip.gameinstance.targetKickflight [1] = _016_ & ~_015_;
	assign _017_ = ~(\mchip.gameinstance.kickflight [1] | \mchip.gameinstance.kickflight [0]);
	assign _018_ = _017_ ^ \mchip.gameinstance.kickflight [2];
	assign \mchip.gameinstance.targetKickflight [2] = _018_ & ~_015_;
	assign _019_ = ~io_in[5];
	assign _020_ = _046_ & ~_019_;
	assign _021_ = _020_ | _006_;
	assign _022_ = _086_ & ~_090_;
	assign _023_ = _051_ & ~_022_;
	assign _024_ = _023_ | \mchip.gameinstance.targetHorsepos [3];
	assign _025_ = _024_ | _021_;
	assign _026_ = _049_ & ~_015_;
	assign \mchip.gameinstance.nextState [0] = _025_ & ~_026_;
	assign _027_ = \mchip.gameinstance.kickflight [0] & ~\mchip.gameinstance.kickflight [1];
	assign _028_ = _027_ & ~_018_;
	assign _029_ = _028_ | _096_;
	assign _030_ = _048_ & ~_029_;
	assign _031_ = ~(_030_ | _020_);
	assign _032_ = _031_ & ~_015_;
	assign \mchip.gameinstance.nextState [1] = ~(_032_ | _026_);
	assign _033_ = ~(_098_[31] | _098_[2]);
	assign _034_ = _098_[1] | \mchip.gameinstance.move [0];
	assign _035_ = _033_ & ~_034_;
	assign _036_ = _035_ | _098_[31];
	assign _037_ = _077_ & _074_;
	assign _038_ = _013_ | _019_;
	assign _039_ = _038_ | _037_;
	assign _040_ = _039_ | _036_;
	assign \mchip.gameinstance.nextState [2] = _026_ & ~_040_;
	assign _100_[1] = \mchip.gameinstance.kickcount [1] ^ \mchip.gameinstance.kickcount [0];
	assign _041_ = \mchip.gameinstance.kickcount [1] & \mchip.gameinstance.kickcount [0];
	assign _100_[2] = _041_ ^ \mchip.gameinstance.kickcount [2];
	always @(posedge io_in[0])
		if (_002_)
			if (\mchip.gameinstance.targetHorsepos [3])
				\mchip.gameinstance.cowboypos [0] <= 1'h0;
			else
				\mchip.gameinstance.cowboypos [0] <= \mchip.gameinstance.move [0];
	always @(posedge io_in[0])
		if (_002_)
			if (\mchip.gameinstance.targetHorsepos [3])
				\mchip.gameinstance.cowboypos [1] <= 1'h0;
			else
				\mchip.gameinstance.cowboypos [1] <= _098_[1];
	always @(posedge io_in[0])
		if (_002_)
			if (\mchip.gameinstance.targetHorsepos [3])
				\mchip.gameinstance.cowboypos [2] <= 1'h0;
			else
				\mchip.gameinstance.cowboypos [2] <= _098_[2];
	always @(posedge io_in[0])
		if (_002_)
			if (\mchip.gameinstance.targetHorsepos [3])
				\mchip.gameinstance.cowboypos [3] <= 1'h0;
			else
				\mchip.gameinstance.cowboypos [3] <= _098_[31];
	always @(posedge io_in[0])
		if (_001_)
			\mchip.gameinstance.kickflight [0] <= \mchip.gameinstance.targetKickflight [0];
	always @(posedge io_in[0])
		if (_001_)
			\mchip.gameinstance.kickflight [1] <= \mchip.gameinstance.targetKickflight [1];
	always @(posedge io_in[0])
		if (_001_)
			\mchip.gameinstance.kickflight [2] <= \mchip.gameinstance.targetKickflight [2];
	always @(posedge io_in[0])
		if (_000_)
			if (\mchip.gameinstance.targetHorsepos [3])
				\mchip.gameinstance.kickcount [0] <= 1'h0;
			else
				\mchip.gameinstance.kickcount [0] <= _099_[0];
	always @(posedge io_in[0])
		if (_000_)
			if (\mchip.gameinstance.targetHorsepos [3])
				\mchip.gameinstance.kickcount [1] <= 1'h0;
			else
				\mchip.gameinstance.kickcount [1] <= _100_[1];
	always @(posedge io_in[0])
		if (_000_)
			if (\mchip.gameinstance.targetHorsepos [3])
				\mchip.gameinstance.kickcount [2] <= 1'h0;
			else
				\mchip.gameinstance.kickcount [2] <= _100_[2];
	reg \mchip.gameinstance.horsepos_reg[1] ;
	always @(posedge io_in[0])
		if (_003_)
			\mchip.gameinstance.horsepos_reg[1]  <= \mchip.gameinstance.targetHorsepos [3];
	assign \mchip.gameinstance.horsepos [1] = \mchip.gameinstance.horsepos_reg[1] ;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.gameinstance.lostwon  <= 1'h1;
		else if (_004_)
			\mchip.gameinstance.lostwon  <= 1'h0;
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.gameinstance.state [0] <= 1'h1;
		else
			\mchip.gameinstance.state [0] <= \mchip.gameinstance.nextState [0];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.gameinstance.state [1] <= 1'h0;
		else
			\mchip.gameinstance.state [1] <= \mchip.gameinstance.nextState [1];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.gameinstance.state [2] <= 1'h0;
		else
			\mchip.gameinstance.state [2] <= \mchip.gameinstance.nextState [2];
	always @(posedge io_in[0])
		if (!io_in[1])
			\mchip.lostwon  <= \mchip.gameinstance.lostwon ;
	assign {_098_[30:3], _098_[0]} = {_098_[31], _098_[31], _098_[31], _098_[31], _098_[31], _098_[31], _098_[31], _098_[31], _098_[31], _098_[31], _098_[31], _098_[31], _098_[31], _098_[31], _098_[31], _098_[31], _098_[31], _098_[31], _098_[31], _098_[31], _098_[31], _098_[31], _098_[31], _098_[31], _098_[31], _098_[31], _098_[31], _098_[31], \mchip.gameinstance.move [0]};
	assign _099_[2:1] = \mchip.gameinstance.kickcount [2:1];
	assign _100_[0] = _099_[0];
	assign io_out = {8'h00, \mchip.lostwon , 5'h10};
	assign \mchip.clock  = io_in[0];
	assign \mchip.cowboypos  = 4'h0;
	assign \mchip.data  = 4'h0;
	assign \mchip.enter  = io_in[5];
	assign \mchip.gameenter  = io_in[5];
	assign \mchip.gamegameover  = 1'h1;
	assign \mchip.gameinstance.boltDest$func$d41_stroucki_corralgame/src/game.sv:154$21.boltStrength  = 32'd0;
	assign \mchip.gameinstance.boltDest$func$d41_stroucki_corralgame/src/game.sv:154$21.cowboyLeftOfHorse  = 1'h0;
	assign \mchip.gameinstance.boltDest$func$d41_stroucki_corralgame/src/game.sv:154$21.horsePos  = 4'h0;
	assign \mchip.gameinstance.boundHorse$func$d41_stroucki_corralgame/src/game.sv:144$17.horsePos  = 32'd0;
	assign \mchip.gameinstance.boundHorse$func$d41_stroucki_corralgame/src/game.sv:144$17.targetHorsePos  = 32'd0;
	assign \mchip.gameinstance.boundHorse$func$d41_stroucki_corralgame/src/game.sv:146$18.horsePos  = 32'd0;
	assign \mchip.gameinstance.boundHorse$func$d41_stroucki_corralgame/src/game.sv:146$18.targetHorsePos  = 32'd0;
	assign \mchip.gameinstance.boundHorse$func$d41_stroucki_corralgame/src/game.sv:151$20.horsePos  = 32'd0;
	assign \mchip.gameinstance.boundHorse$func$d41_stroucki_corralgame/src/game.sv:151$20.targetHorsePos  = 32'd0;
	assign \mchip.gameinstance.boundHorse$func$d41_stroucki_corralgame/src/game.sv:154$22.horsePos  = 32'd0;
	assign \mchip.gameinstance.boundHorse$func$d41_stroucki_corralgame/src/game.sv:154$22.targetHorsePos  = 32'd0;
	assign \mchip.gameinstance.boundHorse$func$d41_stroucki_corralgame/src/game.sv:156$23.horsePos  = 32'd0;
	assign \mchip.gameinstance.boundHorse$func$d41_stroucki_corralgame/src/game.sv:156$23.targetHorsePos  = 32'd0;
	assign \mchip.gameinstance.boundHorse$func$d41_stroucki_corralgame/src/game.sv:175$24.horsePos  = 32'd0;
	assign \mchip.gameinstance.boundHorse$func$d41_stroucki_corralgame/src/game.sv:175$24.targetHorsePos  = 32'd0;
	assign \mchip.gameinstance.clock  = io_in[0];
	assign \mchip.gameinstance.cowboyDest$func$d41_stroucki_corralgame/src/game.sv:150$19.cowboyLeftOfHorse  = 1'h0;
	assign \mchip.gameinstance.cowboyDest$func$d41_stroucki_corralgame/src/game.sv:150$19.cowboyPos  = 4'h0;
	assign \mchip.gameinstance.cowboyDest$func$d41_stroucki_corralgame/src/game.sv:150$19.move  = 4'h0;
	assign \mchip.gameinstance.cowboyHitpoints  = 3'h1;
	assign \mchip.gameinstance.cowboyInBound$func$d41_stroucki_corralgame/src/game.sv:122$16.cowboyLeftOfHorse  = 1'h0;
	assign \mchip.gameinstance.cowboyInBound$func$d41_stroucki_corralgame/src/game.sv:122$16.cowboyPos  = 4'h0;
	assign \mchip.gameinstance.cowboyInBound$func$d41_stroucki_corralgame/src/game.sv:122$16.dest  = 32'd0;
	assign \mchip.gameinstance.cowboyInBound$func$d41_stroucki_corralgame/src/game.sv:122$16.move  = 4'h0;
	assign \mchip.gameinstance.cowboyPos  = 4'h0;
	assign \mchip.gameinstance.distance  = {3'h0, \mchip.gameinstance.cowboypos [0]};
	assign \mchip.gameinstance.enter  = io_in[5];
	assign \mchip.gameinstance.gameover  = 1'h1;
	assign {\mchip.gameinstance.horsepos [3:2], \mchip.gameinstance.horsepos [0]} = {\mchip.gameinstance.horsepos [1], 2'h0};
	assign \mchip.gameinstance.lfsrinstance.i_Clk  = io_in[0];
	assign \mchip.gameinstance.lfsrinstance.i_Enable  = 1'h0;
	assign \mchip.gameinstance.lfsrinstance.o_LFSR_Data  = 5'h00;
	assign \mchip.gameinstance.lfsrinstance.r_LFSR  = 5'h00;
	assign \mchip.gameinstance.lfsrout  = 5'h00;
	assign \mchip.gameinstance.move [2:1] = 2'h0;
	assign \mchip.gameinstance.p  = 31'h2332210f;
	assign \mchip.gameinstance.pVal  = 4'hf;
	assign \mchip.gameinstance.q  = 31'h34543210;
	assign \mchip.gameinstance.qVal  = 4'h0;
	assign \mchip.gameinstance.randomVal  = 5'h00;
	assign \mchip.gameinstance.ready  = 1'h0;
	assign \mchip.gameinstance.targetGameover  = 1'h1;
	assign \mchip.gameinstance.targetHorsepos [2:0] = {1'h0, \mchip.gameinstance.targetHorsepos [3], 1'h0};
	assign \mchip.gameinstance.targetLostwon  = 1'h0;
	assign \mchip.gameinstance.targetMove  = {2'h0, \mchip.gameinstance.move [0]};
	assign \mchip.gamelostwon  = \mchip.gameinstance.lostwon ;
	assign \mchip.gamemove  = {2'h0, \mchip.gameinstance.move [0]};
	assign \mchip.gameover  = 1'h1;
	assign \mchip.gameready  = 1'h0;
	assign \mchip.io_in  = io_in[7:0];
	assign \mchip.io_out  = {2'h0, \mchip.lostwon , 5'h10};
	assign \mchip.move  = io_in[4:2];
	assign \mchip.ready  = 1'h0;
	assign \mchip.reset  = io_in[1];
	assign \mchip.state  = 3'h3;
endmodule
module d42_qilins_sevenseg (
	io_in,
	io_out
);
	wire _00_;
	wire _01_;
	wire _02_;
	wire _03_;
	wire _04_;
	wire _05_;
	wire _06_;
	wire _07_;
	wire _08_;
	wire _09_;
	wire _10_;
	wire _11_;
	wire _12_;
	wire _13_;
	wire _14_;
	wire _15_;
	wire _16_;
	wire _17_;
	wire _18_;
	wire _19_;
	wire _20_;
	wire _21_;
	wire _22_;
	wire _23_;
	wire _24_;
	wire _25_;
	wire _26_;
	wire _27_;
	wire _28_;
	wire _29_;
	wire _30_;
	wire _31_;
	wire _32_;
	wire _33_;
	wire _34_;
	wire _35_;
	wire _36_;
	wire _37_;
	wire _38_;
	wire _39_;
	wire _40_;
	wire _41_;
	wire _42_;
	wire _43_;
	wire _44_;
	input wire [13:0] io_in;
	output wire [13:0] io_out;
	wire \mchip.gate10.in ;
	wire \mchip.gate11.b ;
	wire \mchip.gate15.a ;
	wire \mchip.gate16.a ;
	wire \mchip.gate17.a ;
	wire \mchip.gate17.b ;
	wire \mchip.gate20.out ;
	wire \mchip.gate22.a ;
	wire \mchip.gate24.b ;
	wire \mchip.gate25.b ;
	wire \mchip.gate26.a ;
	wire \mchip.gate27.b ;
	wire \mchip.gate28.a ;
	wire \mchip.gate28.b ;
	wire \mchip.gate34.out ;
	wire \mchip.gate36.b ;
	wire \mchip.gate37.a ;
	wire \mchip.gate38.a ;
	wire \mchip.gate39.a ;
	wire \mchip.gate45.out ;
	wire \mchip.gate47.b ;
	wire \mchip.gate48.b ;
	wire \mchip.gate49.b ;
	wire \mchip.gate50.a ;
	wire \mchip.gate53.out ;
	wire \mchip.gate57.b ;
	wire \mchip.gate58.b ;
	wire \mchip.gate59.a ;
	wire \mchip.gate60.b ;
	wire \mchip.gate61.a ;
	wire \mchip.gate61.b ;
	wire \mchip.gate63.a ;
	wire \mchip.gate68.out ;
	wire \mchip.gate69.a ;
	wire \mchip.gate7.in ;
	wire \mchip.gate70.a ;
	wire \mchip.gate70.b ;
	wire \mchip.gate71.a ;
	wire \mchip.gate71.b ;
	wire \mchip.gate74.out ;
	wire \mchip.gate75.b ;
	wire \mchip.gate77.b ;
	wire \mchip.gate78.a ;
	wire \mchip.gate79.a ;
	wire \mchip.gate8.in ;
	wire \mchip.gate80.a ;
	wire \mchip.gate80.b ;
	wire \mchip.gate83.out ;
	wire \mchip.gate85.a ;
	wire \mchip.gate85.out ;
	wire \mchip.gate9.in ;
	wire [7:0] \mchip.io_in ;
	wire [7:0] \mchip.io_out ;
	wire \mchip.net1 ;
	wire \mchip.net10 ;
	wire \mchip.net11 ;
	wire \mchip.net12 ;
	wire \mchip.net13 ;
	wire \mchip.net14 ;
	wire \mchip.net2 ;
	wire \mchip.net3 ;
	wire \mchip.net4 ;
	wire \mchip.net5 ;
	wire \mchip.net6 ;
	wire \mchip.net7 ;
	wire \mchip.net8 ;
	wire \mchip.net9 ;
	assign _00_ = io_in[2] | ~io_in[0];
	assign _01_ = ~io_in[3];
	assign _02_ = io_in[2] & io_in[1];
	assign _03_ = io_in[1] & ~io_in[2];
	assign _04_ = (io_in[3] ? _03_ : _02_);
	assign _05_ = ~(io_in[1] | io_in[0]);
	assign _06_ = io_in[2] & ~io_in[1];
	assign _07_ = (io_in[3] ? _06_ : _05_);
	assign _08_ = ~(_07_ | _04_);
	assign \mchip.gate68.out  = ~(_08_ & _00_);
	assign _09_ = io_in[0] & ~io_in[1];
	assign _10_ = io_in[1] & ~io_in[0];
	assign _11_ = io_in[3] & ~io_in[2];
	assign _12_ = _11_ | _10_;
	assign _13_ = io_in[3] & ~io_in[0];
	assign _14_ = ~(io_in[2] | io_in[0]);
	assign _15_ = _14_ | _13_;
	assign _16_ = _15_ | _12_;
	assign \mchip.gate53.out  = _16_ | _09_;
	assign _17_ = ~(io_in[1] | io_in[3]);
	assign _18_ = ~(io_in[2] | io_in[1]);
	assign _19_ = io_in[3] & ~_00_;
	assign _20_ = _19_ | _18_;
	assign _21_ = io_in[2] & ~io_in[0];
	assign _22_ = (io_in[3] ? _21_ : _14_);
	assign _23_ = _22_ | _20_;
	assign \mchip.gate45.out  = _23_ | _17_;
	assign _24_ = _17_ | _02_;
	assign _25_ = (io_in[0] ? _01_ : io_in[2]);
	assign _26_ = io_in[0] | ~io_in[1];
	assign _27_ = io_in[3] & ~_26_;
	assign _28_ = _09_ & ~io_in[2];
	assign _29_ = _28_ | _27_;
	assign _30_ = _29_ | _25_;
	assign \mchip.gate34.out  = _30_ | _24_;
	assign _31_ = io_in[2] & io_in[0];
	assign _32_ = (io_in[1] ? _01_ : io_in[0]);
	assign _33_ = _32_ | _31_;
	assign _34_ = ~(io_in[2] | io_in[3]);
	assign _35_ = _10_ & ~io_in[2];
	assign _36_ = _35_ | _34_;
	assign \mchip.gate20.out  = _36_ | _33_;
	assign \mchip.gate85.out  = io_in[0] & ~_18_;
	assign _37_ = io_in[0] & io_in[3];
	assign _38_ = io_in[2] & ~io_in[3];
	assign _39_ = ~(_38_ | _09_);
	assign _40_ = (io_in[2] ? io_in[1] : _26_);
	assign _41_ = ~(_40_ & _39_);
	assign \mchip.gate83.out  = _41_ | _37_;
	assign _42_ = io_in[1] & io_in[0];
	assign _43_ = _42_ | _31_;
	assign _44_ = _38_ | _17_;
	assign \mchip.gate74.out  = _44_ | _43_;
	assign io_out = {6'h00, \mchip.gate85.out , \mchip.gate83.out , \mchip.gate20.out , \mchip.gate74.out , \mchip.gate68.out , \mchip.gate53.out , \mchip.gate45.out , \mchip.gate34.out };
	assign \mchip.gate10.in  = io_in[3];
	assign \mchip.gate11.b  = io_in[1];
	assign \mchip.gate15.a  = io_in[1];
	assign \mchip.gate16.a  = io_in[0];
	assign \mchip.gate17.a  = io_in[0];
	assign \mchip.gate17.b  = io_in[2];
	assign \mchip.gate22.a  = io_in[0];
	assign \mchip.gate24.b  = io_in[1];
	assign \mchip.gate25.b  = io_in[3];
	assign \mchip.gate26.a  = io_in[0];
	assign \mchip.gate27.b  = io_in[2];
	assign \mchip.gate28.a  = io_in[1];
	assign \mchip.gate28.b  = io_in[2];
	assign \mchip.gate36.b  = io_in[2];
	assign \mchip.gate37.a  = io_in[3];
	assign \mchip.gate38.a  = io_in[0];
	assign \mchip.gate39.a  = io_in[3];
	assign \mchip.gate47.b  = io_in[3];
	assign \mchip.gate48.b  = io_in[3];
	assign \mchip.gate49.b  = io_in[1];
	assign \mchip.gate50.a  = io_in[0];
	assign \mchip.gate57.b  = io_in[2];
	assign \mchip.gate58.b  = io_in[3];
	assign \mchip.gate59.a  = io_in[1];
	assign \mchip.gate60.b  = io_in[3];
	assign \mchip.gate61.a  = io_in[1];
	assign \mchip.gate61.b  = io_in[2];
	assign \mchip.gate63.a  = io_in[0];
	assign \mchip.gate69.a  = io_in[2];
	assign \mchip.gate7.in  = io_in[0];
	assign \mchip.gate70.a  = io_in[0];
	assign \mchip.gate70.b  = io_in[2];
	assign \mchip.gate71.a  = io_in[0];
	assign \mchip.gate71.b  = io_in[1];
	assign \mchip.gate75.b  = io_in[1];
	assign \mchip.gate77.b  = io_in[2];
	assign \mchip.gate78.a  = io_in[2];
	assign \mchip.gate79.a  = io_in[0];
	assign \mchip.gate8.in  = io_in[1];
	assign \mchip.gate80.a  = io_in[0];
	assign \mchip.gate80.b  = io_in[3];
	assign \mchip.gate85.a  = io_in[0];
	assign \mchip.gate9.in  = io_in[2];
	assign \mchip.io_in  = io_in[7:0];
	assign \mchip.io_out  = {\mchip.gate85.out , \mchip.gate83.out , \mchip.gate20.out , \mchip.gate74.out , \mchip.gate68.out , \mchip.gate53.out , \mchip.gate45.out , \mchip.gate34.out };
	assign \mchip.net1  = io_in[0];
	assign \mchip.net10  = \mchip.gate20.out ;
	assign \mchip.net11  = \mchip.gate83.out ;
	assign \mchip.net12  = \mchip.gate85.out ;
	assign \mchip.net13  = 1'h0;
	assign \mchip.net14  = 1'h1;
	assign \mchip.net2  = io_in[1];
	assign \mchip.net3  = io_in[2];
	assign \mchip.net4  = io_in[3];
	assign \mchip.net5  = \mchip.gate34.out ;
	assign \mchip.net6  = \mchip.gate45.out ;
	assign \mchip.net7  = \mchip.gate53.out ;
	assign \mchip.net8  = \mchip.gate68.out ;
	assign \mchip.net9  = \mchip.gate74.out ;
endmodule
module d43_mmx_counter (
	io_in,
	io_out
);
	wire _00_;
	wire _01_;
	wire _02_;
	wire _03_;
	wire _04_;
	wire _05_;
	wire _06_;
	wire [6:0] _07_;
	wire [6:0] _08_;
	input wire [13:0] io_in;
	output wire [13:0] io_out;
	wire \mchip.clk ;
	reg [6:0] \mchip.counter ;
	wire [7:0] \mchip.io_in ;
	wire [7:0] \mchip.io_out ;
	wire \mchip.reset ;
	assign _07_[0] = ~\mchip.counter [0];
	assign _08_[1] = \mchip.counter [1] ^ \mchip.counter [0];
	assign _00_ = \mchip.counter [1] & \mchip.counter [0];
	assign _08_[2] = _00_ ^ \mchip.counter [2];
	assign _01_ = _00_ & \mchip.counter [2];
	assign _08_[3] = _01_ ^ \mchip.counter [3];
	assign _02_ = ~(\mchip.counter [3] & \mchip.counter [2]);
	assign _03_ = _00_ & ~_02_;
	assign _08_[4] = _03_ ^ \mchip.counter [4];
	assign _04_ = _03_ & \mchip.counter [4];
	assign _08_[5] = _04_ ^ \mchip.counter [5];
	assign _05_ = ~(\mchip.counter [5] & \mchip.counter [4]);
	assign _06_ = _03_ & ~_05_;
	assign _08_[6] = _06_ ^ \mchip.counter [6];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.counter [0] <= 1'h0;
		else
			\mchip.counter [0] <= _07_[0];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.counter [1] <= 1'h0;
		else
			\mchip.counter [1] <= _08_[1];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.counter [2] <= 1'h0;
		else
			\mchip.counter [2] <= _08_[2];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.counter [3] <= 1'h0;
		else
			\mchip.counter [3] <= _08_[3];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.counter [4] <= 1'h0;
		else
			\mchip.counter [4] <= _08_[4];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.counter [5] <= 1'h0;
		else
			\mchip.counter [5] <= _08_[5];
	always @(posedge io_in[0])
		if (io_in[1])
			\mchip.counter [6] <= 1'h0;
		else
			\mchip.counter [6] <= _08_[6];
	assign _07_[6:1] = \mchip.counter [6:1];
	assign _08_[0] = _07_[0];
	assign io_out = {7'h00, \mchip.counter };
	assign \mchip.clk  = io_in[0];
	assign \mchip.io_in  = io_in[7:0];
	assign \mchip.io_out  = {1'h0, \mchip.counter };
	assign \mchip.reset  = io_in[1];
endmodule
`default_nettype none
module multiplexer (
	io_in,
	io_out,
	des_sel,
	hold_if_not_sel,
	des_io_in,
	des_reset,
	des_io_out,
	clock,
	reset
);
	input wire [11:0] io_in;
	output reg [11:0] io_out;
	input wire [5:0] des_sel;
	input wire hold_if_not_sel;
	output reg [767:0] des_io_in;
	output reg [0:63] des_reset;
	input wire [767:0] des_io_out;
	input wire clock;
	input wire reset;
	reg [63:0] des_sel_dec;
	always @(posedge clock) begin
		des_sel_dec <= 1'sb0;
		des_sel_dec[des_sel] <= 1;
	end
	integer i;
	always @(*) begin
		io_out = 1'sb0;
		for (i = 0; i < 64; i = i + 1)
			begin
				if (des_sel_dec[i])
					io_out = des_io_out[(63 - i) * 12+:12];
				if (hold_if_not_sel && !des_sel_dec[i]) begin
					des_io_in[(63 - i) * 12+:12] = 1'sb0;
					des_reset[i] = 1'sb1;
				end
				else begin
					des_io_in[(63 - i) * 12+:12] = io_in;
					des_reset[i] = reset;
				end
			end
	end
endmodule
`default_nettype none
module design_instantiations (
	io_in,
	io_out,
	des_sel,
	hold_if_not_sel,
	clock,
	reset
);
	input wire [11:0] io_in;
	output wire [11:0] io_out;
	input wire [5:0] des_sel;
	input wire hold_if_not_sel;
	input wire clock;
	input wire reset;
	wire [767:0] des_io_in;
	wire [767:0] des_io_out;
	wire [0:63] des_reset;
	multiplexer mux(
		.io_in(io_in),
		.io_out(io_out),
		.des_sel(des_sel),
		.hold_if_not_sel(hold_if_not_sel),
		.des_io_in(des_io_in),
		.des_reset(des_reset),
		.des_io_out(des_io_out),
		.clock(clock),
		.reset(reset)
	);
	assign des_io_out[756+:12] = 12'h000;
	d01_example_adder inst1(
		.io_in({des_reset[1], clock, des_io_in[744+:12]}),
		.io_out(des_io_out[744+:12])
	);
	d02_example_counter inst2(
		.io_in({des_reset[2], clock, des_io_in[732+:12]}),
		.io_out(des_io_out[732+:12])
	);
	d03_example_beepboop inst3(
		.io_in({des_reset[3], clock, des_io_in[720+:12]}),
		.io_out(des_io_out[720+:12])
	);
	d04_example_aes128sca inst4(
		.io_in({des_reset[4], clock, des_io_in[708+:12]}),
		.io_out(des_io_out[708+:12])
	);
	d05_meta_info inst5(
		.io_in({des_reset[5], clock, des_io_in[696+:12]}),
		.io_out(des_io_out[696+:12])
	);
	assign des_io_out[684+:12] = 12'h000;
	assign des_io_out[672+:12] = 12'h000;
	assign des_io_out[660+:12] = 12'h000;
	assign des_io_out[648+:12] = 12'h000;
	assign des_io_out[636+:12] = 12'h000;
	d11_gbailey_bfchip inst11(
		.io_in({des_reset[11], clock, des_io_in[624+:12]}),
		.io_out(des_io_out[624+:12])
	);
	d12_oball_i2c inst12(
		.io_in({des_reset[12], clock, des_io_in[612+:12]}),
		.io_out(des_io_out[612+:12])
	);
	d13_jrduvall_s444 inst13(
		.io_in({des_reset[13], clock, des_io_in[600+:12]}),
		.io_out(des_io_out[600+:12])
	);
	d14_jessief_trafficlight inst14(
		.io_in({des_reset[14], clock, des_io_in[588+:12]}),
		.io_out(des_io_out[588+:12])
	);
	d15_jerryfen_prng inst15(
		.io_in({des_reset[15], clock, des_io_in[576+:12]}),
		.io_out(des_io_out[576+:12])
	);
	d16_bgonzale_pll inst16(
		.io_in({des_reset[16], clock, des_io_in[564+:12]}),
		.io_out(des_io_out[564+:12])
	);
	d17_njayawar_tetris inst17(
		.io_in({des_reset[17], clock, des_io_in[552+:12]}),
		.io_out(des_io_out[552+:12])
	);
	d18_nikhildj_mac inst18(
		.io_in({des_reset[18], clock, des_io_in[540+:12]}),
		.io_out(des_io_out[540+:12])
	);
	d19_rdkapur_encryptor inst19(
		.io_in({des_reset[19], clock, des_io_in[528+:12]}),
		.io_out(des_io_out[528+:12])
	);
	d20_rashik_tetris inst20(
		.io_in({des_reset[20], clock, des_io_in[516+:12]}),
		.io_out(des_io_out[516+:12])
	);
	d21_varunk2_motorctrl inst21(
		.io_in({des_reset[21], clock, des_io_in[504+:12]}),
		.io_out(des_io_out[504+:12])
	);
	d22_yushuanl_convolution inst22(
		.io_in({des_reset[22], clock, des_io_in[492+:12]}),
		.io_out(des_io_out[492+:12])
	);
	d23_zhiyingm_turing inst23(
		.io_in({des_reset[23], clock, des_io_in[480+:12]}),
		.io_out(des_io_out[480+:12])
	);
	d24_mnguyen2_tpu inst24(
		.io_in({des_reset[24], clock, des_io_in[468+:12]}),
		.io_out(des_io_out[468+:12])
	);
	d25_araghave_huffman inst25(
		.io_in({des_reset[25], clock, des_io_in[456+:12]}),
		.io_out(des_io_out[456+:12])
	);
	d26_cjstange_perceptron inst26(
		.io_in({des_reset[26], clock, des_io_in[444+:12]}),
		.io_out(des_io_out[444+:12])
	);
	d27_svemulap_fpu inst27(
		.io_in({des_reset[27], clock, des_io_in[432+:12]}),
		.io_out(des_io_out[432+:12])
	);
	d28_gvenkata_ucpu inst28(
		.io_in({des_reset[28], clock, des_io_in[420+:12]}),
		.io_out(des_io_out[420+:12])
	);
	d29_bwilhelm_i8008 inst29(
		.io_in({des_reset[29], clock, des_io_in[408+:12]}),
		.io_out(des_io_out[408+:12])
	);
	d30_yuchingw_fpga inst30(
		.io_in({des_reset[30], clock, des_io_in[396+:12]}),
		.io_out(des_io_out[396+:12])
	);
	d31_mdhamank_lfsr inst31(
		.io_in({des_reset[31], clock, des_io_in[384+:12]}),
		.io_out(des_io_out[384+:12])
	);
	d32_ngaertne_cpu inst32(
		.io_in({des_reset[32], clock, des_io_in[372+:12]}),
		.io_out(des_io_out[372+:12])
	);
	d33_mgee3_adder inst33(
		.io_in({des_reset[33], clock, des_io_in[360+:12]}),
		.io_out(des_io_out[360+:12])
	);
	d34_hgrodin_collatz inst34(
		.io_in({des_reset[34], clock, des_io_in[348+:12]}),
		.io_out(des_io_out[348+:12])
	);
	d35_ckasuba_comparator inst35(
		.io_in({des_reset[35], clock, des_io_in[336+:12]}),
		.io_out(des_io_out[336+:12])
	);
	d36_jxli_fpmul inst36(
		.io_in({des_reset[36], clock, des_io_in[324+:12]}),
		.io_out(des_io_out[324+:12])
	);
	d37_sophiali_calculator inst37(
		.io_in({des_reset[37], clock, des_io_in[312+:12]}),
		.io_out(des_io_out[312+:12])
	);
	d38_jxlu_pwm inst38(
		.io_in({des_reset[38], clock, des_io_in[300+:12]}),
		.io_out(des_io_out[300+:12])
	);
	d39_oonyeado_sevenseg inst39(
		.io_in({des_reset[39], clock, des_io_in[288+:12]}),
		.io_out(des_io_out[288+:12])
	);
	d40_jrecta_asyncfifo inst40(
		.io_in({des_reset[40], clock, des_io_in[276+:12]}),
		.io_out(des_io_out[276+:12])
	);
	d41_stroucki_corralgame inst41(
		.io_in({des_reset[41], clock, des_io_in[264+:12]}),
		.io_out(des_io_out[264+:12])
	);
	d42_qilins_sevenseg inst42(
		.io_in({des_reset[42], clock, des_io_in[252+:12]}),
		.io_out(des_io_out[252+:12])
	);
	d43_mmx_counter inst43(
		.io_in({des_reset[43], clock, des_io_in[240+:12]}),
		.io_out(des_io_out[240+:12])
	);
	assign des_io_out[228+:12] = 12'h000;
	assign des_io_out[216+:12] = 12'h000;
	assign des_io_out[204+:12] = 12'h000;
	assign des_io_out[192+:12] = 12'h000;
	assign des_io_out[180+:12] = 12'h000;
	assign des_io_out[168+:12] = 12'h000;
	assign des_io_out[156+:12] = 12'h000;
	assign des_io_out[144+:12] = 12'h000;
	assign des_io_out[132+:12] = 12'h000;
	assign des_io_out[120+:12] = 12'h000;
	assign des_io_out[108+:12] = 12'h000;
	assign des_io_out[96+:12] = 12'h000;
	assign des_io_out[84+:12] = 12'h000;
	assign des_io_out[72+:12] = 12'h000;
	assign des_io_out[60+:12] = 12'h000;
	assign des_io_out[48+:12] = 12'h000;
	assign des_io_out[36+:12] = 12'h000;
	assign des_io_out[24+:12] = 12'h000;
	assign des_io_out[12+:12] = 12'h000;
	assign des_io_out[0+:12] = 12'h000;
endmodule
