`ifndef DEFINES_H
`define DEFINES_H

`define DATA_WIDTH 8

typedef logic [`DATA_WIDTH-1:0] data_t;

`endif
