
`default_nettype none

module my_chip (
    input logic [11:0] io_in,
    input logic clock, reset,
    output logic [11:0] io_out
);

wire [7:0] val;

always_ff @(posedge clock) io_out <= {4'b0000, val};

assign val[0] = (io_in[0] & ~io_in[1] & ~io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[6] & ~io_in[7] & io_in[8] & io_in[10] & ~io_in[11]) | (~io_in[1] & ~io_in[2] & io_in[4] & io_in[6] & io_in[7] & io_in[8] & ~io_in[9] & io_in[11]) | (io_in[0] & io_in[2] & io_in[3] & ~io_in[6] & io_in[7] & io_in[8] & io_in[10] & ~io_in[11]) | (io_in[0] & ~io_in[1] & ~io_in[4] & io_in[6] & io_in[7] & ~io_in[8] & io_in[9] & io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[4] & ~io_in[5] & ~io_in[6] & io_in[7] & ~io_in[8] & ~io_in[9] & ~io_in[10]) | (io_in[0] & ~io_in[1] & ~io_in[3] & io_in[5] & io_in[6] & io_in[7] & ~io_in[8] & io_in[10]) | (~io_in[0] & io_in[1] & ~io_in[3] & io_in[4] & io_in[7] & ~io_in[8] & ~io_in[9] & ~io_in[11]) | (~io_in[1] & ~io_in[2] & io_in[4] & ~io_in[6] & io_in[7] & ~io_in[8] & io_in[9] & io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & io_in[3] & io_in[6] & ~io_in[9] & io_in[11]) | (~io_in[1] & io_in[2] & ~io_in[3] & io_in[6] & io_in[8] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (io_in[0] & ~io_in[2] & io_in[4] & ~io_in[6] & io_in[7] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[1] & io_in[2] & io_in[5] & ~io_in[6] & ~io_in[9] & io_in[10]) | (io_in[0] & ~io_in[1] & ~io_in[2] & io_in[3] & ~io_in[4] & ~io_in[6] & io_in[7] & ~io_in[10] & ~io_in[11]) | (io_in[2] & io_in[3] & ~io_in[4] & ~io_in[6] & io_in[7] & ~io_in[8] & io_in[9] & ~io_in[10]) | (~io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & io_in[4] & io_in[6] & io_in[7] & io_in[8]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & io_in[5] & io_in[6] & ~io_in[8] & io_in[9]) | (~io_in[0] & io_in[1] & ~io_in[2] & io_in[4] & io_in[7] & ~io_in[8] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[3] & ~io_in[6] & io_in[7] & ~io_in[8] & ~io_in[9] & io_in[10] & ~io_in[11]) | (io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[7] & io_in[9] & io_in[10]) | (io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[7] & ~io_in[8] & io_in[9] & ~io_in[11]) | (io_in[0] & ~io_in[2] & ~io_in[3] & io_in[4] & io_in[6] & ~io_in[7] & ~io_in[10] & io_in[11]) | (io_in[0] & io_in[1] & ~io_in[2] & io_in[3] & io_in[6] & ~io_in[7] & io_in[8] & ~io_in[10]) | (io_in[0] & io_in[2] & ~io_in[4] & ~io_in[5] & io_in[6] & io_in[7] & io_in[8] & ~io_in[9] & io_in[11]) | (io_in[0] & io_in[1] & io_in[3] & ~io_in[6] & ~io_in[7] & ~io_in[8] & ~io_in[9]) | (io_in[1] & io_in[2] & ~io_in[3] & io_in[4] & ~io_in[7] & ~io_in[8] & ~io_in[9] & io_in[10]) | (~io_in[0] & io_in[3] & io_in[6] & io_in[7] & io_in[8] & ~io_in[9] & io_in[11]) | (~io_in[0] & ~io_in[3] & io_in[4] & ~io_in[6] & io_in[7] & io_in[8] & io_in[9] & io_in[10] & ~io_in[11]) | (io_in[0] & ~io_in[1] & ~io_in[2] & io_in[4] & ~io_in[7] & io_in[9] & ~io_in[10] & io_in[11]) | (io_in[2] & io_in[3] & io_in[4] & ~io_in[7] & ~io_in[8] & ~io_in[10] & ~io_in[11]) | (io_in[0] & ~io_in[3] & io_in[4] & ~io_in[6] & io_in[7] & ~io_in[8] & ~io_in[9] & io_in[11]) | (io_in[1] & io_in[4] & io_in[6] & io_in[7] & io_in[9] & ~io_in[10] & io_in[11]) | (~io_in[0] & io_in[1] & io_in[2] & ~io_in[4] & io_in[6] & ~io_in[7] & io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & io_in[1] & ~io_in[4] & ~io_in[5] & io_in[6] & io_in[7] & ~io_in[8] & io_in[9] & io_in[10]) | (~io_in[0] & ~io_in[1] & io_in[2] & io_in[4] & ~io_in[7] & ~io_in[8] & ~io_in[10] & ~io_in[11]) | (io_in[0] & ~io_in[1] & io_in[3] & ~io_in[4] & io_in[7] & io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & ~io_in[2] & io_in[4] & ~io_in[6] & io_in[7] & io_in[8] & ~io_in[9] & io_in[10]) | (~io_in[0] & io_in[2] & ~io_in[3] & ~io_in[4] & io_in[6] & ~io_in[7] & io_in[8] & ~io_in[10] & io_in[11]) | (io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & io_in[7] & ~io_in[9] & io_in[11]) | (io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[7] & ~io_in[9] & ~io_in[11]) | (io_in[0] & io_in[1] & io_in[2] & ~io_in[5] & ~io_in[6] & ~io_in[7] & ~io_in[8] & io_in[9] & io_in[11]) | (io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[4] & ~io_in[6] & io_in[7] & io_in[10] & io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[5] & ~io_in[6] & ~io_in[7] & ~io_in[9] & ~io_in[11]) | (~io_in[0] & ~io_in[2] & ~io_in[3] & ~io_in[5] & ~io_in[6] & ~io_in[7] & ~io_in[8] & io_in[9] & ~io_in[10] & io_in[11]) | (io_in[0] & io_in[1] & io_in[2] & ~io_in[3] & io_in[4] & io_in[7] & io_in[8] & io_in[9] & io_in[10]) | (~io_in[0] & io_in[1] & io_in[3] & ~io_in[4] & io_in[6] & ~io_in[7] & io_in[8] & io_in[9] & io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[2] & io_in[3] & ~io_in[4] & io_in[6] & io_in[8] & io_in[9] & io_in[10] & ~io_in[11]) | (io_in[0] & ~io_in[1] & io_in[2] & ~io_in[4] & ~io_in[5] & ~io_in[6] & io_in[7] & ~io_in[8] & io_in[9]) | (io_in[1] & ~io_in[2] & io_in[5] & io_in[7] & io_in[8] & io_in[9] & io_in[10] & ~io_in[11]) | (io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & ~io_in[5] & io_in[6] & io_in[7] & io_in[8] & io_in[9] & ~io_in[10]) | (io_in[0] & ~io_in[1] & io_in[3] & io_in[4] & io_in[6] & ~io_in[8] & io_in[11]) | (~io_in[0] & io_in[1] & io_in[2] & ~io_in[3] & ~io_in[5] & io_in[6] & ~io_in[8] & ~io_in[9] & io_in[11]) | (~io_in[0] & io_in[1] & io_in[2] & io_in[3] & ~io_in[6] & ~io_in[8] & ~io_in[9] & io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[7] & io_in[8] & io_in[10] & ~io_in[11]) | (~io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & io_in[6] & ~io_in[7] & io_in[8] & io_in[9] & ~io_in[11]) | (~io_in[0] & io_in[1] & io_in[2] & ~io_in[3] & io_in[4] & ~io_in[5] & io_in[7] & io_in[9] & io_in[11]) | (~io_in[0] & io_in[2] & io_in[3] & io_in[4] & io_in[6] & ~io_in[7] & io_in[9] & io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & io_in[5] & io_in[7] & ~io_in[9] & ~io_in[10]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & io_in[7] & ~io_in[8] & ~io_in[10] & ~io_in[11]) | (io_in[1] & io_in[2] & ~io_in[3] & io_in[5] & ~io_in[6] & io_in[7] & ~io_in[8] & ~io_in[9] & io_in[10]) | (~io_in[0] & io_in[1] & io_in[2] & io_in[5] & io_in[6] & io_in[9] & ~io_in[10]) | (io_in[0] & io_in[2] & ~io_in[3] & ~io_in[5] & io_in[6] & io_in[7] & ~io_in[8] & io_in[9] & io_in[10]) | (io_in[0] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[6] & ~io_in[7] & ~io_in[8] & ~io_in[9]) | (io_in[0] & io_in[1] & ~io_in[3] & io_in[5] & io_in[6] & ~io_in[7] & io_in[11]) | (io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & io_in[4] & ~io_in[6] & ~io_in[7] & io_in[8] & io_in[10]) | (~io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & io_in[4] & ~io_in[6] & io_in[8] & io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[7] & ~io_in[8] & ~io_in[11]) | (~io_in[0] & ~io_in[2] & io_in[5] & io_in[6] & io_in[8] & io_in[11]) | (~io_in[0] & io_in[2] & io_in[3] & ~io_in[4] & io_in[6] & ~io_in[7] & io_in[8] & io_in[9] & ~io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[8] & io_in[9] & ~io_in[10] & ~io_in[11]) | (io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & ~io_in[5] & io_in[7] & ~io_in[9] & io_in[10]) | (~io_in[0] & ~io_in[1] & io_in[5] & ~io_in[6] & io_in[7] & io_in[9] & ~io_in[10]) | (~io_in[0] & ~io_in[2] & io_in[4] & ~io_in[5] & io_in[6] & io_in[7] & io_in[8] & ~io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & io_in[5] & ~io_in[7] & io_in[8] & ~io_in[10]) | (io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & io_in[6] & ~io_in[7] & ~io_in[10]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & io_in[4] & io_in[6] & io_in[7] & ~io_in[9] & io_in[11]) | (io_in[0] & io_in[1] & ~io_in[2] & ~io_in[4] & io_in[6] & io_in[7] & io_in[8] & io_in[9] & ~io_in[10]) | (~io_in[0] & io_in[1] & io_in[2] & ~io_in[3] & io_in[4] & io_in[6] & ~io_in[7] & io_in[9] & ~io_in[11]) | (io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[7] & io_in[8] & io_in[10]) | (io_in[0] & ~io_in[2] & io_in[3] & ~io_in[4] & io_in[6] & io_in[7] & io_in[9] & io_in[11]) | (io_in[1] & io_in[2] & io_in[3] & ~io_in[6] & io_in[7] & io_in[8] & io_in[9] & ~io_in[11]) | (io_in[0] & ~io_in[1] & io_in[2] & ~io_in[4] & ~io_in[5] & io_in[6] & ~io_in[7] & ~io_in[8] & io_in[10]) | (~io_in[0] & io_in[1] & io_in[2] & ~io_in[3] & io_in[4] & io_in[7] & io_in[8] & ~io_in[10]) | (io_in[1] & ~io_in[2] & io_in[3] & io_in[4] & ~io_in[6] & io_in[7] & io_in[8] & io_in[11]) | (~io_in[0] & ~io_in[1] & io_in[4] & ~io_in[6] & ~io_in[7] & io_in[8] & ~io_in[9] & io_in[10]) | (~io_in[0] & io_in[2] & io_in[3] & io_in[4] & io_in[6] & ~io_in[8] & io_in[9] & io_in[10]) | (~io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & ~io_in[6] & ~io_in[7] & ~io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & io_in[1] & io_in[2] & io_in[3] & ~io_in[7] & ~io_in[8] & ~io_in[10]) | (io_in[0] & ~io_in[1] & io_in[4] & io_in[6] & io_in[7] & ~io_in[8] & io_in[9] & io_in[10]) | (~io_in[0] & ~io_in[1] & io_in[2] & ~io_in[4] & ~io_in[6] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & ~io_in[2] & io_in[3] & io_in[4] & ~io_in[5] & ~io_in[6] & ~io_in[7] & io_in[10] & io_in[11]) | (~io_in[0] & ~io_in[1] & io_in[3] & io_in[5] & ~io_in[7] & ~io_in[8]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[4] & ~io_in[5] & io_in[7] & ~io_in[8] & ~io_in[9] & io_in[10] & ~io_in[11]) | (io_in[0] & io_in[1] & io_in[3] & io_in[5] & ~io_in[6] & ~io_in[7]) | (~io_in[0] & ~io_in[1] & io_in[2] & ~io_in[4] & ~io_in[5] & ~io_in[6] & io_in[10] & io_in[11]) | (~io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & io_in[5] & ~io_in[7]) | (~io_in[0] & ~io_in[1] & io_in[2] & io_in[4] & io_in[6] & io_in[7] & io_in[9] & io_in[11]) | (~io_in[0] & io_in[1] & io_in[2] & ~io_in[4] & ~io_in[6] & ~io_in[7] & ~io_in[8] & ~io_in[9] & io_in[11]) | (~io_in[0] & io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & ~io_in[6] & io_in[7] & io_in[10]) | (io_in[0] & ~io_in[1] & ~io_in[3] & ~io_in[5] & io_in[6] & ~io_in[7] & ~io_in[8] & io_in[9]) | (~io_in[0] & io_in[1] & ~io_in[3] & io_in[4] & io_in[8] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (io_in[0] & ~io_in[1] & io_in[3] & ~io_in[4] & ~io_in[6] & ~io_in[7] & ~io_in[8] & io_in[9]) | (io_in[0] & io_in[1] & ~io_in[2] & io_in[3] & ~io_in[4] & ~io_in[6] & io_in[9] & io_in[10] & ~io_in[11]) | (io_in[0] & io_in[1] & io_in[2] & ~io_in[3] & io_in[4] & io_in[6] & ~io_in[7] & ~io_in[9]) | (~io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & io_in[6] & ~io_in[7] & io_in[8] & ~io_in[9] & ~io_in[10]) | (io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & io_in[6] & io_in[7] & ~io_in[9] & io_in[10]) | (io_in[0] & io_in[3] & ~io_in[4] & ~io_in[6] & io_in[8] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & ~io_in[2] & ~io_in[3] & ~io_in[6] & ~io_in[7] & io_in[8] & io_in[9] & ~io_in[11]) | (~io_in[0] & io_in[2] & io_in[3] & ~io_in[4] & ~io_in[6] & ~io_in[7] & ~io_in[8] & io_in[9] & io_in[10]) | (~io_in[0] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & io_in[7] & ~io_in[8] & ~io_in[10] & io_in[11]) | (~io_in[0] & io_in[2] & io_in[3] & ~io_in[4] & ~io_in[5] & io_in[7] & ~io_in[10] & io_in[11]) | (~io_in[1] & ~io_in[2] & io_in[5] & io_in[6] & ~io_in[7] & io_in[8] & io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[4] & ~io_in[5] & ~io_in[6] & io_in[7] & io_in[9] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[6] & ~io_in[7] & io_in[8] & ~io_in[11]) | (io_in[0] & io_in[1] & ~io_in[2] & io_in[3] & ~io_in[4] & ~io_in[6] & ~io_in[8] & io_in[10]) | (~io_in[0] & io_in[1] & ~io_in[2] & io_in[3] & ~io_in[6] & io_in[7] & io_in[9] & ~io_in[10]) | (io_in[1] & ~io_in[3] & ~io_in[4] & ~io_in[8] & io_in[9] & ~io_in[10] & ~io_in[11]) | (~io_in[1] & ~io_in[3] & io_in[5] & ~io_in[7] & io_in[8] & ~io_in[9] & io_in[10]) | (~io_in[0] & ~io_in[1] & io_in[2] & io_in[5] & io_in[7] & ~io_in[8] & ~io_in[9] & io_in[10]) | (~io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & io_in[4] & ~io_in[8] & io_in[9] & ~io_in[10] & ~io_in[11]) | (io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & io_in[5] & ~io_in[7] & io_in[8] & io_in[11]) | (~io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & ~io_in[6] & ~io_in[7] & ~io_in[8] & io_in[9]) | (~io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & ~io_in[6] & ~io_in[9] & ~io_in[11]) | (io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & io_in[7] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[3] & io_in[5] & ~io_in[7] & ~io_in[8] & ~io_in[9] & io_in[10]) | (~io_in[0] & io_in[1] & ~io_in[3] & ~io_in[4] & io_in[5] & ~io_in[6] & ~io_in[7] & io_in[10] & io_in[11]) | (~io_in[0] & io_in[2] & ~io_in[3] & io_in[4] & ~io_in[5] & io_in[7] & io_in[10] & io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[3] & ~io_in[6] & io_in[7] & io_in[8] & ~io_in[10] & io_in[11]) | (io_in[0] & ~io_in[2] & io_in[3] & io_in[4] & ~io_in[6] & io_in[7] & io_in[8] & ~io_in[9]) | (~io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & io_in[7] & ~io_in[8] & ~io_in[9] & io_in[10]) | (~io_in[0] & io_in[2] & ~io_in[4] & ~io_in[5] & ~io_in[6] & io_in[7] & io_in[8] & ~io_in[9]) | (io_in[0] & ~io_in[1] & ~io_in[2] & io_in[4] & io_in[6] & ~io_in[7] & io_in[9] & ~io_in[10]) | (~io_in[0] & io_in[1] & ~io_in[3] & ~io_in[5] & ~io_in[6] & ~io_in[7] & io_in[8] & io_in[9] & io_in[10] & ~io_in[11]) | (~io_in[0] & ~io_in[2] & io_in[4] & io_in[6] & ~io_in[7] & ~io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & ~io_in[2] & ~io_in[3] & io_in[4] & io_in[6] & ~io_in[7] & io_in[9] & io_in[10] & ~io_in[11]) | (io_in[0] & io_in[1] & ~io_in[2] & io_in[3] & ~io_in[4] & ~io_in[5] & io_in[7] & ~io_in[8] & io_in[10]) | (~io_in[0] & io_in[1] & ~io_in[2] & io_in[4] & io_in[6] & io_in[8] & ~io_in[9] & ~io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & io_in[4] & io_in[6] & io_in[7] & io_in[8] & io_in[9]) | (~io_in[0] & ~io_in[2] & io_in[3] & io_in[4] & io_in[6] & io_in[7] & io_in[9] & ~io_in[10]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & io_in[3] & io_in[8] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[5] & io_in[6] & io_in[7] & ~io_in[8] & ~io_in[9]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[6] & io_in[8] & io_in[10] & ~io_in[11]) | (io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[7] & io_in[8] & ~io_in[10]) | (io_in[0] & io_in[2] & io_in[3] & io_in[5] & ~io_in[8] & io_in[9]) | (~io_in[1] & ~io_in[2] & io_in[3] & io_in[6] & ~io_in[7] & ~io_in[8] & ~io_in[9] & io_in[10]) | (~io_in[0] & ~io_in[1] & io_in[2] & io_in[4] & ~io_in[6] & ~io_in[8] & ~io_in[10] & ~io_in[11]) | (io_in[1] & ~io_in[2] & io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & ~io_in[8] & io_in[9] & io_in[10]) | (io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[7] & ~io_in[8] & ~io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & io_in[3] & ~io_in[4] & ~io_in[6] & ~io_in[8] & io_in[11]) | (~io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & ~io_in[7] & io_in[8] & io_in[9] & ~io_in[10]) | (io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & io_in[5] & io_in[6] & io_in[7] & io_in[10] & ~io_in[11]) | (~io_in[0] & ~io_in[1] & io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & io_in[9] & ~io_in[10] & ~io_in[11]) | (io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & io_in[8] & io_in[10] & ~io_in[11]) | (io_in[0] & ~io_in[1] & ~io_in[3] & io_in[4] & io_in[6] & io_in[7] & ~io_in[8] & ~io_in[9] & ~io_in[11]) | (io_in[0] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[6] & ~io_in[7] & io_in[8] & io_in[9] & ~io_in[10]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & io_in[3] & ~io_in[7] & ~io_in[8] & ~io_in[9] & io_in[11]) | (io_in[0] & ~io_in[2] & ~io_in[3] & io_in[5] & ~io_in[8] & ~io_in[9] & io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & io_in[3] & io_in[4] & io_in[6] & io_in[8] & ~io_in[11]) | (io_in[0] & ~io_in[1] & ~io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[7] & ~io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & ~io_in[3] & ~io_in[4] & ~io_in[6] & ~io_in[8] & io_in[9] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[2] & io_in[3] & io_in[4] & io_in[7] & ~io_in[8] & io_in[9] & io_in[10]) | (io_in[0] & io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[7] & io_in[8] & ~io_in[9] & io_in[10]) | (~io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & io_in[6] & ~io_in[8] & io_in[11]) | (~io_in[0] & io_in[1] & io_in[2] & ~io_in[4] & ~io_in[5] & io_in[6] & ~io_in[7] & io_in[10] & io_in[11]) | (io_in[0] & io_in[1] & io_in[3] & io_in[4] & io_in[6] & io_in[7] & ~io_in[8] & ~io_in[10]) | (~io_in[0] & io_in[1] & io_in[2] & io_in[3] & io_in[4] & ~io_in[6] & ~io_in[7] & ~io_in[9]) | (~io_in[0] & ~io_in[1] & io_in[2] & ~io_in[4] & ~io_in[5] & io_in[6] & io_in[7] & io_in[8] & io_in[9] & io_in[10] & ~io_in[11]) | (io_in[0] & io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & ~io_in[6] & ~io_in[7] & ~io_in[9]) | (io_in[0] & io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & ~io_in[6] & ~io_in[8] & io_in[11]) | (io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[6] & io_in[8] & ~io_in[10] & io_in[11]) | (~io_in[0] & ~io_in[1] & io_in[4] & ~io_in[6] & ~io_in[7] & io_in[8] & io_in[9] & ~io_in[10]) | (io_in[0] & io_in[2] & ~io_in[4] & ~io_in[6] & io_in[7] & ~io_in[8] & io_in[9] & ~io_in[10]) | (io_in[0] & io_in[1] & ~io_in[2] & io_in[3] & ~io_in[5] & ~io_in[6] & ~io_in[9] & io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[4] & io_in[5] & io_in[6] & ~io_in[7] & io_in[10]) | (~io_in[1] & io_in[4] & io_in[6] & io_in[8] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (io_in[0] & ~io_in[1] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[7] & io_in[9] & io_in[11]) | (io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & ~io_in[6] & ~io_in[8] & ~io_in[9] & ~io_in[10]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[7] & io_in[8] & io_in[9] & ~io_in[10] & ~io_in[11]) | (io_in[0] & io_in[1] & ~io_in[4] & ~io_in[6] & io_in[7] & io_in[8] & io_in[9] & io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & io_in[6] & io_in[7] & ~io_in[9] & ~io_in[10]) | (io_in[0] & io_in[1] & ~io_in[2] & io_in[3] & io_in[6] & ~io_in[7] & ~io_in[8] & io_in[9] & io_in[10]) | (io_in[0] & ~io_in[1] & io_in[2] & io_in[4] & io_in[6] & io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & ~io_in[5] & io_in[7] & io_in[8] & io_in[10] & ~io_in[11]) | (io_in[0] & ~io_in[2] & ~io_in[3] & ~io_in[4] & io_in[5] & ~io_in[6] & io_in[10] & io_in[11]) | (~io_in[0] & io_in[2] & ~io_in[4] & io_in[6] & io_in[7] & ~io_in[8] & ~io_in[9] & io_in[11]) | (io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[6] & ~io_in[7] & ~io_in[8]) | (~io_in[0] & io_in[2] & io_in[5] & io_in[6] & ~io_in[7] & ~io_in[11]) | (~io_in[0] & io_in[2] & io_in[3] & io_in[4] & io_in[6] & io_in[7] & ~io_in[8] & io_in[10]) | (io_in[0] & io_in[2] & io_in[3] & io_in[4] & ~io_in[6] & io_in[8] & ~io_in[10] & ~io_in[11]) | (~io_in[1] & io_in[2] & io_in[4] & io_in[5] & ~io_in[6]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & io_in[3] & ~io_in[6] & io_in[7] & ~io_in[8] & io_in[9] & io_in[10]) | (~io_in[0] & ~io_in[2] & io_in[4] & ~io_in[6] & ~io_in[7] & ~io_in[8] & io_in[9] & io_in[10]) | (io_in[1] & ~io_in[2] & io_in[3] & ~io_in[4] & io_in[6] & ~io_in[7] & ~io_in[8] & io_in[9]) | (io_in[0] & ~io_in[1] & ~io_in[2] & io_in[3] & io_in[5] & io_in[6] & ~io_in[9]) | (io_in[0] & ~io_in[1] & ~io_in[2] & io_in[3] & ~io_in[5] & io_in[6] & ~io_in[7] & io_in[9] & io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & ~io_in[6] & io_in[8] & ~io_in[9] & io_in[11]) | (io_in[1] & io_in[3] & io_in[5] & io_in[8] & io_in[10] & ~io_in[11]) | (~io_in[1] & ~io_in[2] & io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[6] & io_in[7] & ~io_in[8] & ~io_in[9]) | (io_in[0] & io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[7] & io_in[8] & io_in[9] & ~io_in[10]) | (io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & ~io_in[7] & io_in[8] & io_in[9] & io_in[10] & ~io_in[11]) | (io_in[1] & io_in[2] & io_in[4] & ~io_in[6] & ~io_in[7] & io_in[8] & ~io_in[9] & io_in[11]) | (io_in[0] & io_in[2] & ~io_in[3] & io_in[6] & io_in[7] & io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & io_in[1] & io_in[2] & io_in[3] & ~io_in[7] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[2] & ~io_in[3] & io_in[5] & io_in[7] & ~io_in[8] & io_in[10]) | (io_in[0] & io_in[1] & ~io_in[2] & ~io_in[4] & io_in[6] & io_in[8] & ~io_in[9] & ~io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[5] & ~io_in[6] & io_in[10] & io_in[11]) | (~io_in[0] & ~io_in[1] & io_in[5] & ~io_in[7] & io_in[9] & ~io_in[11]) | (io_in[0] & io_in[2] & io_in[3] & io_in[4] & ~io_in[6] & ~io_in[7] & io_in[9] & ~io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & io_in[4] & ~io_in[5] & ~io_in[6] & io_in[8] & io_in[9] & io_in[10]) | (io_in[0] & io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[7] & ~io_in[8] & ~io_in[9] & ~io_in[11]) | (io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & ~io_in[6] & ~io_in[7] & io_in[8] & io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[4] & ~io_in[5] & ~io_in[6] & ~io_in[7] & io_in[8] & io_in[11]) | (io_in[0] & io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & io_in[6] & io_in[10] & io_in[11]) | (io_in[0] & io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & io_in[7] & io_in[9] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[1] & io_in[2] & io_in[3] & io_in[4] & ~io_in[8] & io_in[10]) | (~io_in[1] & ~io_in[2] & io_in[3] & io_in[4] & io_in[6] & ~io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & io_in[6] & io_in[7] & ~io_in[8] & ~io_in[11]) | (io_in[0] & io_in[2] & io_in[3] & io_in[4] & ~io_in[6] & io_in[7] & io_in[8] & io_in[9]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[7] & io_in[10] & io_in[11]) | (~io_in[0] & io_in[1] & io_in[2] & io_in[4] & io_in[6] & ~io_in[7] & io_in[9] & ~io_in[10]) | (~io_in[0] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[6] & io_in[8] & io_in[9] & io_in[10] & io_in[11]) | (io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & ~io_in[6] & io_in[8] & io_in[9] & ~io_in[10]) | (~io_in[2] & io_in[3] & io_in[4] & io_in[7] & io_in[9] & ~io_in[10] & io_in[11]) | (io_in[0] & ~io_in[2] & ~io_in[3] & ~io_in[4] & io_in[6] & ~io_in[7] & io_in[8] & ~io_in[9]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & io_in[3] & ~io_in[4] & ~io_in[5] & io_in[7] & ~io_in[9]) | (~io_in[0] & io_in[1] & io_in[3] & ~io_in[5] & ~io_in[6] & io_in[7] & ~io_in[8] & ~io_in[9] & io_in[10]) | (~io_in[0] & ~io_in[1] & io_in[3] & io_in[5] & ~io_in[7] & io_in[11]) | (io_in[0] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & io_in[7] & io_in[8] & ~io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & io_in[3] & io_in[5] & io_in[6] & io_in[10]) | (~io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & io_in[4] & ~io_in[8] & io_in[9] & io_in[11]) | (~io_in[0] & io_in[2] & io_in[3] & ~io_in[7] & ~io_in[8] & ~io_in[10] & ~io_in[11]) | (io_in[0] & io_in[1] & io_in[2] & ~io_in[3] & io_in[6] & ~io_in[7] & ~io_in[9] & io_in[10]) | (io_in[0] & io_in[1] & ~io_in[2] & io_in[3] & io_in[6] & io_in[7] & ~io_in[8] & io_in[11]) | (io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & io_in[6] & ~io_in[7] & ~io_in[9] & io_in[11]) | (io_in[0] & io_in[1] & io_in[2] & io_in[3] & io_in[4] & ~io_in[6] & io_in[7] & io_in[8]) | (io_in[0] & io_in[1] & io_in[2] & ~io_in[8] & io_in[9] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & io_in[5] & io_in[8] & ~io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & io_in[3] & ~io_in[4] & ~io_in[6] & io_in[9] & ~io_in[10]) | (io_in[0] & io_in[3] & io_in[5] & io_in[9] & ~io_in[10]) | (io_in[1] & io_in[2] & ~io_in[4] & ~io_in[7] & ~io_in[8] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & ~io_in[2] & io_in[3] & ~io_in[5] & io_in[6] & ~io_in[7] & ~io_in[8] & ~io_in[9] & io_in[11]) | (~io_in[1] & ~io_in[2] & io_in[3] & ~io_in[5] & io_in[6] & io_in[7] & io_in[8] & io_in[9] & io_in[10] & ~io_in[11]) | (io_in[0] & io_in[1] & ~io_in[5] & ~io_in[6] & ~io_in[7] & io_in[8] & ~io_in[9] & io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & io_in[3] & ~io_in[4] & io_in[6] & ~io_in[9] & ~io_in[10]) | (~io_in[0] & ~io_in[2] & ~io_in[3] & io_in[6] & ~io_in[7] & io_in[8] & io_in[9] & io_in[10] & io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & io_in[3] & io_in[6] & ~io_in[7] & ~io_in[8] & io_in[10]) | (io_in[0] & ~io_in[1] & ~io_in[3] & io_in[4] & ~io_in[5] & io_in[6] & io_in[10] & io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[3] & io_in[4] & ~io_in[5] & ~io_in[6] & io_in[7] & io_in[9] & io_in[10]) | (~io_in[0] & io_in[3] & ~io_in[4] & io_in[6] & io_in[7] & ~io_in[9] & io_in[11]) | (io_in[0] & io_in[1] & ~io_in[2] & io_in[4] & ~io_in[6] & io_in[8] & ~io_in[9] & io_in[10]) | (~io_in[0] & ~io_in[1] & io_in[2] & ~io_in[4] & io_in[5] & io_in[6] & io_in[11]) | (io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & io_in[4] & io_in[8] & ~io_in[9] & ~io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[5] & io_in[6] & io_in[9] & io_in[11]) | (io_in[0] & io_in[1] & io_in[2] & ~io_in[3] & ~io_in[5] & io_in[7] & io_in[10] & io_in[11]) | (io_in[0] & io_in[1] & ~io_in[2] & io_in[3] & io_in[6] & ~io_in[7] & io_in[8] & ~io_in[9]) | (io_in[0] & io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[8] & ~io_in[10] & ~io_in[11]) | (~io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[6] & ~io_in[7] & io_in[8] & io_in[9] & io_in[10] & ~io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[4] & io_in[6] & ~io_in[7] & ~io_in[9] & ~io_in[10] & io_in[11]) | (io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & ~io_in[5] & ~io_in[6] & io_in[7] & ~io_in[9] & io_in[10]) | (io_in[0] & ~io_in[1] & ~io_in[2] & io_in[5] & ~io_in[6] & io_in[7] & io_in[9] & ~io_in[11]) | (~io_in[0] & ~io_in[1] & io_in[2] & io_in[4] & ~io_in[6] & ~io_in[7] & ~io_in[8] & io_in[11]) | (~io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & ~io_in[7] & ~io_in[8] & io_in[10]) | (~io_in[1] & ~io_in[2] & ~io_in[4] & ~io_in[5] & ~io_in[6] & io_in[7] & ~io_in[9] & io_in[10] & ~io_in[11]) | (io_in[0] & ~io_in[1] & io_in[2] & io_in[5] & ~io_in[6] & io_in[8] & ~io_in[9]) | (~io_in[0] & io_in[1] & io_in[2] & io_in[5] & ~io_in[6] & ~io_in[8]) | (io_in[0] & io_in[1] & ~io_in[2] & io_in[3] & ~io_in[6] & io_in[7] & io_in[9] & io_in[10] & ~io_in[11]) | (io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[7] & ~io_in[9] & ~io_in[10]) | (~io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & io_in[4] & io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & io_in[1] & io_in[2] & io_in[3] & ~io_in[6] & io_in[7] & io_in[9] & ~io_in[10]) | (~io_in[0] & io_in[1] & io_in[5] & io_in[7] & io_in[8] & ~io_in[9] & io_in[10]) | (~io_in[1] & io_in[2] & ~io_in[3] & ~io_in[5] & io_in[6] & io_in[7] & io_in[10] & io_in[11]) | (io_in[0] & io_in[2] & ~io_in[3] & ~io_in[6] & ~io_in[8] & io_in[9] & ~io_in[10] & ~io_in[11]) | (io_in[0] & io_in[1] & io_in[4] & io_in[5] & io_in[7]) | (io_in[0] & io_in[1] & io_in[2] & io_in[3] & ~io_in[6] & ~io_in[7] & io_in[11]) | (~io_in[0] & io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[6] & io_in[7] & ~io_in[8] & io_in[11]);

assign val[1] = (io_in[1] & io_in[3] & io_in[4] & io_in[6] & io_in[7] & io_in[10] & io_in[11]) | (~io_in[0] & io_in[1] & io_in[2] & io_in[6] & io_in[7] & ~io_in[8] & io_in[9] & io_in[11]) | (io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & io_in[6] & ~io_in[7] & ~io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & io_in[2] & io_in[3] & ~io_in[4] & io_in[6] & io_in[7] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (io_in[0] & io_in[1] & io_in[2] & io_in[3] & io_in[4] & io_in[9] & ~io_in[10]) | (~io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & ~io_in[6] & ~io_in[7] & io_in[8] & ~io_in[10] & io_in[11]) | (io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & io_in[7] & io_in[8] & io_in[9] & ~io_in[11]) | (~io_in[0] & io_in[2] & io_in[3] & ~io_in[4] & io_in[6] & ~io_in[7] & io_in[8] & io_in[9] & ~io_in[10]) | (io_in[0] & io_in[2] & io_in[4] & ~io_in[6] & ~io_in[7] & io_in[8] & io_in[9] & ~io_in[10]) | (io_in[0] & io_in[1] & ~io_in[2] & io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & io_in[8] & io_in[9] & ~io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & io_in[3] & io_in[6] & ~io_in[7] & ~io_in[8] & io_in[9] & io_in[10]) | (~io_in[0] & io_in[1] & io_in[2] & ~io_in[3] & io_in[4] & io_in[7] & io_in[8] & io_in[9] & io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[4] & ~io_in[5] & ~io_in[7] & ~io_in[8] & io_in[9] & io_in[10]) | (~io_in[0] & io_in[1] & io_in[2] & io_in[3] & ~io_in[7] & ~io_in[8] & io_in[9] & io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & io_in[3] & ~io_in[5] & io_in[6] & io_in[7] & ~io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & ~io_in[1] & ~io_in[2] & io_in[3] & ~io_in[4] & io_in[6] & io_in[7] & ~io_in[9] & io_in[10]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[6] & ~io_in[7] & ~io_in[10]) | (io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & ~io_in[6] & io_in[7] & ~io_in[8] & io_in[9] & io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & io_in[4] & ~io_in[5] & ~io_in[6] & ~io_in[7] & io_in[10] & io_in[11]) | (io_in[0] & io_in[1] & io_in[2] & io_in[3] & io_in[4] & ~io_in[6] & ~io_in[8] & io_in[11]) | (~io_in[1] & io_in[3] & ~io_in[4] & ~io_in[6] & ~io_in[7] & ~io_in[8] & io_in[9] & io_in[10]) | (io_in[0] & ~io_in[1] & ~io_in[2] & io_in[3] & io_in[4] & ~io_in[6] & io_in[7] & ~io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & io_in[5] & io_in[6] & ~io_in[7] & io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[3] & io_in[4] & io_in[6] & ~io_in[8] & io_in[9] & io_in[10]) | (io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & ~io_in[7] & ~io_in[8] & ~io_in[9] & io_in[11]) | (io_in[0] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[7] & io_in[8] & io_in[9] & io_in[10] & ~io_in[11]) | (io_in[1] & ~io_in[2] & io_in[3] & io_in[4] & io_in[6] & ~io_in[7] & io_in[8] & io_in[9] & ~io_in[10]) | (io_in[0] & io_in[1] & ~io_in[3] & ~io_in[6] & io_in[7] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & io_in[4] & io_in[6] & ~io_in[7] & io_in[8] & io_in[9] & ~io_in[11]) | (io_in[0] & ~io_in[1] & ~io_in[2] & io_in[3] & ~io_in[4] & ~io_in[6] & io_in[7] & ~io_in[8] & io_in[9] & ~io_in[10]) | (io_in[0] & io_in[2] & io_in[3] & io_in[4] & ~io_in[8] & io_in[9] & ~io_in[10] & ~io_in[11]) | (io_in[0] & ~io_in[1] & io_in[2] & io_in[5] & io_in[7] & io_in[8] & ~io_in[10]) | (~io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & io_in[4] & ~io_in[7] & ~io_in[8] & io_in[9] & io_in[10]) | (~io_in[0] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & io_in[7] & ~io_in[8] & io_in[9] & io_in[10] & ~io_in[11]) | (~io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & ~io_in[8] & io_in[9] & ~io_in[10] & io_in[11]) | (io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[6] & io_in[7] & io_in[8] & ~io_in[9]) | (~io_in[0] & io_in[2] & ~io_in[3] & io_in[6] & ~io_in[7] & io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & io_in[9] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & io_in[3] & io_in[5] & io_in[6] & io_in[9] & io_in[11]) | (~io_in[0] & ~io_in[2] & io_in[3] & io_in[4] & ~io_in[6] & io_in[8] & ~io_in[10] & io_in[11]) | (io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[7] & io_in[10] & io_in[11]) | (io_in[0] & io_in[2] & io_in[4] & ~io_in[6] & ~io_in[7] & ~io_in[8] & ~io_in[9] & io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & io_in[6] & ~io_in[7] & ~io_in[8] & ~io_in[9] & io_in[10]) | (io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[6] & ~io_in[7] & io_in[9] & io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[2] & ~io_in[3] & io_in[4] & ~io_in[6] & io_in[8] & io_in[9] & io_in[10] & ~io_in[11]) | (~io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & io_in[4] & ~io_in[6] & io_in[7] & io_in[8] & io_in[11]) | (io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[5] & io_in[7] & io_in[10] & io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[3] & io_in[5] & io_in[6] & io_in[7] & ~io_in[9] & io_in[10]) | (io_in[0] & io_in[5] & io_in[7] & io_in[9] & ~io_in[10] & io_in[11]) | (io_in[0] & ~io_in[2] & io_in[3] & ~io_in[4] & io_in[6] & ~io_in[7] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (io_in[0] & ~io_in[1] & io_in[2] & io_in[4] & io_in[6] & io_in[7] & ~io_in[9] & io_in[10]) | (~io_in[0] & ~io_in[1] & io_in[2] & io_in[6] & io_in[7] & io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & io_in[5] & io_in[6] & io_in[7] & ~io_in[8]) | (io_in[0] & ~io_in[1] & ~io_in[2] & io_in[3] & io_in[6] & io_in[7] & io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & ~io_in[1] & io_in[2] & ~io_in[4] & ~io_in[6] & ~io_in[7] & io_in[10] & io_in[11]) | (io_in[0] & ~io_in[2] & io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[6] & io_in[10] & io_in[11]) | (~io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & ~io_in[5] & io_in[6] & ~io_in[7] & ~io_in[8] & ~io_in[9] & io_in[11]) | (~io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & io_in[7] & ~io_in[8] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[4] & ~io_in[5] & io_in[6] & ~io_in[7] & ~io_in[8] & io_in[9] & io_in[10]) | (io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & ~io_in[8] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[2] & io_in[3] & io_in[4] & io_in[6] & ~io_in[7] & io_in[9] & io_in[11]) | (~io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & io_in[5] & io_in[9] & io_in[11]) | (io_in[0] & io_in[1] & io_in[5] & ~io_in[6] & io_in[7] & ~io_in[10]) | (~io_in[0] & io_in[1] & io_in[2] & io_in[4] & ~io_in[6] & ~io_in[7] & ~io_in[8] & ~io_in[9] & io_in[10]) | (~io_in[1] & ~io_in[2] & io_in[4] & ~io_in[6] & ~io_in[7] & io_in[9] & ~io_in[10] & io_in[11]) | (io_in[0] & io_in[2] & ~io_in[4] & ~io_in[6] & io_in[7] & io_in[9] & ~io_in[10] & io_in[11]) | (io_in[0] & io_in[1] & io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[6] & ~io_in[7] & io_in[8] & io_in[9]) | (io_in[0] & ~io_in[2] & io_in[3] & io_in[4] & ~io_in[7] & io_in[8] & io_in[9] & io_in[10] & ~io_in[11]) | (io_in[0] & ~io_in[1] & io_in[2] & ~io_in[4] & ~io_in[6] & io_in[8] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (io_in[1] & ~io_in[2] & io_in[4] & ~io_in[6] & io_in[7] & io_in[8] & ~io_in[9] & io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[3] & io_in[4] & ~io_in[6] & io_in[7] & io_in[8] & ~io_in[9] & io_in[10]) | (~io_in[0] & io_in[1] & ~io_in[2] & io_in[3] & ~io_in[4] & ~io_in[6] & io_in[7] & io_in[8] & ~io_in[11]) | (io_in[0] & io_in[1] & ~io_in[3] & io_in[4] & ~io_in[6] & ~io_in[7] & ~io_in[8] & io_in[9] & io_in[10]) | (io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[6] & io_in[8] & io_in[9] & ~io_in[10]) | (io_in[0] & io_in[1] & ~io_in[2] & ~io_in[4] & ~io_in[5] & io_in[6] & ~io_in[7] & io_in[8] & io_in[11]) | (io_in[0] & io_in[1] & io_in[3] & ~io_in[4] & io_in[6] & io_in[7] & ~io_in[9] & io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & ~io_in[6] & io_in[7] & ~io_in[10] & io_in[11]) | (~io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & io_in[4] & ~io_in[6] & ~io_in[8] & io_in[9] & ~io_in[10] & ~io_in[11]) | (io_in[1] & io_in[2] & ~io_in[3] & io_in[4] & io_in[6] & ~io_in[7] & ~io_in[8] & ~io_in[9] & io_in[11]) | (io_in[0] & io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & ~io_in[7] & ~io_in[8] & ~io_in[9] & ~io_in[11]) | (io_in[0] & io_in[1] & ~io_in[3] & io_in[5] & io_in[6] & ~io_in[9] & io_in[10]) | (io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & io_in[4] & io_in[6] & io_in[7] & ~io_in[9] & io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[3] & io_in[4] & io_in[6] & ~io_in[7] & ~io_in[9] & io_in[11]) | (~io_in[0] & io_in[1] & io_in[2] & ~io_in[3] & io_in[5] & ~io_in[6] & io_in[7] & ~io_in[8] & ~io_in[9]) | (io_in[0] & io_in[1] & io_in[2] & io_in[3] & io_in[4] & io_in[6] & io_in[7] & io_in[8]) | (~io_in[0] & ~io_in[1] & io_in[2] & ~io_in[4] & ~io_in[6] & ~io_in[8] & io_in[9] & io_in[10]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & io_in[5] & ~io_in[6] & ~io_in[7] & io_in[9] & io_in[11]) | (io_in[0] & io_in[1] & io_in[2] & ~io_in[3] & ~io_in[5] & ~io_in[6] & io_in[7] & io_in[10] & io_in[11]) | (~io_in[0] & io_in[1] & io_in[2] & io_in[3] & io_in[4] & io_in[7] & ~io_in[8] & io_in[9] & io_in[10]) | (io_in[1] & ~io_in[2] & io_in[3] & ~io_in[4] & io_in[6] & ~io_in[7] & io_in[8] & ~io_in[9] & ~io_in[11]) | (io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & io_in[5] & ~io_in[6] & ~io_in[8] & ~io_in[9] & io_in[10]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & io_in[3] & io_in[4] & ~io_in[6] & io_in[7] & ~io_in[8] & io_in[9]) | (io_in[0] & ~io_in[2] & io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & io_in[7] & io_in[8] & ~io_in[10]) | (io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[5] & ~io_in[6] & io_in[7] & ~io_in[8] & ~io_in[9] & io_in[11]) | (~io_in[1] & io_in[2] & io_in[5] & ~io_in[7] & ~io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & io_in[4] & ~io_in[6] & io_in[7] & ~io_in[8] & io_in[10]) | (io_in[0] & io_in[1] & ~io_in[2] & io_in[4] & ~io_in[7] & ~io_in[8] & io_in[9] & io_in[11]) | (io_in[0] & io_in[2] & io_in[3] & io_in[4] & ~io_in[7] & io_in[8] & ~io_in[9] & io_in[11]) | (io_in[1] & io_in[3] & io_in[4] & io_in[7] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (io_in[0] & io_in[1] & io_in[2] & io_in[4] & io_in[7] & io_in[8] & io_in[9] & ~io_in[10]) | (~io_in[0] & ~io_in[1] & io_in[2] & io_in[4] & io_in[5] & io_in[7]) | (~io_in[0] & ~io_in[2] & io_in[3] & ~io_in[4] & ~io_in[5] & io_in[7] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (io_in[0] & io_in[1] & io_in[2] & ~io_in[3] & io_in[4] & ~io_in[6] & ~io_in[7] & ~io_in[9] & io_in[10]) | (~io_in[0] & ~io_in[3] & io_in[5] & ~io_in[6] & ~io_in[8] & ~io_in[9] & io_in[11]) | (io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & ~io_in[8] & io_in[9] & ~io_in[10] & ~io_in[11]) | (~io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & ~io_in[6] & ~io_in[8] & io_in[9] & io_in[10]) | (~io_in[0] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[6] & ~io_in[7] & io_in[8] & ~io_in[9] & ~io_in[10] & io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[3] & ~io_in[6] & ~io_in[7] & ~io_in[8] & io_in[9] & ~io_in[10] & io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & io_in[3] & io_in[4] & ~io_in[6] & ~io_in[7] & ~io_in[9] & io_in[10]) | (io_in[0] & ~io_in[1] & ~io_in[2] & io_in[3] & io_in[4] & io_in[7] & io_in[8] & io_in[9] & ~io_in[10]) | (~io_in[0] & io_in[1] & io_in[2] & ~io_in[3] & io_in[6] & ~io_in[7] & io_in[10] & io_in[11]) | (io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & io_in[6] & ~io_in[7] & io_in[8] & ~io_in[10] & io_in[11]) | (io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[6] & io_in[8] & ~io_in[9] & io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[3] & ~io_in[4] & ~io_in[7] & ~io_in[8] & ~io_in[10] & ~io_in[11]) | (io_in[0] & io_in[1] & ~io_in[3] & ~io_in[4] & io_in[6] & ~io_in[7] & ~io_in[9] & io_in[10]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & ~io_in[6] & ~io_in[8] & ~io_in[9] & io_in[11]) | (~io_in[0] & io_in[1] & io_in[3] & ~io_in[4] & ~io_in[6] & io_in[7] & io_in[8] & ~io_in[9] & io_in[10]) | (~io_in[0] & io_in[1] & ~io_in[2] & io_in[4] & ~io_in[6] & ~io_in[7] & io_in[8] & ~io_in[9] & io_in[10]) | (~io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & io_in[4] & ~io_in[6] & ~io_in[7] & io_in[8] & io_in[10]) | (io_in[0] & io_in[1] & ~io_in[2] & io_in[3] & ~io_in[4] & ~io_in[6] & ~io_in[8] & ~io_in[9] & io_in[10]) | (~io_in[0] & ~io_in[1] & ~io_in[3] & ~io_in[4] & io_in[7] & io_in[8] & io_in[9] & io_in[10] & io_in[11]) | (~io_in[0] & ~io_in[1] & io_in[4] & io_in[6] & ~io_in[7] & ~io_in[8] & ~io_in[9] & io_in[11]) | (io_in[0] & ~io_in[2] & ~io_in[3] & io_in[4] & ~io_in[6] & io_in[7] & ~io_in[8] & io_in[9] & io_in[10]) | (io_in[1] & ~io_in[2] & ~io_in[5] & io_in[6] & io_in[7] & ~io_in[8] & ~io_in[9] & io_in[11]) | (~io_in[0] & io_in[1] & io_in[2] & io_in[3] & io_in[4] & io_in[6] & ~io_in[8] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[1] & io_in[3] & io_in[4] & io_in[6] & io_in[7] & io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[6] & ~io_in[7] & ~io_in[8]) | (~io_in[0] & io_in[1] & ~io_in[3] & ~io_in[5] & ~io_in[6] & ~io_in[7] & io_in[8] & io_in[9] & io_in[10] & ~io_in[11]) | (io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[5] & ~io_in[6] & io_in[7] & ~io_in[8] & io_in[9] & io_in[10]) | (io_in[0] & io_in[1] & io_in[2] & io_in[3] & io_in[4] & io_in[8] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[1] & io_in[2] & ~io_in[4] & ~io_in[5] & ~io_in[6] & ~io_in[7] & io_in[8] & ~io_in[9] & io_in[10]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & io_in[4] & io_in[6] & io_in[7] & io_in[9] & io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[7] & ~io_in[8] & io_in[9] & io_in[10]) | (io_in[0] & ~io_in[2] & io_in[5] & ~io_in[7] & ~io_in[8] & io_in[9] & io_in[10]) | (io_in[0] & ~io_in[2] & ~io_in[3] & ~io_in[5] & io_in[6] & io_in[7] & ~io_in[8] & ~io_in[9] & io_in[10]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & io_in[4] & io_in[6] & ~io_in[7] & ~io_in[8] & ~io_in[9] & ~io_in[10]) | (~io_in[1] & ~io_in[3] & ~io_in[4] & io_in[6] & io_in[7] & ~io_in[8] & io_in[9] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & ~io_in[2] & ~io_in[3] & io_in[4] & ~io_in[6] & io_in[7] & io_in[8] & io_in[9] & ~io_in[10]) | (io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & io_in[6] & io_in[8] & io_in[9] & io_in[10] & ~io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & io_in[3] & ~io_in[5] & io_in[6] & ~io_in[7] & ~io_in[8] & ~io_in[9] & io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[5] & io_in[6] & ~io_in[8] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[1] & io_in[2] & io_in[3] & io_in[4] & io_in[6] & ~io_in[7] & io_in[8] & io_in[10]) | (io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[5] & io_in[6] & ~io_in[7] & io_in[8] & io_in[10] & ~io_in[11]) | (~io_in[1] & io_in[2] & io_in[3] & io_in[4] & io_in[6] & io_in[7] & io_in[8] & io_in[9] & ~io_in[10]) | (io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & ~io_in[6] & io_in[7] & io_in[10] & io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[4] & io_in[7] & io_in[8] & io_in[9] & io_in[10] & io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & io_in[4] & io_in[5] & ~io_in[6] & ~io_in[7]) | (io_in[0] & io_in[1] & ~io_in[3] & io_in[5] & io_in[6] & ~io_in[7] & io_in[10] & io_in[11]) | (~io_in[1] & io_in[2] & ~io_in[3] & io_in[5] & io_in[6] & io_in[8] & ~io_in[10]) | (~io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & ~io_in[5] & io_in[7] & ~io_in[8] & io_in[9] & io_in[10]) | (io_in[0] & ~io_in[1] & ~io_in[2] & io_in[3] & io_in[4] & ~io_in[7] & ~io_in[8] & io_in[11]) | (io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & ~io_in[6] & io_in[8] & io_in[9] & ~io_in[10]) | (io_in[0] & ~io_in[1] & ~io_in[3] & ~io_in[5] & io_in[6] & io_in[7] & io_in[8] & io_in[9] & ~io_in[10]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & ~io_in[6] & ~io_in[7] & ~io_in[9] & ~io_in[11]) | (io_in[0] & io_in[3] & io_in[5] & ~io_in[7] & ~io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[4] & ~io_in[6] & io_in[7] & ~io_in[8] & ~io_in[9] & ~io_in[10] & io_in[11]) | (io_in[0] & ~io_in[2] & ~io_in[3] & io_in[4] & io_in[6] & io_in[7] & io_in[9] & ~io_in[10] & ~io_in[11]) | (io_in[0] & io_in[1] & io_in[2] & io_in[5] & ~io_in[6] & io_in[9] & ~io_in[11]) | (~io_in[0] & io_in[2] & ~io_in[3] & io_in[4] & io_in[6] & ~io_in[7] & ~io_in[8] & io_in[9] & io_in[10]) | (io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & io_in[4] & io_in[6] & io_in[7] & io_in[10] & ~io_in[11]) | (io_in[0] & io_in[1] & io_in[3] & io_in[4] & ~io_in[6] & ~io_in[8] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & ~io_in[8] & ~io_in[9] & io_in[10]) | (~io_in[0] & io_in[1] & ~io_in[2] & io_in[3] & ~io_in[5] & ~io_in[6] & ~io_in[7] & io_in[8] & io_in[11]) | (io_in[1] & io_in[2] & io_in[3] & ~io_in[6] & io_in[7] & io_in[8] & io_in[9] & ~io_in[10]) | (io_in[0] & ~io_in[2] & ~io_in[3] & ~io_in[4] & io_in[6] & io_in[9] & ~io_in[10] & io_in[11]) | (io_in[0] & ~io_in[1] & ~io_in[2] & io_in[3] & io_in[4] & ~io_in[7] & io_in[9] & io_in[11]) | (io_in[0] & ~io_in[1] & io_in[5] & io_in[6] & io_in[7] & ~io_in[8] & io_in[11]) | (io_in[0] & io_in[2] & io_in[3] & ~io_in[4] & ~io_in[6] & ~io_in[7] & ~io_in[8] & io_in[9]) | (io_in[1] & ~io_in[2] & ~io_in[3] & io_in[5] & ~io_in[7] & ~io_in[9] & io_in[10]) | (io_in[0] & io_in[1] & io_in[2] & io_in[4] & io_in[6] & io_in[7] & io_in[10] & io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & io_in[3] & io_in[4] & ~io_in[6] & io_in[7] & io_in[8] & ~io_in[9]) | (io_in[0] & io_in[2] & ~io_in[4] & io_in[6] & io_in[7] & io_in[8] & ~io_in[9] & io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & io_in[4] & ~io_in[6] & io_in[7] & ~io_in[8] & io_in[9] & io_in[10]) | (io_in[0] & ~io_in[1] & io_in[3] & io_in[5] & io_in[6] & io_in[7] & ~io_in[9]) | (~io_in[0] & io_in[2] & io_in[4] & io_in[6] & io_in[7] & io_in[9] & ~io_in[10] & io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & io_in[4] & io_in[5] & io_in[7]) | (io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & io_in[5] & ~io_in[7] & io_in[10] & io_in[11]) | (io_in[0] & ~io_in[2] & io_in[3] & ~io_in[4] & io_in[6] & ~io_in[7] & ~io_in[8] & io_in[9] & io_in[10]) | (~io_in[0] & io_in[1] & io_in[2] & io_in[5] & io_in[6] & io_in[7] & io_in[8] & io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & io_in[7] & io_in[10] & ~io_in[11]) | (io_in[0] & io_in[1] & io_in[2] & ~io_in[4] & io_in[6] & ~io_in[7] & ~io_in[9] & io_in[10]) | (io_in[0] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[6] & io_in[7] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & ~io_in[6] & io_in[7] & ~io_in[9] & ~io_in[10]) | (io_in[0] & ~io_in[2] & io_in[3] & ~io_in[4] & io_in[6] & io_in[8] & ~io_in[9] & ~io_in[10]) | (~io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & io_in[6] & ~io_in[7] & io_in[9] & io_in[11]) | (io_in[0] & ~io_in[1] & io_in[2] & io_in[5] & ~io_in[7] & ~io_in[9] & io_in[10]) | (~io_in[0] & io_in[1] & ~io_in[3] & ~io_in[4] & ~io_in[6] & ~io_in[8] & io_in[9] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & ~io_in[6] & ~io_in[8] & io_in[9] & ~io_in[11]) | (io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & io_in[4] & ~io_in[6] & ~io_in[7] & ~io_in[8] & io_in[10]) | (~io_in[0] & io_in[1] & io_in[2] & ~io_in[4] & ~io_in[6] & ~io_in[8] & ~io_in[9] & io_in[11]) | (~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[6] & io_in[7] & io_in[8] & ~io_in[9] & io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & io_in[6] & io_in[7] & io_in[8] & io_in[9]) | (io_in[0] & ~io_in[3] & io_in[4] & ~io_in[5] & ~io_in[6] & ~io_in[7] & io_in[10] & io_in[11]) | (io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & ~io_in[6] & io_in[7] & io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & io_in[8] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[4] & ~io_in[5] & io_in[6] & ~io_in[8] & io_in[9] & io_in[10]) | (io_in[1] & ~io_in[2] & io_in[3] & ~io_in[4] & ~io_in[6] & io_in[7] & ~io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & io_in[4] & io_in[7] & io_in[8] & ~io_in[9]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & io_in[5] & ~io_in[6] & io_in[7] & io_in[9] & io_in[10] & ~io_in[11]) | (io_in[1] & ~io_in[2] & io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[7] & io_in[10] & io_in[11]) | (io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[6] & io_in[7] & io_in[8] & io_in[9] & ~io_in[10]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[4] & io_in[6] & ~io_in[7] & io_in[8] & ~io_in[9] & ~io_in[10] & io_in[11]) | (~io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & io_in[4] & ~io_in[6] & io_in[8] & io_in[9]) | (~io_in[0] & io_in[1] & io_in[2] & io_in[3] & io_in[5] & ~io_in[6] & ~io_in[7]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & io_in[5] & ~io_in[7] & io_in[8] & io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[1] & io_in[2] & io_in[4] & ~io_in[6] & ~io_in[7] & ~io_in[8] & io_in[9] & io_in[11]) | (io_in[0] & io_in[1] & io_in[2] & ~io_in[3] & ~io_in[5] & io_in[6] & io_in[7] & ~io_in[8] & io_in[9] & io_in[10]) | (~io_in[0] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & io_in[10] & io_in[11]) | (io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[4] & ~io_in[6] & io_in[7] & io_in[8] & ~io_in[9] & io_in[10]) | (~io_in[2] & io_in[3] & io_in[5] & io_in[7] & io_in[8] & io_in[11]) | (~io_in[0] & io_in[2] & io_in[3] & io_in[4] & io_in[7] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & io_in[3] & ~io_in[4] & ~io_in[6] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[6] & io_in[8] & io_in[9] & io_in[10] & io_in[11]) | (io_in[0] & io_in[2] & io_in[3] & ~io_in[4] & io_in[7] & io_in[9] & ~io_in[10] & io_in[11]) | (io_in[0] & io_in[1] & ~io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[7] & ~io_in[8] & io_in[9] & io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[6] & ~io_in[7] & io_in[8] & io_in[9] & ~io_in[11]) | (~io_in[0] & io_in[2] & io_in[3] & io_in[4] & ~io_in[6] & io_in[7] & ~io_in[8] & io_in[10]) | (io_in[1] & io_in[2] & io_in[3] & io_in[4] & ~io_in[6] & ~io_in[7] & io_in[11]) | (io_in[0] & io_in[1] & io_in[3] & ~io_in[4] & io_in[7] & io_in[8] & ~io_in[10] & io_in[11]) | (~io_in[0] & ~io_in[1] & io_in[3] & io_in[5] & ~io_in[6] & io_in[7] & ~io_in[11]) | (io_in[0] & io_in[1] & io_in[2] & io_in[3] & io_in[6] & io_in[7] & io_in[8] & ~io_in[9]) | (~io_in[0] & io_in[2] & io_in[4] & io_in[5] & io_in[6]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[6] & ~io_in[7] & io_in[8] & ~io_in[9] & io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & io_in[3] & io_in[4] & io_in[6] & io_in[7] & io_in[8] & io_in[10]) | (~io_in[0] & ~io_in[2] & io_in[3] & io_in[5] & io_in[8] & ~io_in[10]) | (io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & ~io_in[7] & ~io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & io_in[1] & io_in[2] & io_in[3] & io_in[4] & io_in[6] & ~io_in[7] & ~io_in[8] & io_in[10]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & io_in[3] & io_in[4] & io_in[6] & ~io_in[7] & io_in[8] & io_in[9]) | (io_in[1] & io_in[3] & io_in[5] & io_in[8] & ~io_in[10]) | (io_in[0] & io_in[2] & ~io_in[3] & io_in[4] & ~io_in[5] & ~io_in[6] & io_in[10] & io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[4] & io_in[6] & io_in[7] & ~io_in[8] & io_in[9] & ~io_in[10]) | (~io_in[0] & io_in[1] & ~io_in[4] & ~io_in[6] & ~io_in[7] & ~io_in[8] & ~io_in[9] & io_in[11]) | (~io_in[0] & io_in[1] & io_in[2] & io_in[4] & io_in[6] & io_in[7] & ~io_in[8] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[7] & io_in[8] & ~io_in[9] & io_in[10]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & io_in[7] & io_in[8] & io_in[9] & io_in[10] & ~io_in[11]) | (io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[4] & io_in[6] & ~io_in[7] & ~io_in[8] & io_in[9] & io_in[11]) | (io_in[0] & ~io_in[2] & ~io_in[4] & ~io_in[5] & ~io_in[6] & io_in[7] & io_in[10] & io_in[11]) | (io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & io_in[6] & io_in[7] & io_in[8] & ~io_in[9]) | (~io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & io_in[6] & io_in[8] & ~io_in[9] & ~io_in[11]) | (~io_in[0] & io_in[1] & io_in[2] & ~io_in[3] & io_in[4] & io_in[8] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & io_in[6] & io_in[7] & io_in[9] & io_in[10]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[5] & io_in[6] & ~io_in[7] & io_in[8] & io_in[9] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & io_in[3] & io_in[4] & io_in[7] & io_in[8] & io_in[11]) | (~io_in[0] & ~io_in[2] & io_in[3] & io_in[4] & io_in[7] & ~io_in[9] & io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[4] & ~io_in[6] & io_in[7] & io_in[8] & io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[6] & io_in[7] & io_in[8] & ~io_in[10]) | (~io_in[0] & io_in[1] & ~io_in[2] & io_in[5] & io_in[6] & io_in[7] & io_in[9] & ~io_in[10]) | (~io_in[0] & ~io_in[2] & io_in[3] & io_in[6] & ~io_in[7] & io_in[8] & ~io_in[9] & io_in[10]) | (~io_in[0] & io_in[1] & ~io_in[2] & io_in[4] & io_in[6] & io_in[7] & ~io_in[9] & ~io_in[10]) | (io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[7] & ~io_in[8] & io_in[9]) | (io_in[0] & io_in[1] & ~io_in[2] & io_in[3] & ~io_in[4] & ~io_in[6] & io_in[9] & io_in[11]) | (~io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[6] & ~io_in[7] & io_in[9] & io_in[10] & ~io_in[11]) | (io_in[0] & io_in[1] & io_in[2] & ~io_in[3] & io_in[6] & ~io_in[7] & ~io_in[8] & ~io_in[9] & io_in[11]) | (io_in[0] & ~io_in[2] & io_in[3] & io_in[4] & io_in[6] & ~io_in[7] & ~io_in[8] & ~io_in[9] & io_in[10]) | (~io_in[0] & io_in[1] & io_in[3] & ~io_in[4] & io_in[6] & ~io_in[8] & io_in[9] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & ~io_in[7] & ~io_in[8] & io_in[9] & io_in[10]);

assign val[2] = (~io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (io_in[0] & io_in[1] & io_in[2] & io_in[3] & ~io_in[7] & ~io_in[8] & ~io_in[9] & io_in[10]) | (~io_in[1] & io_in[3] & io_in[4] & io_in[6] & io_in[7] & io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & io_in[6] & ~io_in[7] & ~io_in[8] & io_in[11]) | (~io_in[2] & ~io_in[3] & io_in[4] & io_in[6] & io_in[7] & io_in[8] & ~io_in[10] & io_in[11]) | (~io_in[2] & ~io_in[3] & io_in[4] & ~io_in[6] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (io_in[0] & ~io_in[2] & io_in[3] & ~io_in[4] & ~io_in[6] & io_in[7] & io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[3] & io_in[4] & ~io_in[7] & ~io_in[8] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[7] & io_in[9] & io_in[11]) | (io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & ~io_in[7] & ~io_in[8] & ~io_in[9] & io_in[10]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & io_in[9] & io_in[11]) | (io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & io_in[7] & io_in[8] & ~io_in[9] & io_in[11]) | (io_in[0] & io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[7] & io_in[8] & ~io_in[9] & io_in[11]) | (io_in[0] & io_in[1] & io_in[2] & io_in[3] & io_in[4] & io_in[7] & io_in[8] & ~io_in[9]) | (~io_in[1] & io_in[3] & ~io_in[4] & io_in[6] & ~io_in[7] & ~io_in[8] & io_in[9] & io_in[10]) | (io_in[0] & io_in[1] & io_in[5] & io_in[6] & io_in[7] & ~io_in[8] & io_in[9]) | (~io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & ~io_in[6] & ~io_in[7] & io_in[8] & ~io_in[9] & ~io_in[10]) | (~io_in[0] & ~io_in[1] & io_in[2] & ~io_in[4] & io_in[6] & io_in[7] & io_in[8] & ~io_in[9]) | (io_in[0] & ~io_in[1] & io_in[5] & ~io_in[6] & ~io_in[8] & io_in[9] & io_in[10]) | (io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & ~io_in[6] & ~io_in[8] & io_in[9] & io_in[10]) | (io_in[0] & io_in[1] & io_in[2] & io_in[3] & io_in[4] & io_in[6] & ~io_in[9] & io_in[11]) | (io_in[0] & io_in[2] & io_in[3] & ~io_in[4] & ~io_in[6] & ~io_in[7] & io_in[8] & ~io_in[9] & io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & io_in[4] & ~io_in[5] & ~io_in[6] & ~io_in[7] & io_in[9] & io_in[10]) | (~io_in[0] & io_in[2] & io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[6] & ~io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & ~io_in[1] & ~io_in[2] & io_in[3] & ~io_in[5] & io_in[6] & ~io_in[7] & io_in[10] & io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[5] & io_in[7] & ~io_in[8] & io_in[9] & io_in[10] & ~io_in[11]) | (io_in[1] & ~io_in[2] & io_in[3] & io_in[4] & ~io_in[7] & io_in[8] & io_in[9] & io_in[10] & ~io_in[11]) | (~io_in[1] & io_in[2] & io_in[3] & io_in[4] & ~io_in[6] & ~io_in[7] & ~io_in[8] & io_in[9] & io_in[10]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[5] & ~io_in[6] & ~io_in[7] & ~io_in[8] & io_in[10]) | (~io_in[0] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[6] & ~io_in[7] & io_in[8] & io_in[10]) | (io_in[1] & ~io_in[2] & io_in[4] & ~io_in[6] & io_in[7] & ~io_in[8] & io_in[9] & io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[3] & ~io_in[4] & ~io_in[6] & io_in[7] & io_in[8] & ~io_in[9]) | (io_in[0] & io_in[2] & io_in[3] & io_in[4] & ~io_in[7] & io_in[8] & ~io_in[10] & ~io_in[11]) | (io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & ~io_in[6] & io_in[9] & ~io_in[10] & io_in[11]) | (io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[4] & ~io_in[6] & io_in[7] & io_in[8] & ~io_in[9]) | (io_in[1] & ~io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[6] & io_in[7] & io_in[8] & ~io_in[9] & io_in[10]) | (io_in[1] & ~io_in[3] & io_in[4] & ~io_in[6] & io_in[7] & ~io_in[8] & ~io_in[9] & ~io_in[10]) | (~io_in[0] & io_in[2] & ~io_in[3] & io_in[5] & ~io_in[6] & io_in[7] & ~io_in[9] & io_in[11]) | (io_in[0] & io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & ~io_in[6] & io_in[7] & io_in[8] & io_in[9]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & io_in[3] & io_in[5] & io_in[6] & io_in[8]) | (~io_in[0] & io_in[2] & ~io_in[3] & io_in[4] & ~io_in[7] & ~io_in[8] & ~io_in[9] & io_in[11]) | (io_in[0] & io_in[1] & ~io_in[2] & io_in[3] & io_in[4] & io_in[6] & io_in[7] & io_in[9] & io_in[10] & ~io_in[11]) | (io_in[0] & ~io_in[1] & io_in[2] & io_in[4] & ~io_in[7] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & io_in[7] & ~io_in[9] & io_in[11]) | (~io_in[0] & ~io_in[2] & ~io_in[3] & io_in[4] & ~io_in[5] & io_in[6] & ~io_in[7] & io_in[10] & io_in[11]) | (~io_in[1] & io_in[2] & io_in[3] & io_in[4] & ~io_in[6] & io_in[7] & io_in[9] & io_in[11]) | (~io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & ~io_in[9] & io_in[10] & ~io_in[11]) | (io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & ~io_in[8] & io_in[10]) | (~io_in[0] & ~io_in[1] & io_in[3] & ~io_in[4] & ~io_in[5] & io_in[7] & ~io_in[8] & ~io_in[9] & ~io_in[11]) | (io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[5] & io_in[6] & ~io_in[7] & ~io_in[8] & ~io_in[9] & io_in[10]) | (~io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & ~io_in[6] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & io_in[4] & ~io_in[6] & io_in[7] & io_in[9] & io_in[10]) | (~io_in[0] & ~io_in[1] & ~io_in[3] & ~io_in[4] & ~io_in[6] & ~io_in[7] & ~io_in[8] & io_in[10] & ~io_in[11]) | (~io_in[0] & ~io_in[2] & ~io_in[3] & io_in[4] & ~io_in[6] & ~io_in[8] & io_in[9] & io_in[10]) | (~io_in[0] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[7] & io_in[8] & io_in[9] & io_in[10] & ~io_in[11]) | (io_in[0] & ~io_in[1] & io_in[3] & ~io_in[4] & ~io_in[6] & ~io_in[7] & io_in[8] & io_in[10] & ~io_in[11]) | (io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & ~io_in[6] & io_in[7] & ~io_in[8] & io_in[9] & ~io_in[10]) | (~io_in[0] & io_in[2] & io_in[3] & ~io_in[4] & io_in[6] & ~io_in[7] & io_in[8] & ~io_in[9] & io_in[10]) | (~io_in[0] & io_in[1] & io_in[3] & io_in[4] & ~io_in[6] & ~io_in[7] & io_in[9] & ~io_in[11]) | (io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[6] & io_in[11]) | (~io_in[1] & ~io_in[2] & io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & io_in[7] & io_in[8] & io_in[9] & io_in[10] & ~io_in[11]) | (io_in[0] & io_in[1] & ~io_in[2] & io_in[3] & ~io_in[4] & ~io_in[6] & ~io_in[8] & io_in[9] & io_in[10]) | (~io_in[0] & ~io_in[1] & ~io_in[4] & ~io_in[5] & ~io_in[6] & io_in[7] & io_in[9] & ~io_in[10] & ~io_in[11]) | (io_in[0] & ~io_in[2] & ~io_in[4] & io_in[6] & ~io_in[7] & io_in[8] & ~io_in[9] & io_in[10]) | (io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & io_in[7] & io_in[10] & io_in[11]) | (io_in[0] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & ~io_in[7] & io_in[8] & io_in[9] & ~io_in[10]) | (io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & ~io_in[6] & io_in[7] & io_in[10] & io_in[11]) | (io_in[0] & ~io_in[1] & ~io_in[2] & io_in[4] & io_in[6] & ~io_in[8] & io_in[9] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & io_in[5] & io_in[6] & ~io_in[8] & io_in[9]) | (~io_in[0] & io_in[1] & io_in[2] & io_in[3] & io_in[4] & io_in[8] & ~io_in[9] & ~io_in[10]) | (io_in[1] & io_in[3] & io_in[6] & io_in[8] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (io_in[0] & io_in[1] & ~io_in[2] & io_in[4] & io_in[6] & io_in[8] & io_in[9] & io_in[10] & ~io_in[11]) | (io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & ~io_in[7] & io_in[8] & io_in[9] & ~io_in[10]) | (io_in[0] & io_in[1] & io_in[2] & ~io_in[3] & io_in[6] & io_in[8] & ~io_in[9] & io_in[10]) | (io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[6] & io_in[8] & ~io_in[10] & io_in[11]) | (io_in[0] & ~io_in[1] & io_in[2] & io_in[5] & ~io_in[7] & ~io_in[8] & io_in[11]) | (io_in[0] & io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[7] & io_in[9] & io_in[10]) | (~io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & io_in[4] & ~io_in[6] & io_in[8] & io_in[10] & ~io_in[11]) | (~io_in[1] & io_in[2] & ~io_in[3] & io_in[4] & io_in[6] & ~io_in[7] & ~io_in[8] & io_in[9] & io_in[10]) | (io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & io_in[4] & ~io_in[6] & ~io_in[7] & ~io_in[11]) | (~io_in[1] & ~io_in[2] & io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[6] & ~io_in[7] & io_in[8] & io_in[10] & ~io_in[11]) | (~io_in[1] & io_in[2] & ~io_in[3] & io_in[4] & io_in[7] & ~io_in[9] & io_in[10]) | (~io_in[1] & io_in[2] & io_in[3] & io_in[4] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (io_in[2] & ~io_in[3] & io_in[5] & io_in[6] & io_in[7] & ~io_in[8] & io_in[9]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & io_in[3] & ~io_in[4] & ~io_in[8] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[2] & ~io_in[3] & io_in[4] & ~io_in[6] & io_in[7] & io_in[8] & io_in[9] & ~io_in[11]) | (io_in[0] & ~io_in[1] & io_in[5] & ~io_in[7] & io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[6] & io_in[7] & ~io_in[9] & io_in[10]) | (io_in[0] & io_in[1] & io_in[5] & ~io_in[6] & io_in[8] & io_in[9] & ~io_in[11]) | (io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[4] & ~io_in[7] & ~io_in[8] & io_in[9] & io_in[10]) | (~io_in[0] & io_in[1] & ~io_in[2] & io_in[3] & ~io_in[4] & io_in[8] & ~io_in[10] & ~io_in[11]) | (io_in[0] & io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[6] & io_in[8] & io_in[9] & io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[1] & io_in[2] & io_in[3] & ~io_in[6] & ~io_in[7] & ~io_in[8] & ~io_in[9]) | (io_in[1] & io_in[2] & io_in[3] & io_in[5] & ~io_in[6] & ~io_in[7]) | (io_in[0] & io_in[1] & io_in[2] & ~io_in[4] & io_in[6] & ~io_in[7] & ~io_in[8] & ~io_in[9] & ~io_in[11]) | (~io_in[0] & io_in[3] & ~io_in[4] & ~io_in[6] & io_in[7] & ~io_in[8] & io_in[9] & ~io_in[10]) | (~io_in[0] & ~io_in[1] & ~io_in[3] & ~io_in[4] & ~io_in[6] & ~io_in[7] & ~io_in[9] & ~io_in[10] & io_in[11]) | (~io_in[0] & io_in[1] & io_in[2] & io_in[3] & ~io_in[6] & io_in[7] & io_in[9] & io_in[10] & ~io_in[11]) | (~io_in[0] & ~io_in[1] & io_in[3] & io_in[4] & io_in[6] & io_in[7] & io_in[8] & ~io_in[11]) | (~io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & ~io_in[7] & io_in[10] & io_in[11]) | (io_in[0] & ~io_in[1] & ~io_in[2] & io_in[3] & io_in[4] & ~io_in[6] & ~io_in[7] & io_in[9] & io_in[11]) | (io_in[0] & io_in[2] & ~io_in[3] & io_in[4] & ~io_in[6] & io_in[7] & ~io_in[8] & ~io_in[9] & io_in[11]) | (io_in[0] & io_in[1] & io_in[2] & io_in[5] & io_in[6] & ~io_in[8] & ~io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[6] & ~io_in[9] & io_in[10]) | (io_in[1] & ~io_in[2] & io_in[3] & io_in[5] & io_in[7] & io_in[10] & io_in[11]) | (io_in[1] & ~io_in[2] & ~io_in[4] & ~io_in[5] & io_in[6] & io_in[8] & io_in[9] & ~io_in[10]) | (~io_in[1] & io_in[2] & io_in[3] & io_in[4] & io_in[6] & ~io_in[8] & io_in[9] & io_in[11]) | (io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & ~io_in[7] & ~io_in[8] & ~io_in[9]) | (~io_in[0] & io_in[1] & io_in[5] & io_in[6] & ~io_in[7] & ~io_in[11]) | (~io_in[0] & ~io_in[1] & io_in[2] & io_in[4] & io_in[6] & io_in[7] & io_in[9] & io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & io_in[6] & ~io_in[7] & io_in[10]) | (~io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & ~io_in[5] & io_in[7] & ~io_in[9] & ~io_in[10]) | (io_in[0] & ~io_in[1] & ~io_in[2] & io_in[3] & io_in[4] & ~io_in[6] & ~io_in[7] & io_in[8] & io_in[9]) | (~io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & io_in[6] & ~io_in[7] & io_in[8] & ~io_in[9] & ~io_in[10]) | (io_in[0] & io_in[2] & io_in[5] & ~io_in[6] & io_in[9] & ~io_in[11]) | (~io_in[0] & io_in[2] & ~io_in[3] & io_in[4] & ~io_in[6] & ~io_in[7] & ~io_in[8] & io_in[11]) | (io_in[0] & io_in[5] & ~io_in[6] & io_in[7] & io_in[9] & ~io_in[10]) | (~io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & io_in[7] & io_in[8] & ~io_in[9] & io_in[10]) | (io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & io_in[6] & ~io_in[7] & ~io_in[8] & ~io_in[9] & io_in[11]) | (io_in[0] & ~io_in[1] & io_in[2] & ~io_in[6] & ~io_in[7] & io_in[8] & io_in[9] & ~io_in[10]) | (~io_in[0] & ~io_in[1] & io_in[2] & io_in[4] & io_in[7] & ~io_in[9] & io_in[10]) | (io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & io_in[8] & ~io_in[10]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & io_in[3] & ~io_in[4] & io_in[6] & io_in[8] & ~io_in[10] & io_in[11]) | (io_in[1] & ~io_in[3] & io_in[4] & ~io_in[5] & io_in[6] & ~io_in[7] & io_in[10] & io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[3] & io_in[5] & io_in[6] & ~io_in[7] & io_in[8] & io_in[10]) | (~io_in[0] & ~io_in[1] & io_in[5] & ~io_in[6] & ~io_in[7] & ~io_in[8] & io_in[10]) | (io_in[0] & ~io_in[2] & io_in[3] & ~io_in[4] & io_in[6] & ~io_in[7] & ~io_in[8] & io_in[9]) | (io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & io_in[5] & io_in[8] & ~io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[3] & ~io_in[4] & io_in[5] & ~io_in[6] & io_in[7] & io_in[9] & io_in[11]) | (io_in[1] & ~io_in[3] & io_in[4] & ~io_in[6] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (~io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & ~io_in[6] & io_in[8] & ~io_in[9] & io_in[11]) | (io_in[0] & io_in[1] & io_in[3] & ~io_in[4] & ~io_in[6] & ~io_in[7] & ~io_in[8] & io_in[9]) | (~io_in[1] & ~io_in[2] & io_in[3] & ~io_in[4] & ~io_in[6] & ~io_in[8] & ~io_in[10] & ~io_in[11]) | (io_in[0] & io_in[1] & io_in[2] & ~io_in[4] & io_in[6] & io_in[7] & ~io_in[8] & io_in[9] & io_in[10]) | (io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[6] & io_in[7] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[2] & io_in[3] & io_in[4] & ~io_in[7] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (~io_in[2] & ~io_in[3] & io_in[4] & ~io_in[6] & io_in[7] & ~io_in[8] & io_in[9] & io_in[11]) | (io_in[0] & ~io_in[2] & io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & io_in[7] & ~io_in[8] & ~io_in[9] & io_in[10]) | (~io_in[0] & io_in[1] & io_in[2] & io_in[6] & io_in[8] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & io_in[6] & ~io_in[7] & io_in[8] & io_in[9] & io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[4] & ~io_in[5] & io_in[6] & io_in[7] & io_in[9] & io_in[10]) | (~io_in[0] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & ~io_in[8] & io_in[9] & ~io_in[11]) | (io_in[0] & ~io_in[1] & io_in[2] & io_in[4] & ~io_in[6] & io_in[8] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & ~io_in[2] & ~io_in[3] & io_in[4] & io_in[6] & io_in[7] & io_in[8] & ~io_in[10]) | (io_in[0] & io_in[1] & io_in[2] & ~io_in[4] & ~io_in[5] & ~io_in[6] & ~io_in[7] & io_in[9] & ~io_in[10] & io_in[11]) | (io_in[0] & ~io_in[2] & io_in[3] & ~io_in[4] & io_in[6] & ~io_in[7] & io_in[8] & ~io_in[9] & ~io_in[11]) | (io_in[0] & io_in[1] & ~io_in[2] & ~io_in[4] & ~io_in[5] & io_in[7] & ~io_in[8] & ~io_in[9] & io_in[11]) | (io_in[0] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & ~io_in[7] & io_in[9] & ~io_in[11]) | (io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[10] & io_in[11]) | (~io_in[0] & io_in[3] & io_in[4] & io_in[6] & io_in[7] & io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & io_in[1] & ~io_in[2] & io_in[3] & ~io_in[4] & io_in[7] & io_in[11]) | (io_in[1] & io_in[2] & ~io_in[3] & io_in[4] & io_in[6] & ~io_in[7] & ~io_in[8] & ~io_in[10]) | (io_in[0] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[6] & io_in[7] & io_in[8] & io_in[10]) | (io_in[0] & io_in[1] & io_in[2] & io_in[3] & io_in[5] & io_in[11]) | (io_in[0] & ~io_in[2] & io_in[3] & ~io_in[4] & ~io_in[7] & io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & io_in[1] & io_in[2] & io_in[5] & ~io_in[7] & ~io_in[9]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[4] & ~io_in[5] & io_in[6] & io_in[8] & io_in[9]) | (~io_in[1] & io_in[2] & io_in[6] & io_in[7] & io_in[8] & ~io_in[9] & io_in[10]) | (io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[6] & ~io_in[7] & io_in[10] & io_in[11]) | (~io_in[0] & io_in[2] & io_in[3] & io_in[4] & io_in[6] & ~io_in[7] & io_in[8] & io_in[9] & io_in[10]) | (io_in[0] & io_in[2] & ~io_in[3] & io_in[4] & ~io_in[6] & ~io_in[7] & io_in[8] & ~io_in[9] & ~io_in[10]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[5] & ~io_in[6] & io_in[7] & ~io_in[9] & ~io_in[10]) | (io_in[0] & io_in[1] & io_in[3] & io_in[4] & ~io_in[6] & io_in[7] & io_in[8] & ~io_in[9] & io_in[11]) | (~io_in[0] & io_in[1] & io_in[3] & io_in[4] & io_in[6] & ~io_in[7] & io_in[8] & ~io_in[10] & io_in[11]) | (io_in[0] & ~io_in[2] & io_in[3] & ~io_in[4] & io_in[6] & io_in[7] & io_in[8] & ~io_in[10]) | (io_in[0] & io_in[1] & ~io_in[2] & ~io_in[4] & ~io_in[5] & io_in[6] & ~io_in[8] & ~io_in[9] & io_in[11]) | (~io_in[0] & ~io_in[1] & io_in[2] & ~io_in[4] & ~io_in[5] & io_in[7] & io_in[9] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[2] & ~io_in[4] & ~io_in[5] & ~io_in[6] & ~io_in[7] & io_in[10] & io_in[11]) | (~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[6] & io_in[7] & ~io_in[8] & ~io_in[9] & io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[5] & io_in[6] & io_in[10] & io_in[11]) | (io_in[0] & io_in[1] & io_in[2] & io_in[3] & ~io_in[6] & ~io_in[7] & ~io_in[8] & io_in[9] & io_in[11]) | (~io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & io_in[4] & ~io_in[6] & io_in[9] & ~io_in[10] & ~io_in[11]) | (io_in[1] & io_in[2] & io_in[3] & io_in[4] & io_in[6] & io_in[7] & ~io_in[10] & io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & ~io_in[7] & io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & io_in[3] & ~io_in[6] & ~io_in[7] & ~io_in[8] & io_in[11]) | (io_in[0] & io_in[1] & ~io_in[3] & io_in[4] & io_in[7] & io_in[8] & io_in[9] & io_in[10] & ~io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[4] & ~io_in[5] & io_in[6] & io_in[7] & ~io_in[8] & ~io_in[9] & ~io_in[10] & io_in[11]) | (io_in[0] & io_in[1] & ~io_in[3] & ~io_in[4] & ~io_in[6] & ~io_in[8] & io_in[9] & ~io_in[10] & ~io_in[11]) | (io_in[0] & ~io_in[1] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[7] & io_in[9] & io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[6] & ~io_in[7] & io_in[9] & io_in[10] & ~io_in[11]) | (~io_in[1] & ~io_in[3] & io_in[4] & ~io_in[6] & io_in[7] & io_in[8] & io_in[9] & ~io_in[10]) | (io_in[0] & ~io_in[1] & ~io_in[2] & io_in[3] & io_in[5] & ~io_in[6] & io_in[9]) | (~io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[7] & io_in[9] & io_in[10] & ~io_in[11]) | (io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[6] & io_in[7] & io_in[9] & io_in[11]) | (io_in[0] & io_in[1] & io_in[4] & io_in[5] & io_in[6]) | (io_in[1] & io_in[2] & io_in[5] & ~io_in[8] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[2] & io_in[3] & ~io_in[6] & io_in[7] & io_in[8] & ~io_in[9] & io_in[11]) | (io_in[0] & io_in[1] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & io_in[7] & ~io_in[8] & ~io_in[9] & ~io_in[10]) | (io_in[0] & io_in[1] & ~io_in[2] & io_in[3] & io_in[4] & io_in[6] & ~io_in[7] & io_in[8] & io_in[10]) | (~io_in[0] & ~io_in[1] & io_in[2] & io_in[4] & io_in[6] & io_in[7] & io_in[8] & io_in[10]) | (io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & io_in[6] & io_in[7] & ~io_in[9] & io_in[11]) | (~io_in[0] & io_in[2] & io_in[3] & ~io_in[4] & io_in[6] & ~io_in[7] & ~io_in[8] & ~io_in[9] & io_in[11]) | (~io_in[0] & ~io_in[2] & ~io_in[3] & io_in[4] & io_in[5] & ~io_in[6]) | (io_in[2] & io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[6] & io_in[7] & ~io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & io_in[1] & ~io_in[2] & io_in[3] & io_in[6] & io_in[7] & io_in[8] & io_in[9] & ~io_in[10]) | (~io_in[1] & io_in[3] & io_in[4] & io_in[5]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & io_in[5] & io_in[6] & io_in[9] & io_in[11]) | (~io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & io_in[4] & io_in[8] & ~io_in[9] & io_in[10]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[4] & io_in[6] & ~io_in[7] & ~io_in[8] & ~io_in[9] & io_in[10]) | (~io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[7] & ~io_in[8] & io_in[9]) | (io_in[0] & ~io_in[1] & io_in[2] & io_in[5] & ~io_in[7] & io_in[8] & ~io_in[11]) | (~io_in[1] & ~io_in[3] & io_in[4] & ~io_in[6] & io_in[7] & io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & io_in[2] & ~io_in[3] & io_in[4] & io_in[6] & io_in[7] & io_in[8] & io_in[9] & ~io_in[10]) | (~io_in[1] & ~io_in[2] & io_in[3] & io_in[5] & ~io_in[10]) | (~io_in[0] & io_in[1] & ~io_in[3] & io_in[5] & ~io_in[6] & ~io_in[7] & io_in[10] & io_in[11]) | (io_in[0] & io_in[1] & ~io_in[2] & io_in[3] & io_in[5] & io_in[7] & io_in[9]) | (io_in[1] & io_in[2] & io_in[3] & io_in[4] & ~io_in[7] & io_in[8] & ~io_in[10] & ~io_in[11]) | (io_in[0] & ~io_in[1] & io_in[5] & io_in[6] & ~io_in[7] & io_in[9] & ~io_in[10]) | (io_in[0] & io_in[1] & io_in[2] & ~io_in[4] & io_in[6] & ~io_in[8] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & io_in[7] & ~io_in[8] & io_in[10]) | (io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[6] & io_in[7] & io_in[8] & io_in[9] & ~io_in[10]) | (~io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & io_in[6] & ~io_in[7] & io_in[9] & ~io_in[10]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[7] & ~io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & io_in[2] & ~io_in[3] & io_in[4] & ~io_in[6] & ~io_in[8] & ~io_in[9] & io_in[10]) | (io_in[1] & io_in[2] & ~io_in[3] & io_in[4] & io_in[6] & io_in[7] & io_in[8] & io_in[9] & ~io_in[10]) | (io_in[0] & io_in[3] & ~io_in[4] & ~io_in[6] & io_in[7] & ~io_in[8] & ~io_in[9] & io_in[11]) | (~io_in[1] & ~io_in[3] & ~io_in[4] & io_in[5] & io_in[6] & ~io_in[7] & io_in[9] & io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[10] & io_in[11]) | (io_in[0] & io_in[1] & ~io_in[2] & io_in[3] & ~io_in[7] & ~io_in[8] & ~io_in[10] & ~io_in[11]) | (io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & ~io_in[6] & ~io_in[9] & io_in[11]) | (io_in[0] & io_in[1] & ~io_in[2] & io_in[5] & ~io_in[6] & ~io_in[8] & io_in[11]) | (io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & io_in[8] & io_in[9] & ~io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & ~io_in[7] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[4] & ~io_in[5] & ~io_in[6] & ~io_in[7] & io_in[8] & io_in[11]) | (~io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & io_in[4] & io_in[6] & ~io_in[7] & io_in[10]) | (~io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & ~io_in[8] & io_in[9] & io_in[10]) | (io_in[0] & io_in[1] & io_in[5] & io_in[6] & io_in[7] & io_in[8] & io_in[11]) | (io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[7] & ~io_in[8] & io_in[11]) | (~io_in[2] & io_in[3] & ~io_in[6] & io_in[7] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (io_in[1] & io_in[2] & io_in[4] & ~io_in[6] & ~io_in[7] & ~io_in[8] & ~io_in[9]) | (~io_in[0] & ~io_in[1] & io_in[2] & io_in[5] & io_in[6] & io_in[7] & ~io_in[8] & io_in[10]) | (io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & ~io_in[7] & ~io_in[8] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & ~io_in[1] & io_in[3] & io_in[7] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & ~io_in[6] & ~io_in[7] & io_in[8]) | (~io_in[0] & io_in[1] & io_in[2] & ~io_in[4] & ~io_in[5] & io_in[7] & ~io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & io_in[1] & io_in[3] & io_in[4] & io_in[6] & io_in[7] & ~io_in[8] & ~io_in[9] & ~io_in[10]) | (~io_in[1] & ~io_in[2] & io_in[5] & io_in[7] & ~io_in[8] & ~io_in[10] & ~io_in[11]) | (io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & io_in[7] & io_in[9] & ~io_in[10] & io_in[11]) | (io_in[0] & io_in[1] & io_in[2] & io_in[3] & io_in[4] & io_in[6] & ~io_in[7] & ~io_in[8] & io_in[10]) | (io_in[0] & io_in[1] & ~io_in[2] & ~io_in[4] & io_in[8] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & io_in[3] & io_in[4] & io_in[6] & ~io_in[8] & io_in[9] & ~io_in[10]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & ~io_in[6] & ~io_in[8] & ~io_in[9]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & io_in[6] & io_in[8] & io_in[9] & io_in[10]) | (~io_in[1] & ~io_in[2] & io_in[4] & io_in[8] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & io_in[6] & io_in[7] & ~io_in[8] & ~io_in[9]) | (io_in[0] & io_in[1] & ~io_in[2] & io_in[5] & ~io_in[6] & ~io_in[8] & ~io_in[9]) | (io_in[1] & io_in[3] & ~io_in[4] & io_in[6] & io_in[7] & io_in[8] & ~io_in[10]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & io_in[5] & ~io_in[7] & ~io_in[8] & io_in[9]) | (~io_in[0] & io_in[2] & ~io_in[3] & io_in[4] & io_in[6] & io_in[7] & ~io_in[8] & ~io_in[9] & ~io_in[11]) | (io_in[1] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & io_in[7] & ~io_in[8] & ~io_in[9] & io_in[11]) | (~io_in[0] & ~io_in[1] & io_in[3] & io_in[6] & ~io_in[7] & io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & io_in[5] & io_in[7] & ~io_in[8] & io_in[10]) | (io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[5] & ~io_in[6] & ~io_in[7] & io_in[8] & io_in[11]) | (io_in[0] & io_in[1] & io_in[2] & ~io_in[4] & ~io_in[5] & ~io_in[6] & io_in[7] & io_in[8] & io_in[10]) | (~io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & io_in[7] & io_in[9] & ~io_in[10]) | (io_in[0] & io_in[1] & ~io_in[2] & ~io_in[4] & ~io_in[5] & io_in[6] & io_in[7] & ~io_in[8] & io_in[11]) | (~io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & ~io_in[5] & io_in[6] & io_in[10] & io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & io_in[3] & ~io_in[4] & ~io_in[6] & io_in[7] & ~io_in[8] & io_in[9]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[4] & ~io_in[6] & io_in[7] & io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & io_in[1] & ~io_in[2] & io_in[5] & io_in[7] & io_in[8] & ~io_in[10]) | (~io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & io_in[5] & ~io_in[9] & io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & io_in[5] & io_in[6] & ~io_in[7] & io_in[10]) | (~io_in[1] & io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[7] & io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & ~io_in[2] & ~io_in[3] & ~io_in[5] & io_in[6] & ~io_in[7] & io_in[8] & io_in[9] & ~io_in[10]) | (io_in[0] & ~io_in[1] & ~io_in[2] & io_in[4] & io_in[6] & ~io_in[7] & ~io_in[8] & ~io_in[9] & io_in[11]) | (io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[5] & ~io_in[6] & io_in[8] & ~io_in[9] & ~io_in[10]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & io_in[7] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (io_in[0] & io_in[2] & ~io_in[3] & ~io_in[5] & io_in[6] & io_in[7] & io_in[10] & io_in[11]) | (io_in[2] & io_in[4] & io_in[5] & ~io_in[6] & ~io_in[7]);

assign val[3] = (~io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & io_in[6] & io_in[8] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & io_in[6] & ~io_in[7] & ~io_in[8] & io_in[9]) | (io_in[0] & io_in[1] & io_in[2] & io_in[5] & io_in[6] & ~io_in[8] & io_in[10]) | (io_in[0] & io_in[1] & ~io_in[3] & io_in[4] & ~io_in[6] & ~io_in[7] & ~io_in[8] & io_in[9] & io_in[11]) | (io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & io_in[4] & ~io_in[6] & io_in[8] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[1] & io_in[2] & io_in[4] & io_in[6] & io_in[7] & ~io_in[10] & io_in[11]) | (io_in[0] & io_in[1] & io_in[2] & io_in[3] & io_in[4] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (io_in[0] & io_in[1] & io_in[3] & ~io_in[4] & ~io_in[6] & ~io_in[7] & io_in[8] & ~io_in[10] & io_in[11]) | (~io_in[1] & ~io_in[2] & io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & ~io_in[7] & io_in[10] & io_in[11]) | (io_in[0] & io_in[1] & ~io_in[2] & ~io_in[4] & io_in[6] & io_in[8] & ~io_in[9] & io_in[10]) | (~io_in[1] & ~io_in[2] & io_in[3] & io_in[4] & ~io_in[6] & ~io_in[7] & io_in[10] & io_in[11]) | (io_in[0] & io_in[1] & ~io_in[2] & io_in[4] & io_in[6] & ~io_in[7] & io_in[8] & io_in[9] & ~io_in[10]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & io_in[7] & io_in[8] & ~io_in[9] & io_in[10]) | (~io_in[0] & io_in[1] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & io_in[7] & ~io_in[8] & io_in[9] & io_in[10]) | (io_in[0] & io_in[2] & ~io_in[3] & io_in[4] & ~io_in[7] & ~io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & ~io_in[1] & io_in[2] & io_in[5] & ~io_in[6] & io_in[7] & ~io_in[9] & io_in[10]) | (io_in[0] & ~io_in[1] & ~io_in[2] & io_in[3] & io_in[4] & ~io_in[7] & io_in[10] & io_in[11]) | (~io_in[0] & ~io_in[2] & ~io_in[3] & ~io_in[5] & ~io_in[6] & io_in[7] & ~io_in[8] & io_in[9] & ~io_in[10] & io_in[11]) | (io_in[0] & io_in[1] & ~io_in[3] & ~io_in[4] & io_in[6] & io_in[8] & ~io_in[9] & io_in[10]) | (~io_in[0] & io_in[2] & io_in[3] & io_in[4] & ~io_in[6] & ~io_in[7] & io_in[9] & ~io_in[10]) | (~io_in[0] & ~io_in[2] & io_in[3] & ~io_in[4] & ~io_in[6] & ~io_in[7] & ~io_in[8] & io_in[9] & io_in[11]) | (io_in[0] & ~io_in[2] & io_in[3] & io_in[4] & io_in[7] & ~io_in[8] & io_in[9] & io_in[10]) | (~io_in[0] & ~io_in[2] & io_in[3] & io_in[4] & io_in[6] & ~io_in[7] & ~io_in[8] & ~io_in[9] & io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & io_in[5] & ~io_in[6] & ~io_in[7] & io_in[9] & ~io_in[10]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & io_in[3] & io_in[4] & ~io_in[7] & io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & io_in[1] & ~io_in[4] & ~io_in[7] & ~io_in[8] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[2] & io_in[3] & io_in[4] & io_in[6] & io_in[7] & ~io_in[10] & io_in[11]) | (io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & io_in[6] & io_in[9] & ~io_in[10] & io_in[11]) | (~io_in[0] & io_in[1] & io_in[5] & io_in[6] & io_in[8] & io_in[9] & ~io_in[10]) | (io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & io_in[6] & ~io_in[7] & io_in[8] & io_in[10]) | (~io_in[0] & ~io_in[1] & io_in[2] & ~io_in[4] & ~io_in[5] & io_in[6] & io_in[7] & ~io_in[8] & ~io_in[9] & io_in[11]) | (~io_in[0] & io_in[1] & io_in[4] & io_in[5] & io_in[6]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[8] & ~io_in[10] & io_in[11]) | (io_in[0] & io_in[5] & io_in[7] & io_in[9] & ~io_in[10] & io_in[11]) | (~io_in[0] & ~io_in[1] & io_in[2] & io_in[6] & io_in[7] & io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & ~io_in[1] & io_in[3] & ~io_in[6] & ~io_in[7] & io_in[8] & io_in[9] & ~io_in[10]) | (io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & io_in[4] & ~io_in[5] & io_in[7] & io_in[10] & io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & io_in[7] & ~io_in[9] & ~io_in[10] & io_in[11]) | (~io_in[0] & ~io_in[2] & io_in[3] & io_in[5] & io_in[7] & ~io_in[8] & ~io_in[10]) | (~io_in[0] & io_in[1] & io_in[2] & ~io_in[5] & io_in[6] & ~io_in[7] & io_in[10] & io_in[11]) | (io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[8] & ~io_in[9] & io_in[11]) | (~io_in[0] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[7] & io_in[8] & io_in[9] & io_in[10] & ~io_in[11]) | (~io_in[1] & ~io_in[2] & io_in[3] & ~io_in[4] & ~io_in[6] & io_in[7] & io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[6] & ~io_in[7] & ~io_in[8] & ~io_in[9]) | (~io_in[0] & io_in[1] & ~io_in[3] & io_in[4] & ~io_in[6] & io_in[7] & ~io_in[8] & io_in[9]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & ~io_in[5] & ~io_in[6] & io_in[9] & io_in[11]) | (~io_in[0] & ~io_in[1] & io_in[2] & io_in[4] & ~io_in[6] & io_in[7] & io_in[8] & io_in[9] & ~io_in[10]) | (io_in[0] & io_in[1] & ~io_in[2] & io_in[3] & io_in[4] & ~io_in[7] & io_in[8] & io_in[9] & io_in[10] & ~io_in[11]) | (io_in[0] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[6] & ~io_in[8] & ~io_in[9] & io_in[11]) | (~io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[6] & io_in[7] & io_in[9] & io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & io_in[7] & io_in[8] & io_in[9] & ~io_in[10]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & ~io_in[7] & io_in[9] & ~io_in[10]) | (~io_in[1] & io_in[2] & io_in[3] & io_in[5] & ~io_in[8] & io_in[9]) | (io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & ~io_in[6] & io_in[7] & io_in[8] & io_in[9] & ~io_in[11]) | (io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & ~io_in[6] & ~io_in[8] & io_in[9] & io_in[10]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & io_in[6] & io_in[7] & ~io_in[8] & io_in[10]) | (io_in[0] & ~io_in[1] & ~io_in[3] & io_in[5] & io_in[7] & ~io_in[9] & ~io_in[11]) | (io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & io_in[6] & ~io_in[7] & io_in[8] & ~io_in[9]) | (io_in[0] & ~io_in[1] & io_in[3] & ~io_in[4] & ~io_in[6] & io_in[7] & io_in[8] & ~io_in[9] & io_in[11]) | (~io_in[0] & io_in[1] & io_in[2] & ~io_in[3] & io_in[4] & io_in[6] & ~io_in[7] & io_in[8] & io_in[9]) | (~io_in[0] & io_in[1] & io_in[2] & io_in[3] & io_in[4] & ~io_in[6] & io_in[7] & io_in[10]) | (io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[4] & io_in[6] & io_in[7] & ~io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & io_in[1] & io_in[2] & io_in[3] & ~io_in[6] & ~io_in[7] & ~io_in[8] & io_in[9]) | (~io_in[0] & ~io_in[2] & ~io_in[3] & io_in[4] & io_in[6] & ~io_in[7] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[6] & io_in[7] & ~io_in[9] & ~io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & io_in[4] & io_in[6] & ~io_in[7] & io_in[8] & ~io_in[9] & ~io_in[11]) | (~io_in[0] & io_in[1] & io_in[2] & io_in[3] & ~io_in[6] & ~io_in[7] & ~io_in[8] & ~io_in[9]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[6] & ~io_in[7] & io_in[8] & ~io_in[9] & io_in[10]) | (~io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & ~io_in[5] & ~io_in[7] & ~io_in[8] & io_in[9] & io_in[10]) | (io_in[0] & io_in[2] & io_in[3] & ~io_in[5] & ~io_in[6] & io_in[7] & ~io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & ~io_in[6] & io_in[7] & io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & ~io_in[1] & ~io_in[2] & io_in[3] & io_in[4] & ~io_in[6] & ~io_in[7] & io_in[9] & io_in[11]) | (io_in[0] & io_in[1] & ~io_in[2] & io_in[3] & ~io_in[4] & io_in[6] & ~io_in[8] & io_in[9] & io_in[10]) | (io_in[0] & io_in[2] & io_in[3] & io_in[6] & ~io_in[7] & ~io_in[8] & ~io_in[9] & io_in[10]) | (~io_in[0] & io_in[1] & io_in[2] & io_in[4] & io_in[8] & ~io_in[9] & ~io_in[10]) | (~io_in[0] & io_in[1] & io_in[2] & io_in[3] & io_in[5] & ~io_in[6]) | (io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[6] & io_in[7] & io_in[8] & io_in[10]) | (io_in[0] & io_in[1] & ~io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[6] & io_in[7] & ~io_in[8] & io_in[9] & ~io_in[11]) | (~io_in[0] & ~io_in[2] & ~io_in[3] & ~io_in[4] & io_in[6] & io_in[7] & io_in[8] & io_in[9] & io_in[10] & ~io_in[11]) | (io_in[0] & io_in[1] & ~io_in[3] & io_in[4] & io_in[6] & ~io_in[7] & ~io_in[8] & ~io_in[9] & io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & ~io_in[5] & io_in[6] & ~io_in[7] & io_in[10] & io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & io_in[3] & ~io_in[4] & io_in[6] & ~io_in[7] & io_in[8] & ~io_in[9]) | (~io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & io_in[6] & io_in[8] & ~io_in[9] & io_in[10]) | (~io_in[0] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[6] & io_in[7] & ~io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & io_in[1] & ~io_in[3] & io_in[6] & io_in[7] & io_in[8] & ~io_in[9] & io_in[10]) | (io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & ~io_in[6] & ~io_in[7] & ~io_in[8] & io_in[10]) | (io_in[0] & io_in[1] & io_in[2] & ~io_in[3] & io_in[4] & io_in[6] & io_in[7] & io_in[8] & io_in[9] & ~io_in[10]) | (~io_in[0] & io_in[1] & io_in[2] & io_in[4] & ~io_in[5] & ~io_in[6] & io_in[7] & io_in[8] & io_in[11]) | (io_in[0] & ~io_in[1] & ~io_in[2] & io_in[6] & io_in[7] & io_in[9] & ~io_in[10] & io_in[11]) | (io_in[0] & ~io_in[1] & io_in[2] & io_in[4] & io_in[6] & io_in[7] & io_in[10] & io_in[11]) | (~io_in[0] & ~io_in[1] & io_in[5] & io_in[6] & io_in[8] & ~io_in[9]) | (~io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & io_in[6] & ~io_in[8] & io_in[9] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[1] & io_in[2] & io_in[4] & io_in[6] & ~io_in[7] & io_in[8] & io_in[9] & io_in[10]) | (~io_in[0] & ~io_in[1] & io_in[2] & io_in[4] & io_in[7] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (io_in[0] & io_in[1] & io_in[2] & io_in[3] & ~io_in[6] & io_in[7] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (io_in[0] & io_in[5] & io_in[6] & io_in[9] & ~io_in[10] & io_in[11]) | (io_in[0] & ~io_in[2] & io_in[3] & io_in[5] & io_in[7] & io_in[8] & io_in[10]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & ~io_in[6] & ~io_in[7] & ~io_in[8] & ~io_in[9] & io_in[11]) | (~io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & io_in[6] & io_in[7] & ~io_in[8] & io_in[9] & io_in[10]) | (~io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[6] & io_in[7] & io_in[10] & io_in[11]) | (io_in[0] & ~io_in[1] & ~io_in[2] & io_in[3] & io_in[4] & io_in[7] & io_in[8] & io_in[10] & ~io_in[11]) | (io_in[0] & io_in[2] & io_in[5] & ~io_in[6] & io_in[8] & ~io_in[10]) | (io_in[0] & ~io_in[1] & ~io_in[2] & io_in[5] & ~io_in[7] & io_in[9] & ~io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & io_in[3] & io_in[4] & io_in[6] & ~io_in[7] & io_in[8] & io_in[9] & ~io_in[10]) | (io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & io_in[4] & ~io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[6] & ~io_in[7] & io_in[9] & ~io_in[10]) | (io_in[1] & io_in[2] & io_in[3] & ~io_in[7] & ~io_in[8] & ~io_in[10] & ~io_in[11]) | (io_in[0] & ~io_in[1] & ~io_in[3] & io_in[4] & ~io_in[6] & ~io_in[7] & ~io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & io_in[4] & io_in[6] & ~io_in[7] & ~io_in[8] & ~io_in[11]) | (io_in[0] & io_in[1] & io_in[2] & io_in[3] & io_in[6] & ~io_in[8] & io_in[9] & ~io_in[10]) | (~io_in[0] & io_in[1] & ~io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[6] & io_in[7] & ~io_in[8] & ~io_in[9] & io_in[11]) | (io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[6] & io_in[7] & ~io_in[8] & io_in[9] & io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[3] & ~io_in[4] & ~io_in[6] & io_in[7] & ~io_in[8] & ~io_in[9] & io_in[10] & ~io_in[11]) | (io_in[0] & io_in[1] & io_in[2] & io_in[5] & io_in[7] & ~io_in[8] & io_in[9]) | (io_in[0] & io_in[1] & ~io_in[2] & io_in[3] & io_in[5] & io_in[6] & io_in[9] & io_in[10]) | (io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[7] & io_in[8] & ~io_in[10]) | (io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[6] & ~io_in[7] & ~io_in[10] & io_in[11]) | (io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[4] & ~io_in[5] & io_in[6] & ~io_in[7] & io_in[8] & io_in[9] & io_in[10]) | (io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[8] & io_in[9] & io_in[10] & ~io_in[11]) | (~io_in[0] & ~io_in[1] & io_in[2] & io_in[4] & ~io_in[6] & ~io_in[7] & io_in[9] & io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[2] & io_in[4] & io_in[5] & ~io_in[7]) | (~io_in[0] & io_in[1] & ~io_in[2] & io_in[3] & io_in[4] & ~io_in[6] & io_in[8] & io_in[9] & ~io_in[10]) | (~io_in[1] & io_in[2] & ~io_in[3] & io_in[5] & ~io_in[8] & ~io_in[9] & io_in[10]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & io_in[3] & ~io_in[4] & io_in[6] & ~io_in[8] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & ~io_in[1] & io_in[2] & io_in[4] & io_in[6] & ~io_in[8] & io_in[9] & io_in[11]) | (~io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & io_in[8] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (io_in[0] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[7] & ~io_in[8] & ~io_in[10] & ~io_in[11]) | (io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[8] & io_in[9] & ~io_in[10] & ~io_in[11]) | (io_in[1] & ~io_in[2] & io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[6] & ~io_in[7] & io_in[8] & io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[6] & io_in[7] & ~io_in[9]) | (io_in[0] & ~io_in[1] & ~io_in[2] & io_in[3] & ~io_in[4] & ~io_in[7] & ~io_in[8] & io_in[10]) | (io_in[0] & io_in[1] & ~io_in[2] & io_in[3] & io_in[6] & io_in[7] & ~io_in[10] & io_in[11]) | (~io_in[1] & ~io_in[2] & io_in[3] & io_in[4] & io_in[6] & io_in[7] & ~io_in[8] & io_in[9] & ~io_in[10]) | (io_in[0] & io_in[1] & ~io_in[2] & io_in[4] & ~io_in[6] & ~io_in[7] & io_in[8] & ~io_in[9] & ~io_in[10]) | (io_in[1] & io_in[2] & ~io_in[3] & io_in[4] & ~io_in[6] & ~io_in[8] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & io_in[6] & ~io_in[7] & ~io_in[9] & ~io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & io_in[4] & io_in[7] & io_in[9] & ~io_in[10] & io_in[11]) | (~io_in[0] & io_in[1] & io_in[2] & io_in[3] & io_in[4] & ~io_in[6] & io_in[8] & ~io_in[9]) | (io_in[0] & io_in[1] & io_in[3] & io_in[4] & io_in[6] & io_in[8] & ~io_in[9] & io_in[11]) | (io_in[2] & io_in[3] & io_in[4] & ~io_in[6] & io_in[7] & ~io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & ~io_in[1] & ~io_in[2] & io_in[4] & ~io_in[5] & io_in[6] & io_in[7] & io_in[9] & io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & io_in[7] & io_in[8] & io_in[9] & io_in[10] & ~io_in[11]) | (io_in[0] & io_in[3] & io_in[4] & io_in[6] & io_in[7] & ~io_in[8] & io_in[9]) | (~io_in[0] & io_in[1] & ~io_in[2] & io_in[3] & ~io_in[5] & io_in[6] & ~io_in[7] & ~io_in[8] & ~io_in[9] & ~io_in[10]) | (io_in[0] & ~io_in[1] & ~io_in[3] & io_in[4] & io_in[6] & io_in[7] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (io_in[0] & ~io_in[1] & ~io_in[2] & io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & ~io_in[7] & ~io_in[8] & ~io_in[9] & io_in[11]) | (io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & io_in[4] & ~io_in[5] & io_in[6] & io_in[10] & io_in[11]) | (io_in[0] & io_in[1] & io_in[3] & ~io_in[4] & ~io_in[6] & io_in[7] & io_in[8] & io_in[9] & ~io_in[11]) | (io_in[1] & ~io_in[2] & io_in[3] & io_in[5] & ~io_in[6] & io_in[7] & ~io_in[9]) | (io_in[0] & io_in[1] & ~io_in[2] & io_in[3] & ~io_in[4] & ~io_in[8] & io_in[9] & io_in[11]) | (~io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & io_in[5] & ~io_in[6] & io_in[7] & io_in[11]) | (io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[6] & ~io_in[7] & io_in[8] & io_in[11]) | (io_in[0] & io_in[1] & io_in[3] & io_in[5] & io_in[7] & io_in[11]) | (io_in[0] & io_in[1] & io_in[2] & ~io_in[3] & io_in[4] & io_in[6] & ~io_in[7] & ~io_in[8] & io_in[10]) | (io_in[0] & io_in[2] & io_in[3] & ~io_in[6] & io_in[7] & io_in[8] & io_in[9] & io_in[10] & ~io_in[11]) | (~io_in[1] & io_in[2] & ~io_in[3] & io_in[5] & io_in[7] & io_in[8] & io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[1] & io_in[5] & io_in[6] & ~io_in[7] & io_in[8] & ~io_in[11]) | (io_in[0] & io_in[2] & io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & ~io_in[7] & io_in[10] & io_in[11]) | (io_in[0] & ~io_in[1] & ~io_in[3] & io_in[6] & io_in[7] & ~io_in[8] & io_in[9] & io_in[10]) | (io_in[0] & ~io_in[1] & ~io_in[2] & io_in[3] & io_in[8] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & ~io_in[6] & ~io_in[7] & io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & ~io_in[2] & io_in[3] & io_in[4] & io_in[6] & io_in[7] & ~io_in[8] & io_in[10]) | (io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & io_in[4] & io_in[7] & ~io_in[8] & io_in[11]) | (~io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & ~io_in[7] & io_in[8] & ~io_in[9] & io_in[11]) | (io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & io_in[8] & io_in[9] & io_in[10]) | (~io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & io_in[4] & io_in[6] & ~io_in[7] & ~io_in[10] & io_in[11]) | (io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & io_in[6] & ~io_in[8] & io_in[9] & io_in[10]) | (io_in[0] & io_in[1] & io_in[2] & ~io_in[3] & io_in[4] & ~io_in[6] & ~io_in[7] & io_in[8] & io_in[9] & io_in[10] & ~io_in[11]) | (io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & io_in[6] & ~io_in[7] & io_in[8] & ~io_in[10]) | (io_in[0] & io_in[1] & io_in[2] & io_in[4] & io_in[6] & ~io_in[7] & ~io_in[10] & io_in[11]) | (io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[6] & io_in[8] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[1] & io_in[3] & io_in[4] & ~io_in[6] & io_in[7] & ~io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & ~io_in[1] & ~io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[6] & io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & io_in[1] & ~io_in[2] & io_in[3] & io_in[6] & ~io_in[7] & io_in[8] & ~io_in[10] & ~io_in[11]) | (~io_in[1] & io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & io_in[7] & ~io_in[8] & ~io_in[9] & io_in[10]) | (~io_in[0] & io_in[2] & io_in[3] & io_in[4] & io_in[6] & ~io_in[7] & io_in[10] & io_in[11]) | (io_in[1] & io_in[3] & io_in[4] & io_in[6] & ~io_in[7] & io_in[8] & ~io_in[9] & io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & ~io_in[7] & io_in[9] & io_in[10] & ~io_in[11]) | (io_in[0] & io_in[1] & io_in[5] & ~io_in[6] & ~io_in[7] & ~io_in[8] & io_in[10]) | (io_in[0] & io_in[1] & io_in[2] & ~io_in[4] & ~io_in[6] & ~io_in[7] & io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & io_in[1] & ~io_in[2] & io_in[3] & io_in[4] & ~io_in[6] & ~io_in[7] & ~io_in[8] & ~io_in[9]) | (~io_in[0] & ~io_in[1] & io_in[3] & io_in[4] & io_in[7] & io_in[8] & ~io_in[9] & io_in[11]) | (io_in[1] & io_in[2] & io_in[4] & io_in[5] & ~io_in[7]) | (~io_in[0] & ~io_in[1] & io_in[2] & io_in[5] & io_in[6] & ~io_in[7] & io_in[9] & io_in[11]) | (io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & ~io_in[6] & ~io_in[8] & ~io_in[9] & io_in[11]) | (~io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & io_in[6] & ~io_in[8] & ~io_in[9] & io_in[10]) | (~io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & io_in[4] & ~io_in[6] & io_in[9] & ~io_in[10] & ~io_in[11]) | (io_in[0] & ~io_in[1] & ~io_in[3] & io_in[4] & ~io_in[6] & ~io_in[7] & io_in[8] & ~io_in[9] & ~io_in[10]) | (io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & io_in[4] & ~io_in[6] & ~io_in[7] & ~io_in[9] & io_in[10]) | (io_in[0] & io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[7] & ~io_in[8] & ~io_in[9] & io_in[10]) | (~io_in[0] & io_in[1] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & io_in[10] & io_in[11]) | (io_in[0] & ~io_in[2] & io_in[3] & ~io_in[4] & ~io_in[5] & io_in[7] & io_in[8] & io_in[9] & ~io_in[10]) | (~io_in[0] & ~io_in[1] & ~io_in[3] & io_in[5] & ~io_in[6] & ~io_in[7] & ~io_in[9] & ~io_in[11]) | (io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & ~io_in[6] & io_in[7] & ~io_in[8] & ~io_in[9] & ~io_in[10]) | (io_in[0] & io_in[1] & io_in[2] & io_in[4] & io_in[7] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (~io_in[1] & ~io_in[2] & io_in[5] & io_in[7] & ~io_in[8] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[1] & io_in[2] & ~io_in[3] & ~io_in[5] & ~io_in[6] & ~io_in[7] & io_in[8] & ~io_in[9] & ~io_in[10]) | (~io_in[0] & ~io_in[2] & io_in[3] & io_in[4] & ~io_in[6] & ~io_in[7] & ~io_in[8] & io_in[9] & io_in[10]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & io_in[5] & ~io_in[6] & io_in[7] & io_in[8] & io_in[9]) | (io_in[0] & io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[6] & io_in[7] & io_in[8] & io_in[11]) | (io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & io_in[4] & ~io_in[7] & ~io_in[9] & io_in[11]) | (~io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[6] & ~io_in[8] & io_in[9] & io_in[10]) | (~io_in[0] & io_in[1] & io_in[2] & io_in[4] & io_in[7] & ~io_in[8] & ~io_in[9] & io_in[10]) | (~io_in[0] & io_in[1] & io_in[2] & io_in[3] & io_in[4] & io_in[7] & io_in[8] & io_in[11]) | (io_in[0] & io_in[1] & ~io_in[2] & io_in[3] & io_in[4] & io_in[7] & io_in[8] & io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & io_in[5] & io_in[7] & io_in[9] & ~io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & io_in[3] & ~io_in[4] & ~io_in[5] & io_in[7] & ~io_in[8] & ~io_in[9] & ~io_in[11]) | (~io_in[0] & io_in[2] & io_in[3] & ~io_in[4] & ~io_in[6] & io_in[8] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (io_in[0] & ~io_in[2] & ~io_in[3] & ~io_in[6] & io_in[7] & io_in[8] & io_in[9] & io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & io_in[3] & ~io_in[4] & io_in[7] & io_in[8] & ~io_in[9] & io_in[10]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[6] & ~io_in[7] & ~io_in[8] & io_in[9]) | (~io_in[0] & ~io_in[1] & io_in[3] & io_in[4] & ~io_in[6] & io_in[7] & io_in[8] & io_in[11]) | (io_in[0] & ~io_in[1] & ~io_in[2] & io_in[3] & ~io_in[4] & ~io_in[6] & io_in[9] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & io_in[6] & io_in[7] & io_in[8] & io_in[9] & ~io_in[11]) | (~io_in[1] & ~io_in[2] & io_in[3] & ~io_in[4] & ~io_in[6] & io_in[7] & io_in[8] & io_in[9] & ~io_in[10]) | (io_in[0] & ~io_in[1] & io_in[2] & io_in[5] & ~io_in[7] & ~io_in[9] & io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & io_in[5] & ~io_in[7] & io_in[8] & io_in[11]) | (io_in[0] & io_in[1] & io_in[2] & io_in[4] & ~io_in[7] & ~io_in[8] & io_in[11]) | (io_in[0] & ~io_in[1] & ~io_in[2] & io_in[5] & io_in[6] & io_in[7] & ~io_in[8] & ~io_in[9]) | (~io_in[0] & ~io_in[2] & io_in[3] & ~io_in[6] & io_in[7] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & ~io_in[7] & io_in[8] & ~io_in[9] & ~io_in[10]) | (~io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & ~io_in[5] & io_in[6] & io_in[7] & io_in[8] & ~io_in[10]) | (io_in[1] & ~io_in[2] & io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & io_in[7] & ~io_in[8] & io_in[9] & io_in[10]) | (~io_in[0] & ~io_in[2] & ~io_in[3] & io_in[5] & io_in[6] & ~io_in[7] & ~io_in[9] & io_in[11]) | (~io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[6] & ~io_in[7] & ~io_in[8] & io_in[9]) | (io_in[1] & io_in[2] & io_in[3] & io_in[6] & io_in[7] & ~io_in[8] & io_in[9] & io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & ~io_in[7] & io_in[9] & io_in[11]) | (~io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & ~io_in[7] & io_in[8] & io_in[10] & ~io_in[11]) | (io_in[0] & io_in[1] & ~io_in[2] & ~io_in[4] & ~io_in[5] & io_in[6] & io_in[7] & ~io_in[8] & io_in[11]) | (~io_in[0] & io_in[1] & io_in[2] & ~io_in[3] & ~io_in[5] & ~io_in[6] & ~io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[6] & ~io_in[8] & io_in[9] & ~io_in[10] & ~io_in[11]) | (io_in[0] & io_in[1] & ~io_in[2] & io_in[3] & io_in[4] & ~io_in[6] & io_in[7] & io_in[8] & io_in[10]) | (io_in[0] & io_in[1] & ~io_in[2] & io_in[3] & io_in[4] & io_in[7] & ~io_in[9] & ~io_in[10]) | (~io_in[0] & ~io_in[2] & ~io_in[3] & io_in[4] & io_in[6] & io_in[7] & io_in[8] & ~io_in[9]) | (~io_in[0] & ~io_in[1] & io_in[2] & io_in[5] & io_in[8] & ~io_in[9]) | (io_in[0] & io_in[1] & ~io_in[2] & io_in[3] & ~io_in[6] & io_in[7] & io_in[10] & io_in[11]) | (io_in[0] & io_in[1] & ~io_in[2] & io_in[5] & io_in[8] & io_in[9] & io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & io_in[3] & ~io_in[4] & io_in[6] & ~io_in[7] & io_in[8] & io_in[9] & ~io_in[11]) | (io_in[0] & io_in[1] & ~io_in[2] & io_in[3] & ~io_in[6] & ~io_in[7] & ~io_in[9] & io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[5] & ~io_in[6] & ~io_in[7] & io_in[8] & io_in[9] & ~io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & io_in[7] & io_in[11]) | (io_in[0] & ~io_in[1] & io_in[2] & io_in[5] & io_in[8] & io_in[9] & io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & ~io_in[6] & ~io_in[8] & io_in[9] & ~io_in[10] & ~io_in[11]) | (io_in[0] & ~io_in[1] & ~io_in[2] & io_in[4] & io_in[5] & ~io_in[6] & ~io_in[7]) | (io_in[0] & io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & io_in[7] & ~io_in[9] & ~io_in[11]);

assign val[4] = (~io_in[0] & io_in[2] & ~io_in[3] & ~io_in[4] & io_in[6] & io_in[7] & io_in[9] & ~io_in[10] & io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[6] & ~io_in[8] & io_in[9] & io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[1] & io_in[2] & ~io_in[3] & ~io_in[6] & io_in[7] & io_in[8] & io_in[10] & ~io_in[11]) | (~io_in[1] & ~io_in[2] & ~io_in[4] & ~io_in[5] & ~io_in[6] & ~io_in[7] & io_in[8] & io_in[9] & io_in[10] & io_in[11]) | (io_in[0] & io_in[2] & io_in[3] & ~io_in[4] & io_in[6] & io_in[7] & ~io_in[8] & ~io_in[9] & io_in[11]) | (io_in[0] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & io_in[8] & io_in[9] & ~io_in[10]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[4] & io_in[6] & ~io_in[7] & io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & ~io_in[1] & ~io_in[2] & io_in[5] & ~io_in[7] & io_in[8] & ~io_in[9] & io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & ~io_in[7] & io_in[8] & io_in[9] & ~io_in[11]) | (io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & io_in[5] & io_in[6] & ~io_in[8] & ~io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & io_in[7] & io_in[8] & ~io_in[9]) | (io_in[0] & ~io_in[1] & io_in[2] & ~io_in[4] & io_in[6] & ~io_in[7] & ~io_in[8] & ~io_in[9] & io_in[10]) | (~io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[8] & ~io_in[9] & io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & io_in[3] & io_in[4] & io_in[6] & ~io_in[7] & ~io_in[8] & io_in[9]) | (io_in[0] & io_in[1] & ~io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[6] & io_in[7] & ~io_in[9] & io_in[10]) | (~io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & ~io_in[6] & io_in[7] & ~io_in[8] & io_in[9] & io_in[10]) | (io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & io_in[6] & io_in[10] & io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & io_in[4] & ~io_in[6] & ~io_in[7] & io_in[8] & ~io_in[10] & io_in[11]) | (~io_in[0] & io_in[1] & io_in[2] & ~io_in[3] & io_in[5] & io_in[6] & io_in[7] & io_in[9] & ~io_in[11]) | (~io_in[1] & io_in[2] & io_in[3] & io_in[4] & ~io_in[6] & io_in[7] & io_in[9] & io_in[10] & ~io_in[11]) | (io_in[0] & io_in[1] & ~io_in[2] & ~io_in[4] & ~io_in[6] & ~io_in[7] & io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & io_in[1] & io_in[2] & io_in[3] & ~io_in[6] & io_in[7] & io_in[8] & ~io_in[9] & io_in[11]) | (io_in[0] & ~io_in[1] & ~io_in[2] & io_in[3] & ~io_in[4] & io_in[6] & ~io_in[7] & io_in[8] & io_in[10] & ~io_in[11]) | (io_in[0] & io_in[1] & io_in[2] & ~io_in[3] & ~io_in[5] & ~io_in[6] & io_in[7] & ~io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[7] & ~io_in[8] & ~io_in[9] & io_in[11]) | (io_in[0] & ~io_in[2] & io_in[3] & io_in[4] & io_in[6] & io_in[7] & io_in[8] & io_in[9] & ~io_in[10]) | (io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & io_in[5] & io_in[6] & io_in[7] & ~io_in[8]) | (io_in[0] & ~io_in[1] & io_in[3] & io_in[4] & io_in[6] & ~io_in[7] & ~io_in[8] & io_in[11]) | (io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & io_in[5] & ~io_in[7] & io_in[10] & io_in[11]) | (io_in[0] & io_in[1] & ~io_in[2] & io_in[3] & io_in[4] & io_in[6] & ~io_in[7] & ~io_in[9] & io_in[10]) | (io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & io_in[6] & io_in[7] & ~io_in[9] & io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & io_in[5] & ~io_in[6] & io_in[7] & ~io_in[8] & io_in[9] & io_in[10]) | (io_in[0] & ~io_in[1] & ~io_in[2] & io_in[4] & io_in[6] & ~io_in[7] & ~io_in[8] & ~io_in[9] & io_in[10]) | (~io_in[0] & io_in[1] & ~io_in[2] & io_in[3] & ~io_in[5] & ~io_in[6] & io_in[7] & ~io_in[8] & io_in[9] & io_in[10]) | (io_in[0] & io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & ~io_in[7] & io_in[8] & io_in[9] & io_in[10]) | (io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & io_in[6] & ~io_in[7] & io_in[9] & io_in[11]) | (~io_in[0] & io_in[1] & io_in[2] & io_in[3] & io_in[4] & io_in[6] & io_in[7] & ~io_in[8] & io_in[9]) | (~io_in[0] & io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & io_in[6] & io_in[7] & ~io_in[8] & io_in[9] & ~io_in[10]) | (io_in[2] & io_in[3] & io_in[4] & io_in[6] & io_in[7] & io_in[10] & io_in[11]) | (~io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & io_in[6] & io_in[7] & ~io_in[8] & ~io_in[10] & ~io_in[11]) | (io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & ~io_in[5] & io_in[6] & ~io_in[7] & io_in[8] & io_in[9] & io_in[10]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & ~io_in[6] & io_in[7] & io_in[9] & ~io_in[10] & ~io_in[11]) | (io_in[0] & io_in[2] & io_in[4] & ~io_in[5] & ~io_in[6] & ~io_in[7] & io_in[10] & io_in[11]) | (~io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & ~io_in[6] & ~io_in[8] & io_in[9] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[1] & io_in[2] & ~io_in[3] & io_in[4] & io_in[6] & ~io_in[7] & io_in[9] & ~io_in[11]) | (~io_in[0] & ~io_in[1] & io_in[2] & ~io_in[4] & ~io_in[5] & io_in[6] & io_in[7] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & io_in[4] & ~io_in[5] & ~io_in[6] & io_in[7] & io_in[10] & io_in[11]) | (~io_in[0] & io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & ~io_in[7] & io_in[10] & io_in[11]) | (~io_in[0] & io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & ~io_in[6] & ~io_in[7] & io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & io_in[7] & ~io_in[8] & io_in[9] & io_in[10]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & io_in[6] & io_in[7] & ~io_in[8] & io_in[10]) | (~io_in[0] & io_in[1] & ~io_in[2] & io_in[3] & io_in[4] & io_in[7] & ~io_in[8] & ~io_in[9] & io_in[10]) | (~io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & io_in[4] & io_in[7] & ~io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & io_in[1] & ~io_in[2] & ~io_in[4] & ~io_in[6] & io_in[7] & io_in[8] & io_in[9] & io_in[10] & ~io_in[11]) | (io_in[0] & io_in[1] & ~io_in[3] & ~io_in[4] & ~io_in[6] & ~io_in[7] & ~io_in[8] & io_in[9] & io_in[10]) | (io_in[0] & ~io_in[1] & ~io_in[2] & io_in[3] & io_in[4] & ~io_in[7] & io_in[8] & io_in[9] & io_in[10] & ~io_in[11]) | (~io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & ~io_in[7] & ~io_in[8] & ~io_in[10]) | (~io_in[0] & io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[6] & ~io_in[7] & io_in[9] & io_in[11]) | (io_in[0] & io_in[2] & io_in[3] & io_in[4] & ~io_in[6] & io_in[7] & ~io_in[8] & io_in[9] & io_in[10]) | (~io_in[0] & io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & io_in[6] & ~io_in[7] & ~io_in[8] & io_in[9] & io_in[10]) | (io_in[0] & ~io_in[1] & io_in[2] & ~io_in[4] & ~io_in[5] & io_in[6] & io_in[7] & ~io_in[8] & ~io_in[9] & io_in[11]) | (~io_in[0] & io_in[2] & ~io_in[3] & io_in[4] & ~io_in[6] & io_in[7] & io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & io_in[6] & io_in[8] & ~io_in[10] & io_in[11]) | (~io_in[0] & io_in[1] & io_in[2] & ~io_in[3] & io_in[5] & io_in[6] & ~io_in[7] & io_in[8] & io_in[11]) | (~io_in[0] & io_in[1] & io_in[2] & ~io_in[3] & ~io_in[5] & io_in[7] & ~io_in[8] & ~io_in[9] & io_in[11]) | (io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[6] & io_in[7] & ~io_in[8] & ~io_in[9]) | (~io_in[1] & ~io_in[2] & io_in[3] & ~io_in[4] & io_in[6] & ~io_in[7] & io_in[8] & io_in[9] & io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[3] & ~io_in[4] & io_in[8] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & ~io_in[6] & io_in[8] & io_in[9] & io_in[10] & ~io_in[11]) | (io_in[0] & io_in[1] & ~io_in[3] & io_in[4] & ~io_in[5] & ~io_in[7] & io_in[10] & io_in[11]) | (~io_in[0] & io_in[1] & io_in[2] & ~io_in[5] & ~io_in[6] & ~io_in[7] & io_in[10] & io_in[11]) | (io_in[0] & io_in[1] & io_in[2] & ~io_in[3] & io_in[5] & ~io_in[6] & io_in[7] & io_in[11]) | (io_in[0] & ~io_in[1] & ~io_in[2] & io_in[3] & ~io_in[4] & io_in[6] & io_in[8] & ~io_in[10] & io_in[11]) | (~io_in[0] & io_in[1] & io_in[2] & ~io_in[3] & io_in[4] & ~io_in[8] & ~io_in[9] & io_in[11]) | (~io_in[0] & ~io_in[1] & io_in[2] & io_in[5] & io_in[6] & io_in[7] & ~io_in[8] & io_in[11]) | (io_in[1] & ~io_in[2] & io_in[3] & io_in[4] & io_in[6] & io_in[7] & io_in[8] & io_in[9] & io_in[10]) | (~io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & ~io_in[6] & io_in[7] & ~io_in[8] & io_in[10]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[4] & ~io_in[5] & io_in[6] & io_in[8] & io_in[9] & io_in[10] & io_in[11]) | (io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & ~io_in[7] & io_in[8] & io_in[9] & io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[6] & io_in[10] & io_in[11]) | (~io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & io_in[4] & ~io_in[8] & io_in[9] & ~io_in[10] & ~io_in[11]) | (io_in[0] & io_in[1] & ~io_in[2] & ~io_in[4] & io_in[6] & io_in[7] & ~io_in[8] & ~io_in[9] & io_in[10]) | (~io_in[0] & io_in[1] & io_in[3] & io_in[4] & ~io_in[6] & io_in[7] & io_in[8] & io_in[9] & ~io_in[10]) | (io_in[0] & ~io_in[1] & io_in[3] & ~io_in[4] & io_in[5] & ~io_in[6] & ~io_in[7]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[6] & io_in[7] & ~io_in[8] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[1] & io_in[2] & io_in[3] & io_in[4] & ~io_in[6] & ~io_in[7] & io_in[9] & io_in[10]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & io_in[5] & io_in[6] & io_in[7] & io_in[8]) | (io_in[0] & ~io_in[1] & ~io_in[4] & ~io_in[6] & io_in[7] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (io_in[0] & ~io_in[1] & io_in[2] & ~io_in[4] & io_in[5] & ~io_in[7] & io_in[9] & io_in[11]) | (io_in[0] & ~io_in[2] & ~io_in[3] & io_in[5] & io_in[6] & io_in[7] & ~io_in[9] & io_in[10]) | (io_in[0] & io_in[2] & io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & io_in[7] & ~io_in[8] & io_in[9] & io_in[10]) | (~io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & io_in[5] & ~io_in[6] & ~io_in[7] & io_in[10] & io_in[11]) | (~io_in[0] & io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & ~io_in[5] & io_in[7] & ~io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & io_in[1] & io_in[2] & io_in[3] & io_in[4] & ~io_in[6] & io_in[7] & ~io_in[10]) | (io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[5] & ~io_in[6] & io_in[7] & ~io_in[8] & io_in[10]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & ~io_in[6] & ~io_in[7] & ~io_in[8] & io_in[9] & io_in[10]) | (io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & io_in[6] & io_in[7] & ~io_in[8] & ~io_in[9] & io_in[10]) | (~io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & io_in[6] & ~io_in[7] & io_in[8] & ~io_in[9] & io_in[10]) | (~io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[6] & io_in[7] & io_in[8] & ~io_in[9] & ~io_in[10] & io_in[11]) | (~io_in[0] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[6] & ~io_in[7] & ~io_in[10] & ~io_in[11]) | (io_in[0] & io_in[1] & ~io_in[2] & io_in[4] & ~io_in[6] & io_in[7] & ~io_in[8] & io_in[9] & io_in[11]) | (~io_in[0] & io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & io_in[6] & ~io_in[7] & ~io_in[9] & io_in[11]) | (io_in[0] & io_in[1] & io_in[3] & io_in[4] & ~io_in[6] & ~io_in[7] & ~io_in[9] & io_in[11]) | (~io_in[0] & io_in[1] & io_in[2] & ~io_in[3] & io_in[4] & io_in[7] & ~io_in[10] & io_in[11]) | (~io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & io_in[4] & ~io_in[6] & io_in[8] & ~io_in[9] & io_in[10]) | (~io_in[0] & ~io_in[2] & ~io_in[3] & io_in[4] & ~io_in[6] & ~io_in[7] & io_in[8] & ~io_in[10] & io_in[11]) | (io_in[0] & io_in[1] & ~io_in[2] & io_in[3] & ~io_in[5] & ~io_in[6] & ~io_in[8] & ~io_in[9] & ~io_in[10]) | (io_in[0] & io_in[3] & io_in[4] & ~io_in[6] & io_in[7] & io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & ~io_in[1] & io_in[3] & ~io_in[4] & ~io_in[5] & io_in[7] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & io_in[6] & io_in[7] & ~io_in[8] & io_in[11]) | (io_in[0] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[6] & ~io_in[7] & ~io_in[8] & io_in[9] & io_in[10]) | (io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & io_in[4] & io_in[6] & io_in[7] & ~io_in[9] & ~io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & ~io_in[6] & ~io_in[7] & io_in[8] & io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & io_in[6] & io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & ~io_in[1] & ~io_in[2] & io_in[3] & ~io_in[4] & io_in[6] & io_in[7] & ~io_in[8] & io_in[9] & io_in[10]) | (io_in[0] & io_in[1] & ~io_in[2] & io_in[3] & ~io_in[6] & ~io_in[7] & ~io_in[8] & ~io_in[9]) | (~io_in[0] & ~io_in[2] & ~io_in[3] & io_in[5] & ~io_in[6] & ~io_in[8] & ~io_in[9] & io_in[11]) | (io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[6] & io_in[7] & io_in[10] & io_in[11]) | (io_in[0] & io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & io_in[6] & ~io_in[7] & io_in[8] & ~io_in[9] & io_in[10]) | (~io_in[1] & io_in[2] & ~io_in[3] & io_in[4] & ~io_in[6] & io_in[7] & ~io_in[8] & ~io_in[9] & io_in[11]) | (io_in[0] & io_in[2] & io_in[5] & io_in[6] & io_in[8] & ~io_in[9]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[6] & io_in[7] & io_in[9] & ~io_in[11]) | (io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & ~io_in[8] & ~io_in[9] & io_in[10]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & io_in[3] & ~io_in[5] & io_in[6] & ~io_in[7] & io_in[10] & io_in[11]) | (io_in[0] & io_in[1] & io_in[3] & ~io_in[4] & io_in[6] & ~io_in[7] & ~io_in[8] & ~io_in[9] & io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & io_in[3] & io_in[4] & ~io_in[6] & io_in[7] & io_in[8] & io_in[11]) | (~io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & ~io_in[6] & ~io_in[7] & ~io_in[8] & io_in[9] & io_in[11]) | (io_in[1] & ~io_in[2] & io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[6] & io_in[7] & ~io_in[8] & ~io_in[9] & io_in[11]) | (io_in[0] & io_in[1] & io_in[2] & ~io_in[3] & io_in[4] & ~io_in[6] & io_in[7] & io_in[8] & io_in[9]) | (~io_in[0] & io_in[1] & ~io_in[2] & io_in[5] & ~io_in[6] & ~io_in[7] & ~io_in[8] & io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & io_in[3] & io_in[4] & io_in[6] & io_in[7] & ~io_in[8] & io_in[11]) | (io_in[1] & io_in[2] & io_in[3] & io_in[6] & io_in[7] & io_in[10] & io_in[11]) | (io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & io_in[4] & ~io_in[7] & ~io_in[8] & io_in[9] & io_in[10]) | (io_in[0] & ~io_in[1] & io_in[2] & io_in[5] & ~io_in[7] & ~io_in[9] & io_in[10]) | (~io_in[0] & io_in[1] & io_in[2] & io_in[3] & io_in[4] & io_in[7] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[1] & io_in[2] & io_in[4] & ~io_in[6] & io_in[8] & io_in[9] & io_in[10] & ~io_in[11]) | (io_in[0] & ~io_in[1] & io_in[3] & ~io_in[4] & io_in[7] & ~io_in[8] & io_in[9] & io_in[11]) | (~io_in[0] & io_in[1] & io_in[2] & ~io_in[6] & io_in[7] & io_in[8] & io_in[9] & io_in[10] & ~io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[6] & ~io_in[8] & ~io_in[9] & io_in[11]) | (~io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & io_in[4] & ~io_in[6] & ~io_in[7] & io_in[9] & io_in[11]) | (~io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & io_in[6] & io_in[7] & io_in[8] & ~io_in[9] & io_in[10] & ~io_in[11]) | (io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & ~io_in[6] & ~io_in[7] & io_in[8] & io_in[10] & ~io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[5] & ~io_in[6] & ~io_in[7] & io_in[8] & ~io_in[9] & io_in[10] & ~io_in[11]) | (io_in[0] & io_in[1] & ~io_in[2] & io_in[3] & ~io_in[4] & ~io_in[6] & ~io_in[7] & io_in[8] & io_in[9] & ~io_in[10]) | (io_in[1] & io_in[2] & io_in[4] & io_in[6] & io_in[7] & io_in[10] & io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & io_in[6] & io_in[7] & io_in[8] & io_in[10]) | (io_in[0] & io_in[1] & ~io_in[2] & io_in[4] & io_in[6] & io_in[7] & io_in[9] & ~io_in[10] & ~io_in[11]) | (io_in[1] & ~io_in[2] & io_in[5] & io_in[6] & io_in[7] & io_in[9] & io_in[11]) | (~io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & ~io_in[7] & io_in[11]) | (io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[6] & io_in[7] & io_in[9] & io_in[11]) | (io_in[0] & io_in[1] & ~io_in[5] & io_in[6] & ~io_in[7] & io_in[10] & io_in[11]) | (io_in[0] & io_in[3] & io_in[4] & io_in[6] & io_in[7] & io_in[10] & io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & io_in[3] & ~io_in[5] & ~io_in[6] & ~io_in[7] & ~io_in[8] & io_in[10]) | (~io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[6] & ~io_in[7] & ~io_in[8] & ~io_in[9]) | (io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[8] & io_in[9] & ~io_in[10]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & io_in[5] & io_in[6] & io_in[8] & io_in[10] & ~io_in[11]) | (io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[6] & io_in[8] & io_in[10] & ~io_in[11]) | (io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[5] & ~io_in[6] & io_in[7] & io_in[8] & ~io_in[10]) | (io_in[0] & io_in[1] & ~io_in[2] & io_in[3] & io_in[4] & io_in[6] & io_in[9] & io_in[11]) | (io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & io_in[6] & ~io_in[8] & ~io_in[9] & io_in[10]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[7] & ~io_in[8] & io_in[9] & io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & io_in[7] & io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & io_in[1] & io_in[2] & io_in[3] & io_in[4] & ~io_in[7] & ~io_in[8] & io_in[9] & io_in[10]) | (~io_in[0] & ~io_in[2] & io_in[3] & io_in[4] & ~io_in[6] & ~io_in[7] & io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & io_in[8] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & ~io_in[7] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (io_in[0] & io_in[1] & io_in[2] & io_in[3] & ~io_in[5] & ~io_in[7] & io_in[10] & io_in[11]) | (io_in[0] & io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[6] & io_in[7] & io_in[9] & ~io_in[10] & io_in[11]) | (~io_in[1] & io_in[2] & io_in[5] & ~io_in[6] & ~io_in[8] & io_in[9] & io_in[10]) | (io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & io_in[9] & ~io_in[10] & ~io_in[11]) | (io_in[0] & io_in[1] & io_in[3] & io_in[6] & ~io_in[8] & io_in[9] & ~io_in[10] & ~io_in[11]) | (io_in[0] & io_in[1] & io_in[2] & ~io_in[3] & io_in[4] & io_in[6] & ~io_in[7] & ~io_in[9] & io_in[10]) | (io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & io_in[4] & ~io_in[6] & ~io_in[8] & ~io_in[9] & io_in[11]) | (io_in[0] & io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & io_in[6] & ~io_in[7] & ~io_in[8] & io_in[11]) | (io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & ~io_in[6] & ~io_in[7] & io_in[8] & io_in[9] & ~io_in[10]) | (io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & io_in[7] & io_in[8] & ~io_in[10] & io_in[11]) | (~io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & io_in[8] & io_in[9] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & io_in[7] & ~io_in[8] & io_in[10]) | (~io_in[0] & ~io_in[1] & ~io_in[3] & io_in[4] & ~io_in[6] & ~io_in[7] & io_in[8] & ~io_in[9] & io_in[11]) | (~io_in[0] & ~io_in[1] & io_in[3] & io_in[5] & ~io_in[6] & io_in[7] & ~io_in[9] & io_in[10]) | (~io_in[0] & io_in[1] & io_in[2] & io_in[4] & io_in[6] & ~io_in[7] & io_in[8] & ~io_in[9] & io_in[10]) | (io_in[1] & io_in[2] & io_in[3] & io_in[4] & ~io_in[7] & io_in[8] & io_in[9] & ~io_in[10]) | (io_in[0] & io_in[2] & ~io_in[3] & io_in[4] & io_in[6] & io_in[7] & ~io_in[8] & io_in[9] & io_in[10]) | (~io_in[1] & io_in[2] & ~io_in[3] & io_in[5] & io_in[6] & io_in[9] & ~io_in[10]) | (io_in[0] & ~io_in[1] & io_in[3] & ~io_in[4] & ~io_in[6] & ~io_in[7] & io_in[8] & ~io_in[10] & io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[4] & ~io_in[6] & io_in[7] & ~io_in[8] & io_in[9] & ~io_in[10] & ~io_in[11]) | (io_in[0] & ~io_in[1] & io_in[3] & io_in[4] & ~io_in[7] & ~io_in[8] & ~io_in[9] & io_in[11]) | (io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & ~io_in[5] & io_in[6] & io_in[8] & io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & ~io_in[6] & ~io_in[7] & io_in[9] & ~io_in[10]) | (~io_in[0] & io_in[1] & io_in[2] & ~io_in[4] & ~io_in[5] & io_in[6] & io_in[7] & ~io_in[8] & ~io_in[9] & io_in[10]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & io_in[3] & ~io_in[4] & ~io_in[6] & ~io_in[7] & ~io_in[10] & ~io_in[11]) | (io_in[0] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & ~io_in[7] & io_in[10] & io_in[11]) | (~io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[6] & io_in[7] & io_in[9] & io_in[11]) | (~io_in[1] & io_in[2] & io_in[3] & io_in[5] & io_in[6] & ~io_in[9]) | (~io_in[0] & ~io_in[1] & io_in[5] & io_in[7] & io_in[9] & ~io_in[10] & io_in[11]) | (~io_in[0] & io_in[2] & ~io_in[3] & io_in[4] & io_in[6] & io_in[7] & io_in[8] & io_in[9] & io_in[10]) | (io_in[0] & ~io_in[1] & io_in[3] & ~io_in[4] & io_in[6] & io_in[7] & io_in[8] & ~io_in[10] & io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[3] & ~io_in[4] & ~io_in[6] & ~io_in[7] & ~io_in[8] & ~io_in[9] & ~io_in[10] & io_in[11]) | (~io_in[0] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & ~io_in[7] & ~io_in[8] & ~io_in[9] & io_in[10] & ~io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & io_in[6] & ~io_in[7] & ~io_in[8] & ~io_in[9] & io_in[11]) | (~io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & ~io_in[6] & ~io_in[7] & io_in[9] & io_in[10] & ~io_in[11]) | (io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & io_in[7] & io_in[8] & io_in[9] & io_in[10] & ~io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & io_in[3] & io_in[4] & io_in[6] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & io_in[3] & io_in[4] & io_in[6] & io_in[7] & ~io_in[8] & io_in[9] & io_in[10]) | (io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & io_in[4] & io_in[6] & io_in[7] & io_in[8] & io_in[9]) | (~io_in[0] & io_in[1] & io_in[2] & ~io_in[3] & io_in[4] & ~io_in[6] & io_in[7] & io_in[9] & io_in[10] & ~io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & io_in[3] & ~io_in[4] & io_in[7] & io_in[10] & io_in[11]) | (io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & ~io_in[8] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & io_in[3] & io_in[4] & ~io_in[6] & io_in[7] & ~io_in[8] & io_in[11]) | (io_in[0] & ~io_in[1] & ~io_in[3] & io_in[4] & io_in[6] & ~io_in[7] & io_in[8] & ~io_in[10] & io_in[11]) | (~io_in[0] & io_in[1] & io_in[3] & io_in[6] & io_in[7] & io_in[10] & io_in[11]) | (~io_in[0] & ~io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & ~io_in[6] & io_in[7] & io_in[8] & io_in[9] & ~io_in[10]) | (io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[5] & io_in[6] & ~io_in[7] & ~io_in[8] & io_in[9] & io_in[10]) | (io_in[0] & io_in[1] & io_in[2] & ~io_in[4] & ~io_in[5] & io_in[6] & io_in[7] & io_in[8] & io_in[9] & ~io_in[10]);

assign val[5] = (~io_in[0] & ~io_in[2] & io_in[3] & ~io_in[5] & io_in[7] & ~io_in[9] & io_in[10]) | (io_in[1] & ~io_in[2] & io_in[3] & io_in[5] & io_in[6] & io_in[7] & io_in[10]) | (~io_in[0] & io_in[1] & io_in[4] & io_in[7] & ~io_in[8] & io_in[10]) | (io_in[0] & io_in[1] & ~io_in[2] & ~io_in[4] & ~io_in[7] & ~io_in[8]) | (io_in[1] & io_in[4] & ~io_in[8] & ~io_in[9] & io_in[10]) | (~io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[10]) | (io_in[1] & ~io_in[2] & ~io_in[5] & ~io_in[6] & ~io_in[7] & io_in[8] & io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[4] & ~io_in[5] & ~io_in[7] & io_in[11]) | (~io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & io_in[6] & ~io_in[9]) | (io_in[0] & ~io_in[4] & ~io_in[5] & io_in[6] & ~io_in[7] & io_in[8] & io_in[10]) | (~io_in[1] & ~io_in[2] & io_in[3] & ~io_in[5] & io_in[8] & ~io_in[9] & io_in[10]) | (~io_in[0] & ~io_in[5] & io_in[6] & ~io_in[7] & ~io_in[8] & io_in[9] & ~io_in[10] & io_in[11]) | (io_in[1] & ~io_in[3] & io_in[4] & ~io_in[5] & io_in[7] & io_in[11]) | (io_in[0] & io_in[2] & ~io_in[4] & ~io_in[5] & io_in[6] & ~io_in[7] & io_in[11]) | (~io_in[1] & io_in[2] & ~io_in[3] & ~io_in[8] & ~io_in[9] & io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[3] & io_in[6] & ~io_in[8] & io_in[10]) | (io_in[0] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[9] & ~io_in[11]) | (io_in[2] & ~io_in[5] & io_in[6] & ~io_in[7] & ~io_in[8] & io_in[9]) | (io_in[2] & ~io_in[3] & io_in[5] & io_in[6] & io_in[7] & ~io_in[11]) | (~io_in[0] & io_in[1] & io_in[2] & io_in[4] & ~io_in[9] & ~io_in[11]) | (~io_in[0] & io_in[1] & io_in[2] & ~io_in[4] & ~io_in[5] & io_in[8] & io_in[11]) | (io_in[2] & ~io_in[4] & ~io_in[5] & io_in[6] & io_in[9] & io_in[11]) | (~io_in[1] & ~io_in[2] & io_in[5] & ~io_in[8] & io_in[9]) | (~io_in[1] & io_in[2] & io_in[3] & io_in[6] & io_in[10]) | (~io_in[1] & ~io_in[2] & io_in[5] & ~io_in[6] & io_in[7] & io_in[10]) | (io_in[0] & ~io_in[1] & ~io_in[2] & io_in[3] & ~io_in[10] & ~io_in[11]) | (io_in[1] & ~io_in[2] & io_in[4] & io_in[6] & io_in[9] & ~io_in[10]) | (io_in[0] & ~io_in[1] & ~io_in[2] & io_in[3] & io_in[7] & ~io_in[10]) | (~io_in[0] & io_in[3] & ~io_in[5] & io_in[6] & io_in[7] & io_in[10]) | (~io_in[1] & io_in[2] & io_in[4] & io_in[7] & io_in[8] & ~io_in[9]) | (~io_in[0] & ~io_in[1] & ~io_in[3] & io_in[4] & ~io_in[10] & io_in[11]) | (io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[6] & ~io_in[7]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & io_in[5] & ~io_in[8] & io_in[10]) | (io_in[0] & ~io_in[3] & io_in[5] & ~io_in[6] & ~io_in[7] & io_in[10]) | (io_in[0] & io_in[2] & ~io_in[5] & ~io_in[6] & io_in[7] & ~io_in[8] & io_in[10]) | (io_in[0] & ~io_in[2] & io_in[6] & io_in[7] & io_in[8] & ~io_in[10]) | (io_in[0] & io_in[2] & ~io_in[5] & io_in[6] & io_in[7] & ~io_in[8] & ~io_in[9]) | (io_in[0] & io_in[1] & ~io_in[5] & io_in[10] & io_in[11]) | (io_in[0] & ~io_in[2] & io_in[3] & io_in[4] & ~io_in[9] & ~io_in[10]) | (~io_in[1] & io_in[3] & io_in[4] & io_in[6] & ~io_in[9] & ~io_in[11]) | (~io_in[1] & io_in[3] & ~io_in[5] & io_in[6] & ~io_in[9] & io_in[10]) | (~io_in[0] & io_in[1] & io_in[2] & ~io_in[6] & io_in[7] & ~io_in[9] & ~io_in[11]) | (~io_in[0] & ~io_in[1] & io_in[4] & ~io_in[6] & ~io_in[7] & ~io_in[9]) | (io_in[0] & io_in[1] & io_in[4] & io_in[7] & ~io_in[9] & ~io_in[10]) | (~io_in[0] & ~io_in[2] & io_in[5] & ~io_in[7] & io_in[8] & ~io_in[10]) | (~io_in[0] & ~io_in[3] & io_in[5] & io_in[6] & io_in[7] & ~io_in[8]) | (~io_in[0] & ~io_in[2] & io_in[5] & io_in[6] & io_in[7] & ~io_in[9]) | (io_in[0] & ~io_in[1] & ~io_in[3] & ~io_in[4] & io_in[7] & ~io_in[8] & io_in[9]) | (io_in[1] & io_in[2] & io_in[4] & ~io_in[6] & ~io_in[7] & ~io_in[9]) | (~io_in[1] & io_in[3] & ~io_in[5] & io_in[6] & io_in[7] & io_in[8] & io_in[9]) | (io_in[0] & io_in[3] & ~io_in[5] & io_in[10] & io_in[11]) | (io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[6] & ~io_in[7] & ~io_in[9] & ~io_in[11]) | (io_in[1] & ~io_in[2] & io_in[3] & io_in[7] & io_in[8] & io_in[9] & ~io_in[11]) | (io_in[0] & ~io_in[2] & io_in[3] & io_in[6] & ~io_in[7] & ~io_in[11]) | (~io_in[1] & io_in[3] & io_in[6] & ~io_in[7] & ~io_in[8] & ~io_in[9]) | (io_in[1] & ~io_in[2] & ~io_in[4] & io_in[6] & io_in[8] & ~io_in[9] & ~io_in[11]) | (~io_in[0] & io_in[2] & ~io_in[3] & ~io_in[4] & io_in[6] & io_in[7] & io_in[9] & ~io_in[11]) | (~io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & io_in[6] & io_in[7] & ~io_in[11]) | (~io_in[0] & io_in[2] & ~io_in[5] & io_in[7] & ~io_in[8] & io_in[11]) | (~io_in[0] & ~io_in[1] & io_in[2] & io_in[6] & ~io_in[7] & io_in[9]) | (~io_in[1] & io_in[2] & ~io_in[3] & ~io_in[5] & ~io_in[7] & ~io_in[10] & io_in[11]) | (~io_in[1] & ~io_in[3] & ~io_in[6] & ~io_in[7] & ~io_in[8] & ~io_in[9] & ~io_in[10] & io_in[11]) | (~io_in[0] & io_in[2] & ~io_in[6] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (io_in[1] & ~io_in[2] & ~io_in[5] & io_in[7] & io_in[8] & io_in[9] & ~io_in[11]) | (~io_in[1] & ~io_in[3] & ~io_in[4] & io_in[5] & io_in[6] & io_in[7] & ~io_in[11]) | (~io_in[0] & ~io_in[2] & ~io_in[3] & io_in[4] & io_in[7] & ~io_in[10]) | (~io_in[1] & ~io_in[2] & io_in[5] & ~io_in[6] & ~io_in[8]) | (~io_in[0] & io_in[3] & ~io_in[4] & ~io_in[5] & io_in[8] & io_in[11]) | (~io_in[1] & io_in[2] & ~io_in[4] & ~io_in[5] & ~io_in[8] & io_in[10]) | (~io_in[1] & io_in[3] & io_in[4] & io_in[8] & ~io_in[9] & ~io_in[11]) | (~io_in[1] & io_in[2] & ~io_in[4] & ~io_in[5] & ~io_in[7] & io_in[8] & io_in[11]) | (io_in[0] & ~io_in[1] & io_in[4] & ~io_in[5] & io_in[7] & io_in[10]) | (~io_in[0] & ~io_in[4] & io_in[5] & ~io_in[6] & io_in[10] & io_in[11]) | (io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[6] & io_in[11]) | (io_in[0] & io_in[1] & io_in[4] & ~io_in[6] & ~io_in[7] & io_in[10]) | (~io_in[0] & io_in[2] & ~io_in[4] & ~io_in[5] & io_in[6] & io_in[7] & io_in[10]) | (~io_in[0] & io_in[1] & io_in[2] & ~io_in[5] & ~io_in[6] & ~io_in[7] & io_in[8]) | (io_in[0] & io_in[2] & io_in[3] & io_in[4] & io_in[9] & io_in[10]) | (~io_in[0] & ~io_in[2] & ~io_in[4] & io_in[7] & ~io_in[8] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[1] & io_in[2] & ~io_in[3] & ~io_in[8] & io_in[10]) | (io_in[0] & io_in[2] & io_in[6] & ~io_in[8] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & ~io_in[2] & ~io_in[3] & io_in[4] & io_in[6] & ~io_in[7] & ~io_in[9]) | (io_in[0] & ~io_in[2] & ~io_in[3] & ~io_in[6] & io_in[8] & io_in[10]) | (~io_in[0] & io_in[2] & io_in[5] & ~io_in[7] & ~io_in[8]) | (~io_in[1] & ~io_in[2] & io_in[5] & ~io_in[7] & io_in[11]) | (io_in[0] & io_in[1] & ~io_in[3] & io_in[4] & ~io_in[8] & ~io_in[9]) | (io_in[1] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & ~io_in[8] & io_in[9]) | (~io_in[0] & ~io_in[1] & io_in[2] & ~io_in[4] & ~io_in[5] & io_in[7] & io_in[8] & io_in[9]) | (io_in[1] & ~io_in[2] & ~io_in[3] & io_in[6] & io_in[7] & ~io_in[9] & ~io_in[10]) | (io_in[1] & ~io_in[3] & ~io_in[5] & ~io_in[6] & io_in[7] & io_in[9] & ~io_in[10] & ~io_in[11]) | (io_in[0] & ~io_in[1] & ~io_in[2] & io_in[6] & io_in[8] & ~io_in[10]) | (io_in[0] & io_in[1] & ~io_in[2] & io_in[3] & ~io_in[6] & ~io_in[8]) | (io_in[2] & ~io_in[3] & io_in[4] & io_in[6] & ~io_in[7] & io_in[9] & ~io_in[11]) | (io_in[0] & io_in[1] & io_in[4] & io_in[7] & io_in[8] & io_in[9]) | (~io_in[1] & ~io_in[4] & ~io_in[5] & io_in[6] & ~io_in[7] & ~io_in[8] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (io_in[0] & ~io_in[2] & ~io_in[3] & ~io_in[5] & io_in[7] & io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & io_in[7] & ~io_in[8] & ~io_in[9]) | (~io_in[1] & io_in[3] & ~io_in[7] & io_in[10] & io_in[11]) | (~io_in[1] & ~io_in[2] & io_in[3] & ~io_in[4] & ~io_in[6] & ~io_in[7] & io_in[9]) | (~io_in[1] & ~io_in[2] & io_in[4] & ~io_in[7] & ~io_in[9]) | (io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & io_in[8] & io_in[10]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & io_in[5] & ~io_in[7] & io_in[8]) | (io_in[0] & ~io_in[2] & ~io_in[3] & ~io_in[4] & io_in[8] & io_in[10] & ~io_in[11]) | (io_in[0] & io_in[3] & ~io_in[4] & io_in[6] & io_in[8] & ~io_in[11]) | (io_in[0] & io_in[1] & io_in[2] & io_in[3] & io_in[7] & io_in[8]) | (io_in[2] & ~io_in[5] & io_in[6] & ~io_in[7] & io_in[9] & io_in[10] & ~io_in[11]) | (~io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[7] & io_in[8] & io_in[10]) | (~io_in[0] & ~io_in[1] & io_in[4] & ~io_in[5] & ~io_in[6] & ~io_in[7] & io_in[8]) | (~io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & ~io_in[5] & io_in[6] & io_in[9]) | (io_in[0] & ~io_in[1] & io_in[8] & ~io_in[9] & io_in[10]) | (io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & io_in[6] & ~io_in[9] & io_in[11]) | (io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[5] & ~io_in[6] & io_in[7] & io_in[9]) | (io_in[1] & io_in[2] & io_in[3] & ~io_in[6] & io_in[9] & io_in[10]) | (io_in[0] & ~io_in[2] & ~io_in[3] & ~io_in[5] & ~io_in[9] & io_in[10]) | (~io_in[2] & io_in[4] & io_in[6] & io_in[10] & io_in[11]) | (~io_in[1] & io_in[2] & ~io_in[3] & io_in[4] & io_in[9] & io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[2] & io_in[3] & ~io_in[4] & ~io_in[7] & ~io_in[10]) | (~io_in[0] & io_in[2] & ~io_in[5] & io_in[6] & ~io_in[8] & io_in[10]) | (io_in[1] & io_in[3] & ~io_in[4] & io_in[7] & io_in[8] & io_in[10]) | (io_in[0] & ~io_in[1] & io_in[2] & ~io_in[4] & io_in[7] & ~io_in[8] & ~io_in[9]) | (io_in[1] & io_in[3] & ~io_in[7] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[3] & io_in[5] & io_in[6] & io_in[7] & ~io_in[11]) | (~io_in[1] & ~io_in[3] & io_in[4] & ~io_in[8] & io_in[9] & io_in[10]) | (~io_in[1] & ~io_in[2] & io_in[4] & io_in[10] & io_in[11]) | (io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & ~io_in[8] & ~io_in[10]) | (io_in[0] & io_in[1] & io_in[2] & io_in[4] & io_in[8] & io_in[11]) | (~io_in[0] & io_in[3] & ~io_in[4] & ~io_in[5] & io_in[9] & io_in[11]) | (io_in[1] & ~io_in[2] & io_in[4] & io_in[7] & ~io_in[10] & io_in[11]) | (io_in[0] & io_in[1] & io_in[2] & io_in[3] & ~io_in[5] & ~io_in[7] & io_in[9]) | (io_in[0] & ~io_in[4] & ~io_in[5] & ~io_in[6] & io_in[9] & ~io_in[10] & ~io_in[11]) | (io_in[0] & ~io_in[1] & ~io_in[3] & ~io_in[4] & ~io_in[6] & ~io_in[8]) | (~io_in[1] & ~io_in[2] & io_in[4] & ~io_in[9] & ~io_in[11]) | (io_in[0] & io_in[2] & ~io_in[6] & io_in[7] & io_in[8] & ~io_in[10]) | (io_in[1] & ~io_in[2] & ~io_in[5] & ~io_in[7] & io_in[9] & io_in[11]) | (io_in[0] & ~io_in[2] & ~io_in[3] & ~io_in[6] & ~io_in[7] & io_in[11]) | (io_in[1] & ~io_in[2] & ~io_in[4] & ~io_in[5] & io_in[6] & io_in[9] & io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[2] & io_in[5] & io_in[6] & ~io_in[7]) | (io_in[0] & io_in[4] & io_in[7] & io_in[8] & io_in[11]) | (~io_in[0] & io_in[3] & ~io_in[5] & io_in[6] & ~io_in[7] & ~io_in[8] & ~io_in[10]) | (io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[7] & io_in[10] & io_in[11]) | (io_in[0] & ~io_in[4] & ~io_in[6] & io_in[7] & ~io_in[8] & ~io_in[9] & io_in[11]) | (~io_in[0] & ~io_in[1] & io_in[3] & ~io_in[4] & io_in[6] & io_in[11]) | (~io_in[2] & ~io_in[5] & io_in[6] & ~io_in[7] & io_in[8] & io_in[9] & io_in[10] & io_in[11]) | (io_in[0] & ~io_in[2] & io_in[3] & ~io_in[5] & ~io_in[8] & ~io_in[9] & ~io_in[10]) | (~io_in[1] & ~io_in[2] & io_in[4] & ~io_in[7] & ~io_in[8] & ~io_in[11]) | (io_in[0] & io_in[1] & io_in[2] & io_in[3] & ~io_in[5] & ~io_in[6] & ~io_in[11]) | (~io_in[0] & io_in[1] & io_in[3] & io_in[4] & io_in[8] & io_in[9] & ~io_in[11]) | (io_in[0] & ~io_in[1] & ~io_in[3] & ~io_in[6] & io_in[9] & ~io_in[10]) | (io_in[1] & io_in[3] & ~io_in[4] & ~io_in[6] & ~io_in[8] & ~io_in[10]) | (io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & io_in[11]) | (~io_in[1] & ~io_in[2] & io_in[5] & ~io_in[6] & io_in[9]) | (~io_in[0] & ~io_in[3] & io_in[4] & io_in[8] & ~io_in[9] & ~io_in[10]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[6] & io_in[7] & ~io_in[11]) | (io_in[2] & ~io_in[4] & io_in[6] & ~io_in[7] & io_in[8] & ~io_in[9] & ~io_in[10]) | (io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[5] & io_in[6] & io_in[9] & ~io_in[10]) | (~io_in[0] & io_in[2] & ~io_in[3] & io_in[4] & io_in[8] & ~io_in[10]) | (io_in[2] & ~io_in[3] & io_in[5] & ~io_in[8] & ~io_in[9] & ~io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & ~io_in[7] & io_in[10]) | (~io_in[1] & ~io_in[3] & io_in[5] & ~io_in[6] & io_in[7] & io_in[8] & io_in[9]) | (io_in[0] & io_in[1] & ~io_in[4] & ~io_in[5] & ~io_in[7] & io_in[9] & io_in[11]) | (~io_in[0] & io_in[1] & io_in[3] & ~io_in[4] & ~io_in[6] & ~io_in[7] & io_in[8]) | (~io_in[1] & ~io_in[2] & io_in[3] & io_in[6] & ~io_in[8] & ~io_in[10] & ~io_in[11]) | (io_in[0] & ~io_in[5] & io_in[6] & io_in[7] & ~io_in[8] & ~io_in[9] & io_in[11]) | (io_in[0] & ~io_in[2] & ~io_in[5] & ~io_in[6] & io_in[7] & io_in[9]) | (io_in[0] & ~io_in[2] & io_in[3] & io_in[6] & io_in[8] & io_in[9]) | (io_in[1] & io_in[2] & ~io_in[5] & ~io_in[6] & ~io_in[7] & io_in[8] & io_in[10]) | (~io_in[0] & io_in[4] & ~io_in[6] & io_in[7] & ~io_in[8] & ~io_in[9] & ~io_in[10]) | (~io_in[0] & ~io_in[1] & io_in[3] & ~io_in[4] & io_in[7] & ~io_in[8] & io_in[10]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[4] & ~io_in[5] & ~io_in[7] & io_in[10]) | (io_in[1] & io_in[2] & ~io_in[3] & ~io_in[5] & ~io_in[6] & io_in[8] & ~io_in[9]) | (io_in[2] & ~io_in[6] & ~io_in[7] & io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & ~io_in[2] & ~io_in[5] & ~io_in[7] & ~io_in[8] & ~io_in[9]) | (io_in[1] & io_in[2] & ~io_in[3] & io_in[4] & ~io_in[7] & io_in[10]) | (~io_in[1] & ~io_in[2] & io_in[5] & io_in[9] & io_in[11]) | (~io_in[1] & ~io_in[2] & io_in[4] & ~io_in[6] & ~io_in[10] & ~io_in[11]) | (~io_in[1] & io_in[2] & io_in[3] & io_in[4] & ~io_in[6] & io_in[7] & ~io_in[8] & io_in[9]) | (~io_in[1] & io_in[2] & io_in[3] & io_in[4] & io_in[9] & io_in[11]) | (io_in[0] & ~io_in[6] & io_in[7] & ~io_in[8] & io_in[9] & ~io_in[11]);

assign val[6] = (~io_in[0] & ~io_in[2] & ~io_in[3] & io_in[4] & io_in[5]) | (~io_in[1] & io_in[2] & io_in[3] & io_in[6] & ~io_in[8] & ~io_in[9]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[5] & ~io_in[6] & io_in[8]) | (io_in[0] & io_in[2] & io_in[3] & io_in[7] & ~io_in[8] & io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & io_in[4] & ~io_in[5] & ~io_in[6] & io_in[8] & io_in[9]) | (~io_in[1] & io_in[2] & ~io_in[4] & ~io_in[7] & io_in[8] & ~io_in[9] & io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[7] & ~io_in[9]) | (io_in[1] & io_in[2] & io_in[4] & ~io_in[6] & ~io_in[8] & ~io_in[9]) | (io_in[0] & io_in[1] & ~io_in[2] & io_in[3] & io_in[4] & io_in[6] & ~io_in[8] & ~io_in[11]) | (~io_in[1] & ~io_in[2] & ~io_in[5] & ~io_in[7] & io_in[8] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (io_in[0] & io_in[2] & io_in[3] & ~io_in[4] & ~io_in[6] & io_in[11]) | (io_in[1] & io_in[2] & ~io_in[3] & io_in[4] & ~io_in[7] & ~io_in[9] & ~io_in[10]) | (io_in[0] & io_in[2] & ~io_in[6] & io_in[7] & io_in[10] & io_in[11]) | (~io_in[1] & ~io_in[2] & io_in[3] & io_in[4] & ~io_in[7] & io_in[10] & io_in[11]) | (~io_in[0] & io_in[3] & ~io_in[7] & ~io_in[8] & io_in[9] & io_in[10]) | (io_in[2] & io_in[3] & io_in[4] & ~io_in[8] & io_in[9] & io_in[10]) | (io_in[0] & ~io_in[1] & ~io_in[4] & ~io_in[6] & io_in[8] & io_in[11]) | (io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & ~io_in[6] & io_in[9] & io_in[11]) | (io_in[1] & ~io_in[2] & io_in[3] & io_in[4] & ~io_in[7] & ~io_in[9] & io_in[10]) | (io_in[2] & io_in[4] & io_in[6] & ~io_in[7] & ~io_in[8] & io_in[9]) | (io_in[0] & io_in[1] & ~io_in[3] & ~io_in[4] & io_in[7] & ~io_in[8] & ~io_in[9] & ~io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & io_in[4] & io_in[7] & ~io_in[8] & ~io_in[9]) | (io_in[0] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & io_in[9] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & io_in[3] & io_in[7] & ~io_in[8] & ~io_in[10]) | (io_in[0] & io_in[2] & io_in[3] & ~io_in[6] & ~io_in[7] & io_in[8] & ~io_in[10]) | (io_in[0] & ~io_in[1] & ~io_in[4] & io_in[7] & io_in[8] & ~io_in[9]) | (io_in[0] & ~io_in[1] & io_in[3] & io_in[4] & io_in[8] & io_in[9] & ~io_in[11]) | (~io_in[0] & ~io_in[2] & io_in[5] & io_in[6] & io_in[8] & ~io_in[10]) | (io_in[2] & ~io_in[3] & ~io_in[4] & io_in[7] & ~io_in[8] & io_in[10]) | (~io_in[1] & ~io_in[3] & ~io_in[4] & io_in[7] & ~io_in[8] & io_in[9] & ~io_in[10]) | (io_in[1] & ~io_in[2] & io_in[4] & io_in[6] & io_in[9] & ~io_in[10]) | (io_in[0] & ~io_in[1] & ~io_in[3] & ~io_in[5] & ~io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & io_in[2] & ~io_in[3] & io_in[4] & ~io_in[6] & ~io_in[7] & ~io_in[9]) | (~io_in[0] & io_in[2] & ~io_in[4] & ~io_in[5] & io_in[6] & io_in[7] & ~io_in[8] & ~io_in[9]) | (~io_in[1] & ~io_in[2] & io_in[3] & ~io_in[4] & ~io_in[6] & io_in[7] & ~io_in[10]) | (io_in[0] & io_in[1] & ~io_in[2] & io_in[8] & io_in[9] & io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[2] & io_in[4] & ~io_in[5] & ~io_in[6] & io_in[7] & io_in[8] & io_in[9]) | (io_in[2] & io_in[3] & ~io_in[4] & io_in[6] & ~io_in[7] & io_in[8] & io_in[10] & ~io_in[11]) | (io_in[0] & ~io_in[2] & ~io_in[4] & io_in[6] & ~io_in[7] & ~io_in[10] & io_in[11]) | (io_in[0] & ~io_in[2] & io_in[4] & ~io_in[6] & io_in[7] & io_in[8] & ~io_in[9]) | (io_in[0] & ~io_in[1] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[7] & io_in[9]) | (io_in[1] & io_in[2] & ~io_in[4] & ~io_in[7] & io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & ~io_in[2] & ~io_in[4] & ~io_in[6] & ~io_in[7] & io_in[8] & io_in[10]) | (io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[7] & ~io_in[8]) | (io_in[0] & ~io_in[2] & io_in[3] & io_in[4] & io_in[6] & ~io_in[7] & io_in[8] & io_in[9]) | (io_in[1] & ~io_in[2] & ~io_in[4] & ~io_in[5] & ~io_in[6] & ~io_in[7] & io_in[11]) | (io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & io_in[7] & io_in[10] & io_in[11]) | (io_in[0] & ~io_in[1] & ~io_in[3] & ~io_in[6] & ~io_in[7] & io_in[8] & io_in[11]) | (io_in[1] & io_in[3] & io_in[4] & io_in[8] & ~io_in[10] & io_in[11]) | (~io_in[0] & ~io_in[2] & io_in[3] & io_in[4] & io_in[6] & ~io_in[9] & io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[3] & io_in[4] & io_in[7] & ~io_in[10]) | (io_in[0] & ~io_in[1] & ~io_in[3] & io_in[4] & io_in[6] & ~io_in[7] & ~io_in[11]) | (io_in[0] & io_in[2] & io_in[4] & ~io_in[7] & ~io_in[8] & io_in[10]) | (io_in[1] & io_in[4] & ~io_in[7] & ~io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & io_in[5] & io_in[7] & io_in[11]) | (~io_in[1] & io_in[5] & ~io_in[7] & io_in[8] & io_in[9] & ~io_in[11]) | (io_in[0] & io_in[1] & io_in[2] & io_in[3] & ~io_in[8] & io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & io_in[8] & io_in[10] & ~io_in[11]) | (io_in[0] & io_in[1] & ~io_in[3] & ~io_in[5] & io_in[6] & io_in[7] & io_in[8] & ~io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & io_in[4] & ~io_in[7] & ~io_in[9] & ~io_in[10]) | (io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[6] & ~io_in[7] & io_in[8] & io_in[9] & ~io_in[11]) | (io_in[1] & ~io_in[2] & io_in[3] & io_in[5] & io_in[6] & io_in[10]) | (io_in[0] & io_in[2] & ~io_in[6] & ~io_in[7] & io_in[9] & ~io_in[11]) | (io_in[0] & io_in[2] & ~io_in[3] & io_in[4] & ~io_in[7] & ~io_in[9] & ~io_in[11]) | (io_in[1] & ~io_in[4] & ~io_in[5] & io_in[6] & ~io_in[8] & ~io_in[9] & io_in[11]) | (io_in[1] & ~io_in[2] & io_in[3] & ~io_in[4] & io_in[8] & ~io_in[10] & ~io_in[11]) | (~io_in[2] & ~io_in[3] & ~io_in[5] & ~io_in[6] & io_in[7] & io_in[9] & io_in[10] & ~io_in[11]) | (~io_in[2] & ~io_in[4] & ~io_in[6] & io_in[7] & ~io_in[8] & ~io_in[9] & ~io_in[10] & io_in[11]) | (~io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & io_in[6] & ~io_in[9] & ~io_in[10]) | (~io_in[0] & io_in[2] & ~io_in[5] & io_in[6] & ~io_in[8] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (io_in[0] & ~io_in[1] & ~io_in[3] & io_in[6] & io_in[7] & ~io_in[9] & io_in[11]) | (~io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & io_in[7] & io_in[9] & ~io_in[10]) | (~io_in[0] & ~io_in[1] & io_in[3] & io_in[4] & ~io_in[6] & ~io_in[8] & io_in[9]) | (~io_in[0] & io_in[1] & io_in[2] & ~io_in[6] & io_in[7] & io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & io_in[7] & ~io_in[11]) | (~io_in[1] & ~io_in[2] & ~io_in[3] & io_in[5] & io_in[7] & ~io_in[8] & ~io_in[11]) | (io_in[1] & io_in[2] & io_in[4] & io_in[6] & ~io_in[7] & io_in[9] & io_in[11]) | (io_in[2] & io_in[3] & ~io_in[5] & ~io_in[6] & io_in[7] & ~io_in[9] & io_in[10]) | (~io_in[0] & io_in[1] & ~io_in[3] & ~io_in[6] & ~io_in[7] & io_in[9] & io_in[11]) | (~io_in[1] & io_in[3] & ~io_in[4] & ~io_in[6] & ~io_in[7] & io_in[8] & io_in[9]) | (io_in[1] & ~io_in[3] & ~io_in[5] & ~io_in[6] & ~io_in[7] & ~io_in[10] & io_in[11]) | (io_in[0] & ~io_in[2] & ~io_in[3] & io_in[6] & ~io_in[8] & io_in[11]) | (~io_in[1] & io_in[2] & ~io_in[6] & io_in[8] & ~io_in[9] & io_in[10]) | (~io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[5] & io_in[7] & io_in[9] & io_in[10] & ~io_in[11]) | (~io_in[1] & ~io_in[2] & ~io_in[5] & io_in[7] & io_in[8] & ~io_in[9] & ~io_in[10] & io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[4] & ~io_in[5] & ~io_in[6] & io_in[7] & io_in[9] & ~io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[4] & ~io_in[5] & ~io_in[7] & ~io_in[8]) | (~io_in[0] & ~io_in[1] & io_in[2] & ~io_in[4] & io_in[6] & io_in[7] & io_in[10]) | (~io_in[0] & ~io_in[2] & io_in[6] & io_in[7] & io_in[8] & io_in[10] & ~io_in[11]) | (~io_in[1] & io_in[5] & ~io_in[6] & io_in[9] & ~io_in[11]) | (~io_in[0] & io_in[1] & io_in[2] & io_in[6] & ~io_in[7] & ~io_in[10] & ~io_in[11]) | (~io_in[1] & ~io_in[3] & ~io_in[7] & io_in[8] & ~io_in[9] & ~io_in[10] & io_in[11]) | (~io_in[1] & io_in[3] & io_in[4] & io_in[6] & io_in[7] & io_in[8] & ~io_in[11]) | (~io_in[1] & io_in[2] & io_in[3] & ~io_in[6] & io_in[7] & ~io_in[8] & ~io_in[11]) | (~io_in[2] & ~io_in[4] & io_in[6] & ~io_in[7] & io_in[8] & ~io_in[9] & ~io_in[11]) | (~io_in[2] & io_in[3] & ~io_in[4] & io_in[6] & io_in[7] & io_in[8]) | (io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & io_in[4] & ~io_in[5] & ~io_in[7] & io_in[8]) | (~io_in[0] & io_in[1] & ~io_in[3] & io_in[6] & io_in[7] & ~io_in[8] & ~io_in[10]) | (~io_in[0] & io_in[2] & io_in[3] & io_in[4] & io_in[6] & ~io_in[7] & io_in[10]) | (~io_in[1] & io_in[3] & io_in[4] & ~io_in[7] & ~io_in[8] & ~io_in[9] & io_in[11]) | (io_in[2] & ~io_in[4] & ~io_in[5] & ~io_in[6] & io_in[7] & io_in[8] & ~io_in[9]) | (~io_in[0] & ~io_in[2] & ~io_in[3] & io_in[4] & ~io_in[6] & io_in[8] & ~io_in[11]) | (~io_in[0] & ~io_in[1] & io_in[2] & io_in[8] & ~io_in[9] & io_in[10]) | (io_in[1] & io_in[2] & ~io_in[3] & io_in[4] & io_in[7] & ~io_in[10] & ~io_in[11]) | (io_in[0] & io_in[2] & io_in[6] & io_in[7] & ~io_in[8] & io_in[9] & io_in[10]) | (io_in[0] & ~io_in[1] & ~io_in[5] & io_in[6] & ~io_in[8] & ~io_in[9] & io_in[10]) | (~io_in[0] & ~io_in[1] & io_in[4] & io_in[5]) | (~io_in[0] & io_in[3] & ~io_in[4] & ~io_in[5] & io_in[7] & io_in[9] & ~io_in[10] & ~io_in[11]) | (io_in[0] & io_in[1] & io_in[3] & ~io_in[5] & ~io_in[6] & io_in[7] & io_in[11]) | (io_in[2] & io_in[3] & ~io_in[6] & ~io_in[8] & io_in[9] & io_in[10]) | (~io_in[1] & ~io_in[3] & io_in[6] & ~io_in[7] & io_in[8] & ~io_in[9] & ~io_in[10]) | (~io_in[0] & io_in[1] & io_in[2] & io_in[4] & io_in[6] & ~io_in[7] & ~io_in[11]) | (io_in[1] & io_in[5] & ~io_in[6] & io_in[7] & ~io_in[9] & io_in[11]) | (io_in[1] & io_in[2] & io_in[6] & io_in[7] & ~io_in[8] & ~io_in[10] & ~io_in[11]) | (io_in[0] & io_in[2] & io_in[6] & ~io_in[7] & ~io_in[8] & ~io_in[9] & io_in[10]) | (io_in[1] & io_in[2] & ~io_in[3] & io_in[4] & ~io_in[7] & io_in[11]) | (io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & io_in[6] & io_in[8] & ~io_in[10]) | (~io_in[1] & io_in[3] & ~io_in[4] & ~io_in[8] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[2] & ~io_in[3] & io_in[5] & ~io_in[7] & io_in[9] & io_in[11]) | (io_in[1] & ~io_in[2] & ~io_in[4] & ~io_in[5] & ~io_in[8] & io_in[9] & io_in[10]) | (io_in[1] & ~io_in[2] & io_in[6] & io_in[7] & io_in[9] & ~io_in[10] & ~io_in[11]) | (io_in[0] & ~io_in[2] & io_in[4] & ~io_in[8] & io_in[9] & io_in[11]) | (~io_in[0] & io_in[2] & io_in[3] & io_in[4] & ~io_in[6] & io_in[8] & ~io_in[11]) | (~io_in[0] & ~io_in[1] & io_in[3] & ~io_in[5] & io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & io_in[3] & io_in[4] & io_in[6] & io_in[9] & ~io_in[10]) | (io_in[0] & ~io_in[3] & ~io_in[4] & ~io_in[5] & ~io_in[6] & io_in[7] & io_in[10]) | (io_in[0] & ~io_in[3] & ~io_in[5] & ~io_in[7] & io_in[8] & ~io_in[10] & io_in[11]) | (~io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[10] & ~io_in[11]) | (io_in[0] & ~io_in[2] & io_in[6] & ~io_in[8] & io_in[9] & io_in[11]) | (io_in[0] & ~io_in[1] & ~io_in[4] & ~io_in[5] & io_in[6] & ~io_in[8] & io_in[10]) | (~io_in[0] & ~io_in[1] & io_in[2] & io_in[6] & io_in[7] & io_in[10] & ~io_in[11]) | (io_in[0] & io_in[2] & io_in[3] & io_in[4] & io_in[7] & io_in[9] & ~io_in[11]) | (~io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & ~io_in[7] & io_in[9] & ~io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[4] & io_in[6] & io_in[7] & io_in[8]) | (io_in[0] & ~io_in[1] & ~io_in[3] & ~io_in[5] & ~io_in[6] & io_in[7] & io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & io_in[3] & ~io_in[5] & io_in[6] & ~io_in[9]) | (io_in[0] & ~io_in[1] & ~io_in[5] & io_in[7] & ~io_in[8] & ~io_in[9] & io_in[10]) | (~io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & io_in[6] & ~io_in[8] & io_in[9]) | (io_in[0] & io_in[1] & ~io_in[3] & io_in[4] & ~io_in[5] & ~io_in[6] & ~io_in[7]) | (io_in[0] & io_in[3] & io_in[4] & io_in[7] & io_in[9] & io_in[10] & ~io_in[11]) | (io_in[1] & ~io_in[2] & io_in[3] & ~io_in[4] & ~io_in[6] & io_in[7] & ~io_in[8] & ~io_in[9]) | (~io_in[0] & io_in[2] & ~io_in[3] & ~io_in[5] & ~io_in[7] & ~io_in[10] & io_in[11]) | (io_in[0] & io_in[1] & io_in[5] & io_in[6] & io_in[8] & io_in[11]) | (~io_in[0] & io_in[2] & ~io_in[4] & ~io_in[6] & ~io_in[9] & io_in[10]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[5] & ~io_in[6] & io_in[7] & io_in[9]) | (~io_in[0] & io_in[2] & io_in[6] & ~io_in[8] & io_in[9] & io_in[11]) | (~io_in[1] & ~io_in[4] & ~io_in[5] & ~io_in[6] & io_in[8] & io_in[9] & io_in[10] & io_in[11]) | (~io_in[0] & io_in[2] & ~io_in[3] & ~io_in[6] & ~io_in[8] & ~io_in[9] & io_in[11]) | (io_in[1] & io_in[2] & io_in[3] & io_in[7] & ~io_in[9] & io_in[11]) | (~io_in[0] & io_in[3] & io_in[4] & ~io_in[6] & io_in[7] & io_in[8] & io_in[11]) | (~io_in[1] & io_in[5] & ~io_in[7] & ~io_in[9] & io_in[11]) | (io_in[0] & io_in[1] & ~io_in[2] & io_in[5] & io_in[6] & io_in[10]) | (~io_in[1] & io_in[2] & ~io_in[4] & ~io_in[5] & ~io_in[6] & io_in[7] & ~io_in[9]) | (io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & io_in[7] & ~io_in[8]) | (~io_in[1] & ~io_in[3] & ~io_in[4] & io_in[5] & ~io_in[6] & io_in[7] & io_in[10]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[7] & ~io_in[8] & io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[3] & ~io_in[5] & ~io_in[6] & ~io_in[8] & io_in[9] & io_in[10]) | (~io_in[0] & ~io_in[1] & io_in[5] & io_in[6] & ~io_in[7] & io_in[9]) | (~io_in[0] & ~io_in[2] & ~io_in[3] & io_in[4] & ~io_in[6] & ~io_in[9] & ~io_in[11]) | (~io_in[0] & io_in[2] & io_in[6] & ~io_in[7] & ~io_in[8] & io_in[9]) | (~io_in[2] & io_in[4] & io_in[6] & io_in[7] & ~io_in[9] & io_in[11]) | (~io_in[1] & io_in[2] & io_in[7] & ~io_in[9] & io_in[10]) | (~io_in[2] & io_in[3] & io_in[4] & io_in[6] & io_in[8] & io_in[9] & ~io_in[11]) | (~io_in[0] & ~io_in[2] & ~io_in[4] & io_in[7] & io_in[8] & io_in[10] & ~io_in[11]) | (io_in[0] & ~io_in[1] & io_in[2] & io_in[7] & ~io_in[8] & io_in[10]) | (~io_in[0] & ~io_in[3] & io_in[5] & io_in[6] & io_in[8] & ~io_in[11]) | (~io_in[0] & ~io_in[1] & io_in[5] & ~io_in[6] & ~io_in[8] & io_in[10]) | (~io_in[0] & ~io_in[2] & io_in[3] & ~io_in[4] & io_in[7] & io_in[8] & io_in[9]) | (io_in[0] & ~io_in[2] & io_in[6] & io_in[7] & ~io_in[8] & ~io_in[9] & io_in[10]) | (~io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[5] & io_in[6] & ~io_in[8] & io_in[9]) | (io_in[1] & ~io_in[3] & io_in[4] & io_in[7] & io_in[8] & io_in[9] & ~io_in[11]) | (~io_in[0] & ~io_in[3] & ~io_in[4] & ~io_in[6] & io_in[7] & ~io_in[8] & io_in[9] & ~io_in[11]) | (~io_in[0] & ~io_in[1] & io_in[3] & io_in[4] & io_in[6] & io_in[10] & ~io_in[11]) | (io_in[1] & ~io_in[3] & ~io_in[5] & ~io_in[6] & io_in[8] & io_in[9] & io_in[10] & ~io_in[11]) | (~io_in[2] & ~io_in[3] & ~io_in[4] & io_in[6] & ~io_in[7] & io_in[9] & io_in[10] & ~io_in[11]) | (~io_in[0] & io_in[3] & io_in[4] & io_in[6] & io_in[7] & ~io_in[9] & ~io_in[10]) | (io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[3] & io_in[6] & io_in[7] & ~io_in[8]) | (io_in[0] & ~io_in[1] & io_in[2] & io_in[4] & io_in[6] & ~io_in[9] & ~io_in[11]) | (io_in[0] & io_in[1] & ~io_in[4] & ~io_in[7] & ~io_in[8] & ~io_in[9] & ~io_in[10]) | (io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & ~io_in[6] & ~io_in[9] & ~io_in[10]) | (~io_in[0] & io_in[1] & io_in[3] & ~io_in[4] & io_in[7] & io_in[8] & io_in[9] & ~io_in[11]) | (~io_in[0] & io_in[1] & ~io_in[3] & io_in[4] & ~io_in[8] & ~io_in[9] & ~io_in[11]) | (~io_in[0] & ~io_in[1] & io_in[5] & ~io_in[8] & io_in[9]) | (~io_in[2] & ~io_in[3] & ~io_in[5] & io_in[7] & io_in[8] & io_in[9] & ~io_in[11]) | (io_in[0] & io_in[2] & ~io_in[4] & ~io_in[6] & io_in[7] & io_in[9] & io_in[11]) | (io_in[0] & io_in[2] & ~io_in[4] & ~io_in[5] & io_in[7] & io_in[8] & ~io_in[9]) | (~io_in[0] & io_in[1] & ~io_in[2] & ~io_in[3] & io_in[4] & ~io_in[6]) | (io_in[0] & ~io_in[1] & io_in[2] & ~io_in[4] & io_in[7] & io_in[10] & ~io_in[11]) | (io_in[0] & io_in[3] & io_in[5] & io_in[9] & ~io_in[11]) | (io_in[0] & ~io_in[2] & ~io_in[3] & io_in[6] & ~io_in[7] & ~io_in[8] & io_in[9]) | (io_in[1] & io_in[3] & ~io_in[4] & ~io_in[7] & ~io_in[9] & ~io_in[10] & ~io_in[11]) | (~io_in[1] & ~io_in[2] & ~io_in[3] & io_in[5] & io_in[6] & ~io_in[7] & io_in[9]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & ~io_in[5] & ~io_in[7] & io_in[8] & ~io_in[10] & ~io_in[11]) | (io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & io_in[7] & io_in[9] & ~io_in[10]) | (~io_in[0] & ~io_in[1] & ~io_in[3] & ~io_in[4] & ~io_in[7] & io_in[10] & ~io_in[11]) | (~io_in[0] & ~io_in[2] & ~io_in[4] & ~io_in[5] & io_in[7] & io_in[8] & io_in[9] & io_in[10]) | (~io_in[0] & ~io_in[1] & io_in[2] & ~io_in[3] & ~io_in[4] & ~io_in[10] & io_in[11]) | (io_in[1] & ~io_in[2] & io_in[3] & io_in[4] & io_in[7] & ~io_in[8] & ~io_in[10]) | (io_in[0] & ~io_in[2] & io_in[3] & ~io_in[4] & ~io_in[6] & ~io_in[7] & io_in[10]) | (~io_in[1] & io_in[2] & ~io_in[3] & ~io_in[6] & io_in[9] & ~io_in[10] & ~io_in[11]) | (~io_in[0] & ~io_in[1] & ~io_in[2] & io_in[3] & ~io_in[8] & ~io_in[9] & ~io_in[10]) | (~io_in[0] & io_in[1] & io_in[2] & io_in[3] & ~io_in[4] & io_in[6] & ~io_in[10]) | (~io_in[1] & io_in[2] & ~io_in[6] & ~io_in[7] & io_in[9] & ~io_in[11]) | (~io_in[1] & ~io_in[2] & ~io_in[5] & ~io_in[6] & ~io_in[8] & io_in[9] & ~io_in[10] & io_in[11]) | (~io_in[1] & io_in[2] & ~io_in[4] & io_in[5] & ~io_in[7] & io_in[11]) | (~io_in[1] & ~io_in[2] & ~io_in[3] & ~io_in[5] & io_in[6] & ~io_in[9] & ~io_in[10] & io_in[11]) | (io_in[2] & ~io_in[3] & io_in[5] & ~io_in[8] & ~io_in[9] & io_in[10]) | (io_in[0] & io_in[1] & ~io_in[2] & ~io_in[4] & io_in[7] & io_in[8] & io_in[9] & ~io_in[11]) | (io_in[1] & io_in[2] & io_in[3] & ~io_in[6] & ~io_in[7] & ~io_in[8]);

assign val[7] = 0;



endmodule
