module hex_to_sevenseg (
    input logic [3:0] hexdigit,
    output logic [7:0] seg
);

    always_comb begin
        seg = '1;
        if (hexdigit == 4'h0) seg = 8'b1100_0000;
        if (hexdigit == 4'h1) seg = 8'b1111_1001;
        if (hexdigit == 4'h2) seg = 8'b1010_0100;
        if (hexdigit == 4'h3) seg = 8'b1011_0000;
        if (hexdigit == 4'h4) seg = 8'b1001_1001;
        if (hexdigit == 4'h5) seg = 8'b1001_0010;
        if (hexdigit == 4'h6) seg = 8'b1000_0010;
        if (hexdigit == 4'h7) seg = 8'b1111_1000;
        if (hexdigit == 4'h8) seg = 8'b1000_0000;
        if (hexdigit == 4'h9) seg = 8'b1001_0000;
        if (hexdigit == 4'hA) seg = 8'b1000_1000;
        if (hexdigit == 4'hB) seg = 8'b1000_0011;
        if (hexdigit == 4'hC) seg = 8'b1100_0110;
        if (hexdigit == 4'hD) seg = 8'b1010_0001;
        if (hexdigit == 4'hE) seg = 8'b1000_0110;
        if (hexdigit == 4'hF) seg = 8'b1000_1110;
    end

endmodule

module m_design (
    input logic clk100, // 100MHz clock
    input logic reset_n, // Active-low reset

    output logic [7:0] base_led, // LEDs on the far right side of the board
    output logic [23:0] led, // LEDs in the middle of the board

    input logic [23:0] sw, // The tiny slide-switches
    input logic [4:0] btn, // The buttons

    output logic [3:0] display_sel, // Select between the 4 segments
    output logic [7:0] display // Seven-segment display
);

    logic clk; // 25MHz, generated by PLL

    // 100MHz -> 25MHz
    SB_PLL40_CORE #(
        .FEEDBACK_PATH("SIMPLE"),
        .DIVR(4'b0000),         // DIVR =  0
        .DIVF(7'b0000111),      // DIVF =  7
        .DIVQ(3'b101),          // DIVQ =  5
        .FILTER_RANGE(3'b101)   // FILTER_RANGE = 5
    ) pll (
        .LOCK(),
        .RESETB(1'b1),
        .BYPASS(1'b0),
        .REFERENCECLK(clk100),
        .PLLOUTCORE(clk)
    );
    
    logic [5:0] input_data;
    logic clock, reset, Next, Done;
    logic [10:0] display_out;
    logic Compute_done;

    logic [3:0] state;
    logic tape_reg_out, data_reg_out;
    logic [1:0] direction_out;
    logic [5:0] next_state_out, tape_addr_out;

    // Synchronizer sync0 (.async(btn[2]), .sync(clock), .clock(clk));
    Synchronizer sync1 (.async(btn[0]), .sync(Next), .clock(clk));
    Synchronizer sync2 (.async(btn[1]), .sync(Done), .clock(clk));
    Synchronizer sync3 (.async(sw[0]), .sync(input_data[0]), .clock(clk));
    Synchronizer sync4 (.async(sw[1]), .sync(input_data[1]), .clock(clk));
    Synchronizer sync5 (.async(sw[2]), .sync(input_data[2]), .clock(clk));
    Synchronizer sync6 (.async(sw[3]), .sync(input_data[3]), .clock(clk));
    Synchronizer sync7 (.async(sw[4]), .sync(input_data[4]), .clock(clk));
    Synchronizer sync8 (.async(sw[5]), .sync(input_data[5]), .clock(clk));
    
    TuringMachine TM (.*);

    assign clock = clk;
    assign reset = ~reset_n;
    // assign input_data = sw[3:0];
    assign led[10:0] = display_out;
    assign led[11] = Compute_done;

    hex_to_sevenseg hex(.hexdigit(state), .seg(display));
    assign display_sel = 4'b1110;

    assign base_led[0] = tape_reg_out;
    assign base_led[1] = data_reg_out;
    assign base_led[4:3] = direction_out;
    assign base_led[7:5] = next_state_out;
    assign led[23:18] = tape_addr_out;

    // assign led[15] = clock;
    assign led[14] = Done;
    assign led[13] = Next;

endmodule