`default_nettype none

module sbox(
    input logic [7:0] sbox_in,
    output logic [7:0] sbox_out
);

    logic [21 : 0] y;
    logic [67 : 0] t;
    logic [17 : 0] z;

    logic [7:0] s, u;
    assign u = sbox_in;
    assign sbox_out = s;

    always_comb begin
        y[14] = u[3] ^ u[5];
        y[13] = u[0] ^ u[6];
        y[9] = u[0] ^ u[3];
        y[8] = u[0] ^ u[5];
        t[0] = u[1] ^ u[2];
        y[1] = t[0] ^ u[7];
        y[4] = y[1] ^ u[3];
        y[12] = y[13] ^ y[14];
        y[2] = y[1] ^ u[0];
        y[5] = y[1] ^ u[6];
        y[3] = y[5] ^ y[8];
        t[1] = u[4] ^ y[12];
        y[15] = t[1] ^ u[5];
        y[20] = t[1] ^ u[1];
        y[6] = y[15] ^ u[7];
        y[10] = y[15] ^ t[0];
        y[11] = y[20] ^ y[9];
        y[7] = u[7] ^ y[11];
        y[17] = y[10] ^ y[11];
        y[19] = y[10] ^ y[8];
        y[16] = t[0] ^ y[11];
        y[21] = y[13] ^ y[16];
        y[18] = u[0] ^ y[16];
        t[2] = y[12] & y[15];
        t[3] = y[3] & y[6];
        t[4] = t[3] ^ t[2];
        t[5] = y[4] & u[7];
        t[6] = t[5] ^ t[2];
        t[7] = y[13] & y[16];
        t[8] = y[5] & y[1];
        t[9] = t[8] ^ t[7];
        t[10] = y[2] & y[7];
        t[11] = t[10] ^ t[7];
        t[12] = y[9] & y[11];
        t[13] = y[14] & y[17];
        t[14] = t[13] ^ t[12];
        t[15] = y[8] & y[10];
        t[16] = t[15] ^ t[12];
        t[17] = t[4] ^ t[14];
        t[18] = t[6] ^ t[16];
        t[19] = t[9] ^ t[14];
        t[20] = t[11] ^ t[16];
        t[21] = t[17] ^ y[20];
        t[22] = t[18] ^ y[19];
        t[23] = t[19] ^ y[21];
        t[24] = t[20] ^ y[18];
        t[25] = t[21] ^ t[22];
        t[26] = t[21] & t[23];
        t[27] = t[24] ^ t[26];
        t[28] = t[25] & t[27];
        t[29] = t[28] ^ t[22];
        t[30] = t[23] ^ t[24];
        t[31] = t[22] ^ t[26];
        t[32] = t[31] & t[30];
        t[33] = t[32] ^ t[24];
        t[34] = t[23] ^ t[33];
        t[35] = t[27] ^ t[33];
        t[36] = t[24] & t[35];
        t[37] = t[36] ^ t[34];
        t[38] = t[27] ^ t[36];
        t[39] = t[29] & t[38];
        t[40] = t[25] ^ t[39];
        t[41] = t[40] ^ t[37];
        t[42] = t[29] ^ t[33];
        t[43] = t[29] ^ t[40];
        t[44] = t[33] ^ t[37];
        t[45] = t[42] ^ t[41];
        z[0] = t[44] & y[15];
        z[1] = t[37] & y[6];
        z[2] = t[33] & u[7];
        z[3] = t[43] & y[16];
        z[4] = t[40] & y[1];
        z[5] = t[29] & y[7];
        z[6] = t[42] & y[11];
        z[7] = t[45] & y[17];
        z[8] = t[41] & y[10];
        z[9] = t[44] & y[12];
        z[10] = t[37] & y[3];
        z[11] = t[33] & y[4];
        z[12] = t[43] & y[13];
        z[13] = t[40] & y[5];
        z[14] = t[29] & y[2];
        z[15] = t[42] & y[9];
        z[16] = t[45] & y[14];
        z[17] = t[41] & y[8];
        t[46] = z[15] ^ z[16];
        t[47] = z[10] ^ z[11];
        t[48] = z[5] ^ z[13];
        t[49] = z[9] ^ z[10];
        t[50] = z[2] ^ z[12];
        t[51] = z[2] ^ z[5];
        t[52] = z[7] ^ z[8];
        t[53] = z[0] ^ z[3];
        t[54] = z[6] ^ z[7];
        t[55] = z[16] ^ z[17];
        t[56] = z[12] ^ t[48];
        t[57] = t[50] ^ t[53];
        t[58] = z[4] ^ t[46];
        t[59] = z[3] ^ t[54];
        t[60] = t[46] ^ t[57];
        t[61] = z[14] ^ t[57];
        t[62] = t[52] ^ t[58];
        t[63] = t[49] ^ t[58];
        t[64] = z[4] ^ t[59];
        t[65] = t[61] ^ t[62];
        t[66] = z[1] ^ t[63];
        s[0] = t[59] ^ t[63];
        s[6] = ~t[56] ^ t[62];
        s[7] = ~t[48] ^ t[60];
        t[67] = t[64] ^ t[65];
        s[3] = t[53] ^ t[66];
        s[4] = t[51] ^ t[66];
        s[5] = t[47] ^ t[65];
        s[1] = ~t[64] ^ s[3];
        s[2] = ~t[55] ^ t[67];
    end

endmodule

